module Queue(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_head,
  input         io_enq_bits_tail,
  input  [63:0] io_enq_bits_payload,
  input         io_enq_bits_flow_ingress_node,
  input         io_enq_bits_flow_egress_node,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_head,
  output        io_deq_bits_tail,
  output [63:0] io_deq_bits_payload,
  output        io_deq_bits_flow_ingress_node,
  output        io_deq_bits_flow_egress_node
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg  ram_head [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_head_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_head_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_head_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_tail [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_tail_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_tail_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_tail_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_en; // @[Decoupled.scala 273:95]
  reg [63:0] ram_payload [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_payload_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_payload_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [63:0] ram_payload_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [63:0] ram_payload_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_payload_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_payload_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_payload_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_flow_ingress_node [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_flow_ingress_node_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_flow_ingress_node_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_flow_ingress_node_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_flow_ingress_node_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_flow_ingress_node_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_flow_ingress_node_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_flow_ingress_node_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_flow_egress_node [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_flow_egress_node_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_flow_egress_node_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_flow_egress_node_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_flow_egress_node_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_flow_egress_node_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_flow_egress_node_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_flow_egress_node_MPORT_en; // @[Decoupled.scala 273:95]
  reg  enq_ptr_value; // @[Counter.scala 61:40]
  reg  deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  assign ram_head_io_deq_bits_MPORT_en = 1'h1;
  assign ram_head_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_head_io_deq_bits_MPORT_data = ram_head[ram_head_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_head_MPORT_data = io_enq_bits_head;
  assign ram_head_MPORT_addr = enq_ptr_value;
  assign ram_head_MPORT_mask = 1'h1;
  assign ram_head_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tail_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tail_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_tail_io_deq_bits_MPORT_data = ram_tail[ram_tail_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_tail_MPORT_data = io_enq_bits_tail;
  assign ram_tail_MPORT_addr = enq_ptr_value;
  assign ram_tail_MPORT_mask = 1'h1;
  assign ram_tail_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_payload_io_deq_bits_MPORT_en = 1'h1;
  assign ram_payload_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_payload_io_deq_bits_MPORT_data = ram_payload[ram_payload_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_payload_MPORT_data = io_enq_bits_payload;
  assign ram_payload_MPORT_addr = enq_ptr_value;
  assign ram_payload_MPORT_mask = 1'h1;
  assign ram_payload_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_flow_ingress_node_io_deq_bits_MPORT_en = 1'h1;
  assign ram_flow_ingress_node_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_flow_ingress_node_io_deq_bits_MPORT_data =
    ram_flow_ingress_node[ram_flow_ingress_node_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_flow_ingress_node_MPORT_data = io_enq_bits_flow_ingress_node;
  assign ram_flow_ingress_node_MPORT_addr = enq_ptr_value;
  assign ram_flow_ingress_node_MPORT_mask = 1'h1;
  assign ram_flow_ingress_node_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_flow_egress_node_io_deq_bits_MPORT_en = 1'h1;
  assign ram_flow_egress_node_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_flow_egress_node_io_deq_bits_MPORT_data = ram_flow_egress_node[ram_flow_egress_node_io_deq_bits_MPORT_addr]
    ; // @[Decoupled.scala 273:95]
  assign ram_flow_egress_node_MPORT_data = io_enq_bits_flow_egress_node;
  assign ram_flow_egress_node_MPORT_addr = enq_ptr_value;
  assign ram_flow_egress_node_MPORT_mask = 1'h1;
  assign ram_flow_egress_node_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_head = ram_head_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_tail = ram_tail_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_payload = ram_payload_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_flow_ingress_node = ram_flow_ingress_node_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_flow_egress_node = ram_flow_egress_node_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  always @(posedge clock) begin
    if (ram_head_MPORT_en & ram_head_MPORT_mask) begin
      ram_head[ram_head_MPORT_addr] <= ram_head_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_tail_MPORT_en & ram_tail_MPORT_mask) begin
      ram_tail[ram_tail_MPORT_addr] <= ram_tail_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_payload_MPORT_en & ram_payload_MPORT_mask) begin
      ram_payload[ram_payload_MPORT_addr] <= ram_payload_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_flow_ingress_node_MPORT_en & ram_flow_ingress_node_MPORT_mask) begin
      ram_flow_ingress_node[ram_flow_ingress_node_MPORT_addr] <= ram_flow_ingress_node_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_flow_egress_node_MPORT_en & ram_flow_egress_node_MPORT_mask) begin
      ram_flow_egress_node[ram_flow_egress_node_MPORT_addr] <= ram_flow_egress_node_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_head[initvar] = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_tail[initvar] = _RAND_1[0:0];
  _RAND_2 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload[initvar] = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_flow_ingress_node[initvar] = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_flow_egress_node[initvar] = _RAND_4[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  enq_ptr_value = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  deq_ptr_value = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  maybe_full = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_1(
  input   clock,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input   io_enq_bits_vc_sel_0_0,
  input   io_enq_bits_vc_sel_0_1,
  input   io_enq_bits_vc_sel_0_2,
  input   io_deq_ready,
  output  io_deq_valid,
  output  io_deq_bits_vc_sel_0_0,
  output  io_deq_bits_vc_sel_0_1,
  output  io_deq_bits_vc_sel_0_2
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg  ram_vc_sel_0_0 [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_0_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_0_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_0_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_0_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_0_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_0_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_vc_sel_0_1 [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_1_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_1_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_1_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_1_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_1_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_1_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_vc_sel_0_2 [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_2_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_2_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_2_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_2_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_2_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_2_MPORT_en; // @[Decoupled.scala 273:95]
  reg  enq_ptr_value; // @[Counter.scala 61:40]
  reg  deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  assign ram_vc_sel_0_0_io_deq_bits_MPORT_en = 1'h1;
  assign ram_vc_sel_0_0_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_vc_sel_0_0_io_deq_bits_MPORT_data = ram_vc_sel_0_0[ram_vc_sel_0_0_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_vc_sel_0_0_MPORT_data = io_enq_bits_vc_sel_0_0;
  assign ram_vc_sel_0_0_MPORT_addr = enq_ptr_value;
  assign ram_vc_sel_0_0_MPORT_mask = 1'h1;
  assign ram_vc_sel_0_0_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_vc_sel_0_1_io_deq_bits_MPORT_en = 1'h1;
  assign ram_vc_sel_0_1_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_vc_sel_0_1_io_deq_bits_MPORT_data = ram_vc_sel_0_1[ram_vc_sel_0_1_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_vc_sel_0_1_MPORT_data = io_enq_bits_vc_sel_0_1;
  assign ram_vc_sel_0_1_MPORT_addr = enq_ptr_value;
  assign ram_vc_sel_0_1_MPORT_mask = 1'h1;
  assign ram_vc_sel_0_1_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_vc_sel_0_2_io_deq_bits_MPORT_en = 1'h1;
  assign ram_vc_sel_0_2_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_vc_sel_0_2_io_deq_bits_MPORT_data = ram_vc_sel_0_2[ram_vc_sel_0_2_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_vc_sel_0_2_MPORT_data = io_enq_bits_vc_sel_0_2;
  assign ram_vc_sel_0_2_MPORT_addr = enq_ptr_value;
  assign ram_vc_sel_0_2_MPORT_mask = 1'h1;
  assign ram_vc_sel_0_2_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_vc_sel_0_0 = ram_vc_sel_0_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_vc_sel_0_1 = ram_vc_sel_0_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_vc_sel_0_2 = ram_vc_sel_0_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  always @(posedge clock) begin
    if (ram_vc_sel_0_0_MPORT_en & ram_vc_sel_0_0_MPORT_mask) begin
      ram_vc_sel_0_0[ram_vc_sel_0_0_MPORT_addr] <= ram_vc_sel_0_0_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_vc_sel_0_1_MPORT_en & ram_vc_sel_0_1_MPORT_mask) begin
      ram_vc_sel_0_1[ram_vc_sel_0_1_MPORT_addr] <= ram_vc_sel_0_1_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_vc_sel_0_2_MPORT_en & ram_vc_sel_0_2_MPORT_mask) begin
      ram_vc_sel_0_2[ram_vc_sel_0_2_MPORT_addr] <= ram_vc_sel_0_2_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_vc_sel_0_0[initvar] = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_vc_sel_0_1[initvar] = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_vc_sel_0_2[initvar] = _RAND_2[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  enq_ptr_value = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  deq_ptr_value = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  maybe_full = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_3(
  input   clock,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input   io_enq_bits_vc_sel_0_0,
  input   io_enq_bits_vc_sel_0_1,
  input   io_enq_bits_vc_sel_0_2,
  input   io_deq_ready,
  output  io_deq_valid,
  output  io_deq_bits_vc_sel_0_0,
  output  io_deq_bits_vc_sel_0_1,
  output  io_deq_bits_vc_sel_0_2
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg  ram_vc_sel_0_0 [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_0_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_0_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_0_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_0_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_0_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_0_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_vc_sel_0_1 [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_1_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_1_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_1_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_1_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_1_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_1_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_vc_sel_0_2 [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_2_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_2_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_2_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_2_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_2_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_2_MPORT_en; // @[Decoupled.scala 273:95]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 278:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  assign ram_vc_sel_0_0_io_deq_bits_MPORT_en = 1'h1;
  assign ram_vc_sel_0_0_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_vc_sel_0_0_io_deq_bits_MPORT_data = ram_vc_sel_0_0[ram_vc_sel_0_0_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_vc_sel_0_0_MPORT_data = io_enq_bits_vc_sel_0_0;
  assign ram_vc_sel_0_0_MPORT_addr = 1'h0;
  assign ram_vc_sel_0_0_MPORT_mask = 1'h1;
  assign ram_vc_sel_0_0_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_vc_sel_0_1_io_deq_bits_MPORT_en = 1'h1;
  assign ram_vc_sel_0_1_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_vc_sel_0_1_io_deq_bits_MPORT_data = ram_vc_sel_0_1[ram_vc_sel_0_1_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_vc_sel_0_1_MPORT_data = io_enq_bits_vc_sel_0_1;
  assign ram_vc_sel_0_1_MPORT_addr = 1'h0;
  assign ram_vc_sel_0_1_MPORT_mask = 1'h1;
  assign ram_vc_sel_0_1_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_vc_sel_0_2_io_deq_bits_MPORT_en = 1'h1;
  assign ram_vc_sel_0_2_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_vc_sel_0_2_io_deq_bits_MPORT_data = ram_vc_sel_0_2[ram_vc_sel_0_2_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_vc_sel_0_2_MPORT_data = io_enq_bits_vc_sel_0_2;
  assign ram_vc_sel_0_2_MPORT_addr = 1'h0;
  assign ram_vc_sel_0_2_MPORT_mask = 1'h1;
  assign ram_vc_sel_0_2_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = io_deq_ready | empty; // @[Decoupled.scala 303:16 323:{24,39}]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_vc_sel_0_0 = ram_vc_sel_0_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_vc_sel_0_1 = ram_vc_sel_0_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_vc_sel_0_2 = ram_vc_sel_0_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  always @(posedge clock) begin
    if (ram_vc_sel_0_0_MPORT_en & ram_vc_sel_0_0_MPORT_mask) begin
      ram_vc_sel_0_0[ram_vc_sel_0_0_MPORT_addr] <= ram_vc_sel_0_0_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_vc_sel_0_1_MPORT_en & ram_vc_sel_0_1_MPORT_mask) begin
      ram_vc_sel_0_1[ram_vc_sel_0_1_MPORT_addr] <= ram_vc_sel_0_1_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_vc_sel_0_2_MPORT_en & ram_vc_sel_0_2_MPORT_mask) begin
      ram_vc_sel_0_2[ram_vc_sel_0_2_MPORT_addr] <= ram_vc_sel_0_2_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_vc_sel_0_0[initvar] = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_vc_sel_0_1[initvar] = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_vc_sel_0_2[initvar] = _RAND_2[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IngressUnit(
  input         clock,
  input         reset,
  output        io_router_req_valid,
  input         io_vcalloc_req_ready,
  output        io_vcalloc_req_valid,
  output        io_vcalloc_req_bits_vc_sel_0_0,
  output        io_vcalloc_req_bits_vc_sel_0_1,
  output        io_vcalloc_req_bits_vc_sel_0_2,
  input         io_vcalloc_resp_vc_sel_0_0,
  input         io_vcalloc_resp_vc_sel_0_1,
  input         io_vcalloc_resp_vc_sel_0_2,
  input         io_out_credit_available_0_0,
  input         io_out_credit_available_0_1,
  input         io_out_credit_available_0_2,
  input         io_salloc_req_0_ready,
  output        io_salloc_req_0_valid,
  output        io_salloc_req_0_bits_vc_sel_0_0,
  output        io_salloc_req_0_bits_vc_sel_0_1,
  output        io_salloc_req_0_bits_vc_sel_0_2,
  output        io_salloc_req_0_bits_tail,
  output        io_out_0_valid,
  output        io_out_0_bits_flit_head,
  output        io_out_0_bits_flit_tail,
  output [63:0] io_out_0_bits_flit_payload,
  output        io_out_0_bits_flit_flow_ingress_node,
  output        io_out_0_bits_flit_flow_egress_node,
  output [1:0]  io_out_0_bits_out_virt_channel,
  output        io_in_ready,
  input         io_in_valid,
  input         io_in_bits_head,
  input         io_in_bits_tail,
  input  [63:0] io_in_bits_payload,
  input         io_in_bits_egress_id
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  route_buffer_clock; // @[IngressUnit.scala 26:28]
  wire  route_buffer_reset; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_enq_ready; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_enq_valid; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_enq_bits_head; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_enq_bits_tail; // @[IngressUnit.scala 26:28]
  wire [63:0] route_buffer_io_enq_bits_payload; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_enq_bits_flow_ingress_node; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_enq_bits_flow_egress_node; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_deq_ready; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_deq_valid; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_deq_bits_head; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_deq_bits_tail; // @[IngressUnit.scala 26:28]
  wire [63:0] route_buffer_io_deq_bits_payload; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_deq_bits_flow_ingress_node; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_deq_bits_flow_egress_node; // @[IngressUnit.scala 26:28]
  wire  route_q_clock; // @[IngressUnit.scala 27:23]
  wire  route_q_reset; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_ready; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_valid; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_0_0; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_0_1; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_0_2; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_ready; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_valid; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_0_0; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_0_1; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_0_2; // @[IngressUnit.scala 27:23]
  wire  vcalloc_buffer_clock; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_reset; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_enq_ready; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_enq_valid; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_enq_bits_head; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_enq_bits_tail; // @[IngressUnit.scala 75:30]
  wire [63:0] vcalloc_buffer_io_enq_bits_payload; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_enq_bits_flow_ingress_node; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_enq_bits_flow_egress_node; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_deq_ready; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_deq_valid; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_deq_bits_head; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_deq_bits_tail; // @[IngressUnit.scala 75:30]
  wire [63:0] vcalloc_buffer_io_deq_bits_payload; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_deq_bits_flow_ingress_node; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_deq_bits_flow_egress_node; // @[IngressUnit.scala 75:30]
  wire  vcalloc_q_clock; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_reset; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_ready; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_valid; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_0_0; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_0_1; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_0_2; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_ready; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_valid; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_0_0; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_0_1; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_0_2; // @[IngressUnit.scala 76:25]
  wire  _T_5 = ~reset; // @[IngressUnit.scala 30:9]
  wire  at_dest = ~route_buffer_io_enq_bits_flow_egress_node; // @[IngressUnit.scala 55:59]
  wire  _T_7 = io_in_ready & io_in_valid; // @[Decoupled.scala 51:35]
  wire  _vcalloc_buffer_io_enq_valid_T = ~route_buffer_io_deq_bits_head; // @[IngressUnit.scala 88:30]
  wire  _vcalloc_buffer_io_enq_valid_T_1 = route_q_io_deq_valid | ~route_buffer_io_deq_bits_head; // @[IngressUnit.scala 88:27]
  wire  _vcalloc_buffer_io_enq_valid_T_2 = route_buffer_io_deq_valid & _vcalloc_buffer_io_enq_valid_T_1; // @[IngressUnit.scala 87:61]
  wire  _vcalloc_buffer_io_enq_valid_T_4 = io_vcalloc_req_ready | _vcalloc_buffer_io_enq_valid_T; // @[IngressUnit.scala 89:27]
  wire  _io_vcalloc_req_valid_T_1 = route_buffer_io_deq_valid & route_q_io_deq_valid & route_buffer_io_deq_bits_head; // @[IngressUnit.scala 91:78]
  wire  _route_buffer_io_deq_ready_T_2 = vcalloc_buffer_io_enq_ready & _vcalloc_buffer_io_enq_valid_T_1; // @[IngressUnit.scala 93:61]
  wire  _route_buffer_io_deq_ready_T_5 = _route_buffer_io_deq_ready_T_2 & _vcalloc_buffer_io_enq_valid_T_4; // @[IngressUnit.scala 94:37]
  wire  _route_buffer_io_deq_ready_T_7 = vcalloc_q_io_enq_ready | _vcalloc_buffer_io_enq_valid_T; // @[IngressUnit.scala 96:29]
  wire  _route_q_io_deq_ready_T = route_buffer_io_deq_ready & route_buffer_io_deq_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _c_T = {vcalloc_q_io_deq_bits_vc_sel_0_2,vcalloc_q_io_deq_bits_vc_sel_0_1,vcalloc_q_io_deq_bits_vc_sel_0_0}
    ; // @[IngressUnit.scala 107:41]
  wire [2:0] _c_T_1 = {io_out_credit_available_0_2,io_out_credit_available_0_1,io_out_credit_available_0_0}; // @[IngressUnit.scala 107:74]
  wire [2:0] _c_T_2 = _c_T & _c_T_1; // @[IngressUnit.scala 107:48]
  wire  c = _c_T_2 != 3'h0; // @[IngressUnit.scala 107:82]
  wire  _vcalloc_q_io_deq_ready_T = vcalloc_buffer_io_deq_ready & vcalloc_buffer_io_deq_valid; // @[Decoupled.scala 51:35]
  reg  out_bundle_valid; // @[IngressUnit.scala 116:8]
  reg  out_bundle_bits_flit_head; // @[IngressUnit.scala 116:8]
  reg  out_bundle_bits_flit_tail; // @[IngressUnit.scala 116:8]
  reg [63:0] out_bundle_bits_flit_payload; // @[IngressUnit.scala 116:8]
  reg  out_bundle_bits_flit_flow_ingress_node; // @[IngressUnit.scala 116:8]
  reg  out_bundle_bits_flit_flow_egress_node; // @[IngressUnit.scala 116:8]
  reg [1:0] out_bundle_bits_out_virt_channel; // @[IngressUnit.scala 116:8]
  wire  out_bundle_bits_out_virt_channel_hi_1 = _c_T[2]; // @[OneHot.scala 30:18]
  wire [1:0] out_bundle_bits_out_virt_channel_lo = _c_T[1:0]; // @[OneHot.scala 31:18]
  wire  _out_bundle_bits_out_virt_channel_T_1 = |out_bundle_bits_out_virt_channel_hi_1; // @[OneHot.scala 32:14]
  wire [1:0] _GEN_4 = {{1'd0}, out_bundle_bits_out_virt_channel_hi_1}; // @[OneHot.scala 32:28]
  wire [1:0] _out_bundle_bits_out_virt_channel_T_2 = _GEN_4 | out_bundle_bits_out_virt_channel_lo; // @[OneHot.scala 32:28]
  Queue route_buffer ( // @[IngressUnit.scala 26:28]
    .clock(route_buffer_clock),
    .reset(route_buffer_reset),
    .io_enq_ready(route_buffer_io_enq_ready),
    .io_enq_valid(route_buffer_io_enq_valid),
    .io_enq_bits_head(route_buffer_io_enq_bits_head),
    .io_enq_bits_tail(route_buffer_io_enq_bits_tail),
    .io_enq_bits_payload(route_buffer_io_enq_bits_payload),
    .io_enq_bits_flow_ingress_node(route_buffer_io_enq_bits_flow_ingress_node),
    .io_enq_bits_flow_egress_node(route_buffer_io_enq_bits_flow_egress_node),
    .io_deq_ready(route_buffer_io_deq_ready),
    .io_deq_valid(route_buffer_io_deq_valid),
    .io_deq_bits_head(route_buffer_io_deq_bits_head),
    .io_deq_bits_tail(route_buffer_io_deq_bits_tail),
    .io_deq_bits_payload(route_buffer_io_deq_bits_payload),
    .io_deq_bits_flow_ingress_node(route_buffer_io_deq_bits_flow_ingress_node),
    .io_deq_bits_flow_egress_node(route_buffer_io_deq_bits_flow_egress_node)
  );
  Queue_1 route_q ( // @[IngressUnit.scala 27:23]
    .clock(route_q_clock),
    .reset(route_q_reset),
    .io_enq_ready(route_q_io_enq_ready),
    .io_enq_valid(route_q_io_enq_valid),
    .io_enq_bits_vc_sel_0_0(route_q_io_enq_bits_vc_sel_0_0),
    .io_enq_bits_vc_sel_0_1(route_q_io_enq_bits_vc_sel_0_1),
    .io_enq_bits_vc_sel_0_2(route_q_io_enq_bits_vc_sel_0_2),
    .io_deq_ready(route_q_io_deq_ready),
    .io_deq_valid(route_q_io_deq_valid),
    .io_deq_bits_vc_sel_0_0(route_q_io_deq_bits_vc_sel_0_0),
    .io_deq_bits_vc_sel_0_1(route_q_io_deq_bits_vc_sel_0_1),
    .io_deq_bits_vc_sel_0_2(route_q_io_deq_bits_vc_sel_0_2)
  );
  Queue vcalloc_buffer ( // @[IngressUnit.scala 75:30]
    .clock(vcalloc_buffer_clock),
    .reset(vcalloc_buffer_reset),
    .io_enq_ready(vcalloc_buffer_io_enq_ready),
    .io_enq_valid(vcalloc_buffer_io_enq_valid),
    .io_enq_bits_head(vcalloc_buffer_io_enq_bits_head),
    .io_enq_bits_tail(vcalloc_buffer_io_enq_bits_tail),
    .io_enq_bits_payload(vcalloc_buffer_io_enq_bits_payload),
    .io_enq_bits_flow_ingress_node(vcalloc_buffer_io_enq_bits_flow_ingress_node),
    .io_enq_bits_flow_egress_node(vcalloc_buffer_io_enq_bits_flow_egress_node),
    .io_deq_ready(vcalloc_buffer_io_deq_ready),
    .io_deq_valid(vcalloc_buffer_io_deq_valid),
    .io_deq_bits_head(vcalloc_buffer_io_deq_bits_head),
    .io_deq_bits_tail(vcalloc_buffer_io_deq_bits_tail),
    .io_deq_bits_payload(vcalloc_buffer_io_deq_bits_payload),
    .io_deq_bits_flow_ingress_node(vcalloc_buffer_io_deq_bits_flow_ingress_node),
    .io_deq_bits_flow_egress_node(vcalloc_buffer_io_deq_bits_flow_egress_node)
  );
  Queue_3 vcalloc_q ( // @[IngressUnit.scala 76:25]
    .clock(vcalloc_q_clock),
    .reset(vcalloc_q_reset),
    .io_enq_ready(vcalloc_q_io_enq_ready),
    .io_enq_valid(vcalloc_q_io_enq_valid),
    .io_enq_bits_vc_sel_0_0(vcalloc_q_io_enq_bits_vc_sel_0_0),
    .io_enq_bits_vc_sel_0_1(vcalloc_q_io_enq_bits_vc_sel_0_1),
    .io_enq_bits_vc_sel_0_2(vcalloc_q_io_enq_bits_vc_sel_0_2),
    .io_deq_ready(vcalloc_q_io_deq_ready),
    .io_deq_valid(vcalloc_q_io_deq_valid),
    .io_deq_bits_vc_sel_0_0(vcalloc_q_io_deq_bits_vc_sel_0_0),
    .io_deq_bits_vc_sel_0_1(vcalloc_q_io_deq_bits_vc_sel_0_1),
    .io_deq_bits_vc_sel_0_2(vcalloc_q_io_deq_bits_vc_sel_0_2)
  );
  assign io_router_req_valid = io_in_valid & route_buffer_io_enq_ready & io_in_bits_head & ~at_dest; // @[IngressUnit.scala 58:86]
  assign io_vcalloc_req_valid = _io_vcalloc_req_valid_T_1 & vcalloc_buffer_io_enq_ready & vcalloc_q_io_enq_ready; // @[IngressUnit.scala 92:41]
  assign io_vcalloc_req_bits_vc_sel_0_0 = route_q_io_deq_bits_vc_sel_0_0; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_0_1 = route_q_io_deq_bits_vc_sel_0_1; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_0_2 = route_q_io_deq_bits_vc_sel_0_2; // @[IngressUnit.scala 81:30]
  assign io_salloc_req_0_valid = vcalloc_buffer_io_deq_valid & vcalloc_q_io_deq_valid & c; // @[IngressUnit.scala 109:83]
  assign io_salloc_req_0_bits_vc_sel_0_0 = vcalloc_q_io_deq_bits_vc_sel_0_0; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_0_1 = vcalloc_q_io_deq_bits_vc_sel_0_1; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_0_2 = vcalloc_q_io_deq_bits_vc_sel_0_2; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_tail = vcalloc_buffer_io_deq_bits_tail; // @[IngressUnit.scala 105:30]
  assign io_out_0_valid = out_bundle_valid; // @[IngressUnit.scala 118:13]
  assign io_out_0_bits_flit_head = out_bundle_bits_flit_head; // @[IngressUnit.scala 118:13]
  assign io_out_0_bits_flit_tail = out_bundle_bits_flit_tail; // @[IngressUnit.scala 118:13]
  assign io_out_0_bits_flit_payload = out_bundle_bits_flit_payload; // @[IngressUnit.scala 118:13]
  assign io_out_0_bits_flit_flow_ingress_node = out_bundle_bits_flit_flow_ingress_node; // @[IngressUnit.scala 118:13]
  assign io_out_0_bits_flit_flow_egress_node = out_bundle_bits_flit_flow_egress_node; // @[IngressUnit.scala 118:13]
  assign io_out_0_bits_out_virt_channel = out_bundle_bits_out_virt_channel; // @[IngressUnit.scala 118:13]
  assign io_in_ready = route_buffer_io_enq_ready; // @[IngressUnit.scala 59:44]
  assign route_buffer_clock = clock;
  assign route_buffer_reset = reset;
  assign route_buffer_io_enq_valid = io_in_valid; // @[IngressUnit.scala 56:44]
  assign route_buffer_io_enq_bits_head = io_in_bits_head; // @[IngressUnit.scala 32:33]
  assign route_buffer_io_enq_bits_tail = io_in_bits_tail; // @[IngressUnit.scala 33:33]
  assign route_buffer_io_enq_bits_payload = io_in_bits_payload; // @[IngressUnit.scala 50:36]
  assign route_buffer_io_enq_bits_flow_ingress_node = 1'h0; // @[IngressUnit.scala 38:51]
  assign route_buffer_io_enq_bits_flow_egress_node = 1'h1; // @[IngressUnit.scala 41:50]
  assign route_buffer_io_deq_ready = _route_buffer_io_deq_ready_T_5 & _route_buffer_io_deq_ready_T_7; // @[IngressUnit.scala 95:37]
  assign route_q_clock = clock;
  assign route_q_reset = reset;
  assign route_q_io_enq_valid = _T_7 & io_in_bits_head & at_dest | io_router_req_valid; // @[IngressUnit.scala 62:24 64:53 65:26]
  assign route_q_io_enq_bits_vc_sel_0_0 = _T_7 & io_in_bits_head & at_dest ? 1'h0 : 1'h1; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_0_1 = _T_7 & io_in_bits_head & at_dest ? 1'h0 : 1'h1; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_0_2 = _T_7 & io_in_bits_head & at_dest ? 1'h0 : 1'h1; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_deq_ready = _route_q_io_deq_ready_T & route_buffer_io_deq_bits_tail; // @[IngressUnit.scala 97:55]
  assign vcalloc_buffer_clock = clock;
  assign vcalloc_buffer_reset = reset;
  assign vcalloc_buffer_io_enq_valid = _vcalloc_buffer_io_enq_valid_T_2 & _vcalloc_buffer_io_enq_valid_T_4; // @[IngressUnit.scala 88:37]
  assign vcalloc_buffer_io_enq_bits_head = route_buffer_io_deq_bits_head; // @[IngressUnit.scala 79:30]
  assign vcalloc_buffer_io_enq_bits_tail = route_buffer_io_deq_bits_tail; // @[IngressUnit.scala 79:30]
  assign vcalloc_buffer_io_enq_bits_payload = route_buffer_io_deq_bits_payload; // @[IngressUnit.scala 79:30]
  assign vcalloc_buffer_io_enq_bits_flow_ingress_node = route_buffer_io_deq_bits_flow_ingress_node; // @[IngressUnit.scala 79:30]
  assign vcalloc_buffer_io_enq_bits_flow_egress_node = route_buffer_io_deq_bits_flow_egress_node; // @[IngressUnit.scala 79:30]
  assign vcalloc_buffer_io_deq_ready = io_salloc_req_0_ready & vcalloc_q_io_deq_valid & c; // @[IngressUnit.scala 110:83]
  assign vcalloc_q_clock = clock;
  assign vcalloc_q_reset = reset;
  assign vcalloc_q_io_enq_valid = io_vcalloc_req_ready & io_vcalloc_req_valid; // @[Decoupled.scala 51:35]
  assign vcalloc_q_io_enq_bits_vc_sel_0_0 = io_vcalloc_resp_vc_sel_0_0; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_0_1 = io_vcalloc_resp_vc_sel_0_1; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_0_2 = io_vcalloc_resp_vc_sel_0_2; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_deq_ready = vcalloc_buffer_io_deq_bits_tail & _vcalloc_q_io_deq_ready_T; // @[IngressUnit.scala 111:42]
  always @(posedge clock) begin
    out_bundle_valid <= vcalloc_buffer_io_deq_ready & vcalloc_buffer_io_deq_valid; // @[Decoupled.scala 51:35]
    out_bundle_bits_flit_head <= vcalloc_buffer_io_deq_bits_head; // @[IngressUnit.scala 121:24]
    out_bundle_bits_flit_tail <= vcalloc_buffer_io_deq_bits_tail; // @[IngressUnit.scala 121:24]
    out_bundle_bits_flit_payload <= vcalloc_buffer_io_deq_bits_payload; // @[IngressUnit.scala 121:24]
    out_bundle_bits_flit_flow_ingress_node <= vcalloc_buffer_io_deq_bits_flow_ingress_node; // @[IngressUnit.scala 121:24]
    out_bundle_bits_flit_flow_egress_node <= vcalloc_buffer_io_deq_bits_flow_egress_node; // @[IngressUnit.scala 121:24]
    out_bundle_bits_out_virt_channel <= {_out_bundle_bits_out_virt_channel_T_1,_out_bundle_bits_out_virt_channel_T_2[1]}
      ; // @[Cat.scala 33:92]
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~(io_in_valid & ~(~io_in_bits_egress_id)))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at IngressUnit.scala:30 assert(!(io.in.valid && !cParam.possibleFlows.toSeq.map(_.egressId.U === io.in.bits.egress_id).orR))\n"
            ); // @[IngressUnit.scala 30:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5 & ~(~(route_q_io_enq_valid & ~route_q_io_enq_ready))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at IngressUnit.scala:73 assert(!(route_q.io.enq.valid && !route_q.io.enq.ready))\n"); // @[IngressUnit.scala 73:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5 & ~(~(vcalloc_q_io_enq_valid & ~vcalloc_q_io_enq_ready))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at IngressUnit.scala:102 assert(!(vcalloc_q.io.enq.valid && !vcalloc_q.io.enq.ready))\n"
            ); // @[IngressUnit.scala 102:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  out_bundle_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  out_bundle_bits_flit_head = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  out_bundle_bits_flit_tail = _RAND_2[0:0];
  _RAND_3 = {2{`RANDOM}};
  out_bundle_bits_flit_payload = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  out_bundle_bits_flit_flow_ingress_node = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  out_bundle_bits_flit_flow_egress_node = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  out_bundle_bits_out_virt_channel = _RAND_6[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(~(io_in_valid & ~(~io_in_bits_egress_id))); // @[IngressUnit.scala 30:9]
    end
    //
    if (_T_5) begin
      assert(~(route_q_io_enq_valid & ~route_q_io_enq_ready)); // @[IngressUnit.scala 73:9]
    end
    //
    if (_T_5) begin
      assert(~(vcalloc_q_io_enq_valid & ~vcalloc_q_io_enq_ready)); // @[IngressUnit.scala 102:9]
    end
  end
endmodule
module OutputUnit(
  input         clock,
  input         reset,
  input         io_in_0_valid,
  input         io_in_0_bits_head,
  input         io_in_0_bits_tail,
  input  [63:0] io_in_0_bits_payload,
  input         io_in_0_bits_flow_ingress_node,
  input         io_in_0_bits_flow_egress_node,
  input  [1:0]  io_in_0_bits_virt_channel_id,
  output        io_credit_available_0,
  output        io_credit_available_1,
  output        io_credit_available_2,
  output        io_channel_status_0_occupied,
  output        io_channel_status_1_occupied,
  output        io_channel_status_2_occupied,
  input         io_allocs_0_alloc,
  input         io_allocs_1_alloc,
  input         io_allocs_2_alloc,
  input         io_credit_alloc_0_alloc,
  input         io_credit_alloc_1_alloc,
  input         io_credit_alloc_2_alloc,
  output        io_out_flit_0_valid,
  output        io_out_flit_0_bits_head,
  output        io_out_flit_0_bits_tail,
  output [63:0] io_out_flit_0_bits_payload,
  output        io_out_flit_0_bits_flow_ingress_node,
  output        io_out_flit_0_bits_flow_egress_node,
  output [1:0]  io_out_flit_0_bits_virt_channel_id,
  input  [2:0]  io_out_credit_return,
  input  [2:0]  io_out_vc_free
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg  states_2_occupied; // @[OutputUnit.scala 66:19]
  reg [1:0] states_2_c; // @[OutputUnit.scala 66:19]
  reg  states_1_occupied; // @[OutputUnit.scala 66:19]
  reg [1:0] states_1_c; // @[OutputUnit.scala 66:19]
  reg  states_0_occupied; // @[OutputUnit.scala 66:19]
  reg [1:0] states_0_c; // @[OutputUnit.scala 66:19]
  wire  _GEN_0 = io_out_vc_free[0] ? 1'h0 : states_0_occupied; // @[OutputUnit.scala 74:30 76:18 66:19]
  wire  _GEN_1 = io_out_vc_free[1] ? 1'h0 : states_1_occupied; // @[OutputUnit.scala 74:30 76:18 66:19]
  wire  _GEN_2 = io_out_vc_free[2] ? 1'h0 : states_2_occupied; // @[OutputUnit.scala 74:30 76:18 66:19]
  wire  _GEN_3 = io_allocs_0_alloc | _GEN_0; // @[OutputUnit.scala 83:20 84:18]
  wire  _GEN_9 = io_allocs_1_alloc | _GEN_1; // @[OutputUnit.scala 83:20 84:18]
  wire  _GEN_15 = io_allocs_2_alloc | _GEN_2; // @[OutputUnit.scala 83:20 84:18]
  wire  free = io_out_credit_return[0]; // @[OutputUnit.scala 94:36]
  wire [1:0] _GEN_4 = {{1'd0}, free}; // @[OutputUnit.scala 97:18]
  wire [2:0] _states_0_c_T = states_0_c + _GEN_4; // @[OutputUnit.scala 97:18]
  wire [2:0] _GEN_6 = {{2'd0}, io_credit_alloc_0_alloc}; // @[OutputUnit.scala 97:26]
  wire [2:0] _states_0_c_T_2 = _states_0_c_T - _GEN_6; // @[OutputUnit.scala 97:26]
  wire  free_1 = io_out_credit_return[1]; // @[OutputUnit.scala 94:36]
  wire [1:0] _GEN_8 = {{1'd0}, free_1}; // @[OutputUnit.scala 97:18]
  wire [2:0] _states_1_c_T = states_1_c + _GEN_8; // @[OutputUnit.scala 97:18]
  wire [2:0] _GEN_10 = {{2'd0}, io_credit_alloc_1_alloc}; // @[OutputUnit.scala 97:26]
  wire [2:0] _states_1_c_T_2 = _states_1_c_T - _GEN_10; // @[OutputUnit.scala 97:26]
  wire  free_2 = io_out_credit_return[2]; // @[OutputUnit.scala 94:36]
  wire [1:0] _GEN_12 = {{1'd0}, free_2}; // @[OutputUnit.scala 97:18]
  wire [2:0] _states_2_c_T = states_2_c + _GEN_12; // @[OutputUnit.scala 97:18]
  wire [2:0] _GEN_14 = {{2'd0}, io_credit_alloc_2_alloc}; // @[OutputUnit.scala 97:26]
  wire [2:0] _states_2_c_T_2 = _states_2_c_T - _GEN_14; // @[OutputUnit.scala 97:26]
  wire [2:0] _GEN_24 = reset ? 3'h3 : _states_0_c_T_2; // @[OutputUnit.scala 103:23 105:29 97:11]
  wire [2:0] _GEN_25 = reset ? 3'h3 : _states_1_c_T_2; // @[OutputUnit.scala 103:23 105:29 97:11]
  wire [2:0] _GEN_26 = reset ? 3'h3 : _states_2_c_T_2; // @[OutputUnit.scala 103:23 105:29 97:11]
  assign io_credit_available_0 = states_0_c != 2'h0; // @[OutputUnit.scala 90:14]
  assign io_credit_available_1 = states_1_c != 2'h0; // @[OutputUnit.scala 90:14]
  assign io_credit_available_2 = states_2_c != 2'h0; // @[OutputUnit.scala 90:14]
  assign io_channel_status_0_occupied = io_out_vc_free[0] ? 1'h0 : states_0_occupied; // @[OutputUnit.scala 74:30 76:18 66:19]
  assign io_channel_status_1_occupied = io_out_vc_free[1] ? 1'h0 : states_1_occupied; // @[OutputUnit.scala 74:30 76:18 66:19]
  assign io_channel_status_2_occupied = io_out_vc_free[2] ? 1'h0 : states_2_occupied; // @[OutputUnit.scala 74:30 76:18 66:19]
  assign io_out_flit_0_valid = io_in_0_valid; // @[OutputUnit.scala 71:15]
  assign io_out_flit_0_bits_head = io_in_0_bits_head; // @[OutputUnit.scala 71:15]
  assign io_out_flit_0_bits_tail = io_in_0_bits_tail; // @[OutputUnit.scala 71:15]
  assign io_out_flit_0_bits_payload = io_in_0_bits_payload; // @[OutputUnit.scala 71:15]
  assign io_out_flit_0_bits_flow_ingress_node = io_in_0_bits_flow_ingress_node; // @[OutputUnit.scala 71:15]
  assign io_out_flit_0_bits_flow_egress_node = io_in_0_bits_flow_egress_node; // @[OutputUnit.scala 71:15]
  assign io_out_flit_0_bits_virt_channel_id = io_in_0_bits_virt_channel_id; // @[OutputUnit.scala 71:15]
  always @(posedge clock) begin
    if (reset) begin // @[OutputUnit.scala 103:23]
      states_2_occupied <= 1'h0; // @[OutputUnit.scala 104:31]
    end else begin
      states_2_occupied <= _GEN_15;
    end
    states_2_c <= _GEN_26[1:0];
    if (reset) begin // @[OutputUnit.scala 103:23]
      states_1_occupied <= 1'h0; // @[OutputUnit.scala 104:31]
    end else begin
      states_1_occupied <= _GEN_9;
    end
    states_1_c <= _GEN_25[1:0];
    if (reset) begin // @[OutputUnit.scala 103:23]
      states_0_occupied <= 1'h0; // @[OutputUnit.scala 104:31]
    end else begin
      states_0_occupied <= _GEN_3;
    end
    states_0_c <= _GEN_24[1:0];
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_out_vc_free[0] & ~reset & ~states_0_occupied) begin
          $fwrite(32'h80000002,"Assertion failed\n    at OutputUnit.scala:75 assert(s.occupied)\n"); // @[OutputUnit.scala 75:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_out_vc_free[1] & ~reset & ~states_1_occupied) begin
          $fwrite(32'h80000002,"Assertion failed\n    at OutputUnit.scala:75 assert(s.occupied)\n"); // @[OutputUnit.scala 75:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_out_vc_free[2] & ~reset & ~states_2_occupied) begin
          $fwrite(32'h80000002,"Assertion failed\n    at OutputUnit.scala:75 assert(s.occupied)\n"); // @[OutputUnit.scala 75:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  states_2_occupied = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  states_2_c = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  states_1_occupied = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  states_1_c = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  states_0_occupied = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  states_0_c = _RAND_5[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (io_out_vc_free[0] & ~reset) begin
      assert(states_0_occupied); // @[OutputUnit.scala 75:13]
    end
    //
    if (io_out_vc_free[1] & ~reset) begin
      assert(states_1_occupied); // @[OutputUnit.scala 75:13]
    end
    //
    if (io_out_vc_free[2] & ~reset) begin
      assert(states_2_occupied); // @[OutputUnit.scala 75:13]
    end
  end
endmodule
module Switch(
  input         clock,
  input         reset,
  input         io_in_0_0_valid,
  input         io_in_0_0_bits_flit_head,
  input         io_in_0_0_bits_flit_tail,
  input  [63:0] io_in_0_0_bits_flit_payload,
  input         io_in_0_0_bits_flit_flow_ingress_node,
  input         io_in_0_0_bits_flit_flow_egress_node,
  input  [1:0]  io_in_0_0_bits_out_virt_channel,
  output        io_out_0_0_valid,
  output        io_out_0_0_bits_head,
  output        io_out_0_0_bits_tail,
  output [63:0] io_out_0_0_bits_payload,
  output        io_out_0_0_bits_flow_ingress_node,
  output        io_out_0_0_bits_flow_egress_node,
  output [1:0]  io_out_0_0_bits_virt_channel_id,
  input         io_sel_0_0_0_0
);
  assign io_out_0_0_valid = io_in_0_0_valid & io_sel_0_0_0_0; // @[Switch.scala 48:67]
  assign io_out_0_0_bits_head = io_in_0_0_bits_flit_head; // @[Switch.scala 36:21 40:18]
  assign io_out_0_0_bits_tail = io_in_0_0_bits_flit_tail; // @[Switch.scala 36:21 40:18]
  assign io_out_0_0_bits_payload = io_in_0_0_bits_flit_payload; // @[Switch.scala 36:21 40:18]
  assign io_out_0_0_bits_flow_ingress_node = io_in_0_0_bits_flit_flow_ingress_node; // @[Switch.scala 36:21 40:18]
  assign io_out_0_0_bits_flow_egress_node = io_in_0_0_bits_flit_flow_egress_node; // @[Switch.scala 36:21 40:18]
  assign io_out_0_0_bits_virt_channel_id = io_in_0_0_bits_out_virt_channel; // @[Switch.scala 36:21 40:18]
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(1'h1); // @[Switch.scala 47:13]
    end
  end
endmodule
module SwitchArbiter(
  input   clock,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input   io_in_0_bits_vc_sel_0_0,
  input   io_in_0_bits_vc_sel_0_1,
  input   io_in_0_bits_vc_sel_0_2,
  input   io_in_0_bits_tail,
  output  io_out_0_valid,
  output  io_out_0_bits_vc_sel_0_0,
  output  io_out_0_bits_vc_sel_0_1,
  output  io_out_0_bits_vc_sel_0_2,
  output  io_chosen_oh_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  lock_0; // @[SwitchAllocator.scala 24:38]
  wire  unassigned = io_in_0_valid & ~lock_0; // @[SwitchAllocator.scala 25:52]
  reg  mask; // @[SwitchAllocator.scala 27:21]
  wire  _sel_T = ~mask; // @[SwitchAllocator.scala 30:60]
  wire  _sel_T_1 = unassigned & ~mask; // @[SwitchAllocator.scala 30:58]
  wire [1:0] _sel_T_2 = {unassigned,_sel_T_1}; // @[Cat.scala 33:92]
  wire [1:0] _sel_T_5 = _sel_T_2[1] ? 2'h2 : 2'h0; // @[Mux.scala 47:70]
  wire [1:0] sel = _sel_T_2[0] ? 2'h1 : _sel_T_5; // @[Mux.scala 47:70]
  wire [1:0] _GEN_3 = {{1'd0}, sel[1]}; // @[SwitchAllocator.scala 32:23]
  wire [1:0] _choices_0_T_1 = sel | _GEN_3; // @[SwitchAllocator.scala 32:23]
  wire  choices_0 = _choices_0_T_1[0]; // @[SwitchAllocator.scala 28:21 32:16]
  wire  chosen = |(io_in_0_valid & lock_0) ? lock_0 : choices_0; // @[SwitchAllocator.scala 42:21]
  wire [1:0] _mask_T_3 = {mask, 1'h0}; // @[SwitchAllocator.scala 60:43]
  wire [1:0] _mask_T_4 = _mask_T_3 | 2'h1; // @[SwitchAllocator.scala 60:49]
  wire [1:0] _mask_T_5 = ~_sel_T ? 2'h0 : _mask_T_4; // @[SwitchAllocator.scala 60:16]
  wire [1:0] _GEN_2 = io_out_0_valid ? {{1'd0}, io_chosen_oh_0} : _mask_T_5; // @[SwitchAllocator.scala 57:27 58:10 60:10]
  wire [1:0] _GEN_4 = reset ? 2'h0 : _GEN_2; // @[SwitchAllocator.scala 27:{21,21}]
  assign io_in_0_ready = |(io_in_0_valid & lock_0) ? lock_0 : choices_0; // @[SwitchAllocator.scala 42:21]
  assign io_out_0_valid = |(io_in_0_valid & chosen); // @[SwitchAllocator.scala 44:45]
  assign io_out_0_bits_vc_sel_0_0 = io_in_0_bits_vc_sel_0_0; // @[SwitchAllocator.scala 45:20]
  assign io_out_0_bits_vc_sel_0_1 = io_in_0_bits_vc_sel_0_1; // @[SwitchAllocator.scala 45:20]
  assign io_out_0_bits_vc_sel_0_2 = io_in_0_bits_vc_sel_0_2; // @[SwitchAllocator.scala 45:20]
  assign io_chosen_oh_0 = |(io_in_0_valid & lock_0) ? lock_0 : choices_0; // @[SwitchAllocator.scala 42:21]
  always @(posedge clock) begin
    if (reset) begin // @[SwitchAllocator.scala 24:38]
      lock_0 <= 1'h0; // @[SwitchAllocator.scala 24:38]
    end else if (io_out_0_valid) begin // @[SwitchAllocator.scala 52:29]
      lock_0 <= chosen & ~io_in_0_bits_tail; // @[SwitchAllocator.scala 53:15]
    end
    mask <= _GEN_4[0]; // @[SwitchAllocator.scala 27:{21,21}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lock_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  mask = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SwitchAllocator(
  input   clock,
  input   reset,
  output  io_req_0_0_ready,
  input   io_req_0_0_valid,
  input   io_req_0_0_bits_vc_sel_0_0,
  input   io_req_0_0_bits_vc_sel_0_1,
  input   io_req_0_0_bits_vc_sel_0_2,
  input   io_req_0_0_bits_tail,
  output  io_credit_alloc_0_0_alloc,
  output  io_credit_alloc_0_1_alloc,
  output  io_credit_alloc_0_2_alloc,
  output  io_switch_sel_0_0_0_0
);
  wire  arbs_0_clock; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_reset; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_0_ready; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_0_valid; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_0_bits_vc_sel_0_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_0_bits_vc_sel_0_1; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_0_bits_vc_sel_0_2; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_0_bits_tail; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_out_0_valid; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_out_0_bits_vc_sel_0_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_out_0_bits_vc_sel_0_1; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_out_0_bits_vc_sel_0_2; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_chosen_oh_0; // @[SwitchAllocator.scala 83:45]
  SwitchArbiter arbs_0 ( // @[SwitchAllocator.scala 83:45]
    .clock(arbs_0_clock),
    .reset(arbs_0_reset),
    .io_in_0_ready(arbs_0_io_in_0_ready),
    .io_in_0_valid(arbs_0_io_in_0_valid),
    .io_in_0_bits_vc_sel_0_0(arbs_0_io_in_0_bits_vc_sel_0_0),
    .io_in_0_bits_vc_sel_0_1(arbs_0_io_in_0_bits_vc_sel_0_1),
    .io_in_0_bits_vc_sel_0_2(arbs_0_io_in_0_bits_vc_sel_0_2),
    .io_in_0_bits_tail(arbs_0_io_in_0_bits_tail),
    .io_out_0_valid(arbs_0_io_out_0_valid),
    .io_out_0_bits_vc_sel_0_0(arbs_0_io_out_0_bits_vc_sel_0_0),
    .io_out_0_bits_vc_sel_0_1(arbs_0_io_out_0_bits_vc_sel_0_1),
    .io_out_0_bits_vc_sel_0_2(arbs_0_io_out_0_bits_vc_sel_0_2),
    .io_chosen_oh_0(arbs_0_io_chosen_oh_0)
  );
  assign io_req_0_0_ready = arbs_0_io_in_0_ready & arbs_0_io_in_0_valid; // @[Decoupled.scala 51:35]
  assign io_credit_alloc_0_0_alloc = arbs_0_io_out_0_valid & arbs_0_io_out_0_bits_vc_sel_0_0; // @[SwitchAllocator.scala 120:33]
  assign io_credit_alloc_0_1_alloc = arbs_0_io_out_0_valid & arbs_0_io_out_0_bits_vc_sel_0_1; // @[SwitchAllocator.scala 120:33]
  assign io_credit_alloc_0_2_alloc = arbs_0_io_out_0_valid & arbs_0_io_out_0_bits_vc_sel_0_2; // @[SwitchAllocator.scala 120:33]
  assign io_switch_sel_0_0_0_0 = arbs_0_io_in_0_valid & arbs_0_io_chosen_oh_0 & arbs_0_io_out_0_valid; // @[SwitchAllocator.scala 108:97]
  assign arbs_0_clock = clock;
  assign arbs_0_reset = reset;
  assign arbs_0_io_in_0_valid = io_req_0_0_valid & (io_req_0_0_bits_vc_sel_0_0 | io_req_0_0_bits_vc_sel_0_1 |
    io_req_0_0_bits_vc_sel_0_2); // @[SwitchAllocator.scala 95:37]
  assign arbs_0_io_in_0_bits_vc_sel_0_0 = io_req_0_0_bits_vc_sel_0_0; // @[SwitchAllocator.scala 96:25]
  assign arbs_0_io_in_0_bits_vc_sel_0_1 = io_req_0_0_bits_vc_sel_0_1; // @[SwitchAllocator.scala 96:25]
  assign arbs_0_io_in_0_bits_vc_sel_0_2 = io_req_0_0_bits_vc_sel_0_2; // @[SwitchAllocator.scala 96:25]
  assign arbs_0_io_in_0_bits_tail = io_req_0_0_bits_tail; // @[SwitchAllocator.scala 96:25]
endmodule
module RotatingSingleVCAllocator(
  input   clock,
  input   reset,
  output  io_req_0_ready,
  input   io_req_0_valid,
  input   io_req_0_bits_vc_sel_0_0,
  input   io_req_0_bits_vc_sel_0_1,
  input   io_req_0_bits_vc_sel_0_2,
  output  io_resp_0_vc_sel_0_0,
  output  io_resp_0_vc_sel_0_1,
  output  io_resp_0_vc_sel_0_2,
  input   io_channel_status_0_0_occupied,
  input   io_channel_status_0_1_occupied,
  input   io_channel_status_0_2_occupied,
  output  io_out_allocs_0_0_alloc,
  output  io_out_allocs_0_1_alloc,
  output  io_out_allocs_0_2_alloc
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  mask; // @[SingleVCAllocator.scala 16:21]
  wire  in_arb_reqs_0_0_0 = io_req_0_bits_vc_sel_0_0 & ~io_channel_status_0_0_occupied; // @[SingleVCAllocator.scala 28:61]
  wire  in_arb_reqs_0_0_1 = io_req_0_bits_vc_sel_0_1 & ~io_channel_status_0_1_occupied; // @[SingleVCAllocator.scala 28:61]
  wire  in_arb_reqs_0_0_2 = io_req_0_bits_vc_sel_0_2 & ~io_channel_status_0_2_occupied; // @[SingleVCAllocator.scala 28:61]
  wire  _in_arb_vals_0_T_1 = in_arb_reqs_0_0_0 | in_arb_reqs_0_0_1 | in_arb_reqs_0_0_2; // @[package.scala 73:59]
  wire  in_arb_vals_0 = io_req_0_valid & _in_arb_vals_0_T_1; // @[SingleVCAllocator.scala 32:39]
  wire  _in_arb_filter_T_1 = in_arb_vals_0 & ~mask; // @[SingleVCAllocator.scala 19:84]
  wire [1:0] _in_arb_filter_T_2 = {in_arb_vals_0,_in_arb_filter_T_1}; // @[Cat.scala 33:92]
  wire [1:0] _in_arb_filter_T_5 = _in_arb_filter_T_2[1] ? 2'h2 : 2'h0; // @[Mux.scala 47:70]
  wire [1:0] in_arb_filter = _in_arb_filter_T_2[0] ? 2'h1 : _in_arb_filter_T_5; // @[Mux.scala 47:70]
  wire  _GEN_0 = in_arb_vals_0 | mask; // @[SingleVCAllocator.scala 21:26 22:10 16:21]
  wire  _in_alloc_T = io_req_0_ready & io_req_0_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _in_alloc_T_1 = {in_arb_reqs_0_0_2,in_arb_reqs_0_0_1,in_arb_reqs_0_0_0}; // @[ISLIP.scala 33:18]
  reg [2:0] in_alloc_mask; // @[ISLIP.scala 17:25]
  wire [2:0] _in_alloc_full_T = ~in_alloc_mask; // @[ISLIP.scala 18:31]
  wire [2:0] _in_alloc_full_T_1 = _in_alloc_T_1 & _in_alloc_full_T; // @[ISLIP.scala 18:29]
  wire [5:0] in_alloc_full = {in_arb_reqs_0_0_2,in_arb_reqs_0_0_1,in_arb_reqs_0_0_0,_in_alloc_full_T_1}; // @[Cat.scala 33:92]
  wire [5:0] _in_alloc_oh_T_6 = in_alloc_full[5] ? 6'h20 : 6'h0; // @[Mux.scala 47:70]
  wire [5:0] _in_alloc_oh_T_7 = in_alloc_full[4] ? 6'h10 : _in_alloc_oh_T_6; // @[Mux.scala 47:70]
  wire [5:0] _in_alloc_oh_T_8 = in_alloc_full[3] ? 6'h8 : _in_alloc_oh_T_7; // @[Mux.scala 47:70]
  wire [5:0] _in_alloc_oh_T_9 = in_alloc_full[2] ? 6'h4 : _in_alloc_oh_T_8; // @[Mux.scala 47:70]
  wire [5:0] _in_alloc_oh_T_10 = in_alloc_full[1] ? 6'h2 : _in_alloc_oh_T_9; // @[Mux.scala 47:70]
  wire [5:0] in_alloc_oh = in_alloc_full[0] ? 6'h1 : _in_alloc_oh_T_10; // @[Mux.scala 47:70]
  wire [2:0] in_alloc_sel = in_alloc_oh[2:0] | in_alloc_oh[5:3]; // @[ISLIP.scala 20:28]
  wire [2:0] _in_alloc_mask_T_6 = in_alloc_sel[2] ? 3'h7 : 3'h0; // @[Mux.scala 101:16]
  wire [2:0] _T = {io_resp_0_vc_sel_0_2,io_resp_0_vc_sel_0_1,io_resp_0_vc_sel_0_0}; // @[SingleVCAllocator.scala 53:39]
  wire [1:0] _T_4 = _T[1] + _T[2]; // @[Bitwise.scala 51:90]
  wire [1:0] _GEN_2 = {{1'd0}, _T[0]}; // @[Bitwise.scala 51:90]
  wire [2:0] _T_6 = _GEN_2 + _T_4; // @[Bitwise.scala 51:90]
  assign io_req_0_ready = in_arb_filter[0] | in_arb_filter[1]; // @[SingleVCAllocator.scala 20:57]
  assign io_resp_0_vc_sel_0_0 = in_arb_vals_0 & in_alloc_sel[0]; // @[SingleVCAllocator.scala 41:18]
  assign io_resp_0_vc_sel_0_1 = in_arb_vals_0 & in_alloc_sel[1]; // @[SingleVCAllocator.scala 41:18]
  assign io_resp_0_vc_sel_0_2 = in_arb_vals_0 & in_alloc_sel[2]; // @[SingleVCAllocator.scala 41:18]
  assign io_out_allocs_0_0_alloc = in_arb_vals_0 & in_alloc_sel[0]; // @[SingleVCAllocator.scala 41:18]
  assign io_out_allocs_0_1_alloc = in_arb_vals_0 & in_alloc_sel[1]; // @[SingleVCAllocator.scala 41:18]
  assign io_out_allocs_0_2_alloc = in_arb_vals_0 & in_alloc_sel[2]; // @[SingleVCAllocator.scala 41:18]
  always @(posedge clock) begin
    if (reset) begin // @[SingleVCAllocator.scala 16:21]
      mask <= 1'h0; // @[SingleVCAllocator.scala 16:21]
    end else begin
      mask <= _GEN_0;
    end
    if (reset) begin // @[ISLIP.scala 17:25]
      in_alloc_mask <= 3'h0; // @[ISLIP.scala 17:25]
    end else if (_in_alloc_T) begin // @[ISLIP.scala 21:19]
      if (in_alloc_sel[0]) begin // @[Mux.scala 101:16]
        in_alloc_mask <= 3'h1;
      end else if (in_alloc_sel[1]) begin // @[Mux.scala 101:16]
        in_alloc_mask <= 3'h3;
      end else begin
        in_alloc_mask <= _in_alloc_mask_T_6;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(_T_6[1:0] <= 2'h1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at SingleVCAllocator.scala:53 assert(PopCount(io.resp(i).vc_sel.asUInt) <= 1.U)\n"); // @[SingleVCAllocator.scala 53:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mask = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  in_alloc_mask = _RAND_1[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(_T_6[1:0] <= 2'h1); // @[SingleVCAllocator.scala 53:11]
    end
  end
endmodule
module Router(
  input         clock,
  input         reset,
  output        auto_ingress_nodes_in_flit_ready,
  input         auto_ingress_nodes_in_flit_valid,
  input         auto_ingress_nodes_in_flit_bits_head,
  input         auto_ingress_nodes_in_flit_bits_tail,
  input  [63:0] auto_ingress_nodes_in_flit_bits_payload,
  input         auto_ingress_nodes_in_flit_bits_egress_id,
  output        auto_source_nodes_out_flit_0_valid,
  output        auto_source_nodes_out_flit_0_bits_head,
  output        auto_source_nodes_out_flit_0_bits_tail,
  output [63:0] auto_source_nodes_out_flit_0_bits_payload,
  output        auto_source_nodes_out_flit_0_bits_flow_ingress_node,
  output        auto_source_nodes_out_flit_0_bits_flow_egress_node,
  output [1:0]  auto_source_nodes_out_flit_0_bits_virt_channel_id,
  input  [2:0]  auto_source_nodes_out_credit_return,
  input  [2:0]  auto_source_nodes_out_vc_free
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  ingress_unit_0_from_0_clock; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_reset; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_router_req_valid; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_vcalloc_req_ready; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_vcalloc_req_valid; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_0; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_1; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_2; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_vcalloc_resp_vc_sel_0_0; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_vcalloc_resp_vc_sel_0_1; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_vcalloc_resp_vc_sel_0_2; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_out_credit_available_0_0; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_out_credit_available_0_1; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_out_credit_available_0_2; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_salloc_req_0_ready; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_salloc_req_0_valid; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_0; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_1; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_2; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_salloc_req_0_bits_tail; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_out_0_valid; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_out_0_bits_flit_head; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_out_0_bits_flit_tail; // @[Router.scala 116:13]
  wire [63:0] ingress_unit_0_from_0_io_out_0_bits_flit_payload; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_out_0_bits_flit_flow_ingress_node; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_out_0_bits_flit_flow_egress_node; // @[Router.scala 116:13]
  wire [1:0] ingress_unit_0_from_0_io_out_0_bits_out_virt_channel; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_in_ready; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_in_valid; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_in_bits_head; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_in_bits_tail; // @[Router.scala 116:13]
  wire [63:0] ingress_unit_0_from_0_io_in_bits_payload; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_in_bits_egress_id; // @[Router.scala 116:13]
  wire  output_unit_0_to_1_clock; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_reset; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_in_0_valid; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_in_0_bits_head; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_in_0_bits_tail; // @[Router.scala 122:13]
  wire [63:0] output_unit_0_to_1_io_in_0_bits_payload; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_in_0_bits_flow_ingress_node; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_in_0_bits_flow_egress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_0_to_1_io_in_0_bits_virt_channel_id; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_credit_available_0; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_credit_available_1; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_credit_available_2; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_channel_status_0_occupied; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_channel_status_1_occupied; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_channel_status_2_occupied; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_allocs_0_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_allocs_1_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_allocs_2_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_credit_alloc_0_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_credit_alloc_1_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_credit_alloc_2_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_out_flit_0_valid; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_out_flit_0_bits_head; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_out_flit_0_bits_tail; // @[Router.scala 122:13]
  wire [63:0] output_unit_0_to_1_io_out_flit_0_bits_payload; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_out_flit_0_bits_flow_ingress_node; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_out_flit_0_bits_flow_egress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_0_to_1_io_out_flit_0_bits_virt_channel_id; // @[Router.scala 122:13]
  wire [2:0] output_unit_0_to_1_io_out_credit_return; // @[Router.scala 122:13]
  wire [2:0] output_unit_0_to_1_io_out_vc_free; // @[Router.scala 122:13]
  wire  switch_clock; // @[Router.scala 129:24]
  wire  switch_reset; // @[Router.scala 129:24]
  wire  switch_io_in_0_0_valid; // @[Router.scala 129:24]
  wire  switch_io_in_0_0_bits_flit_head; // @[Router.scala 129:24]
  wire  switch_io_in_0_0_bits_flit_tail; // @[Router.scala 129:24]
  wire [63:0] switch_io_in_0_0_bits_flit_payload; // @[Router.scala 129:24]
  wire  switch_io_in_0_0_bits_flit_flow_ingress_node; // @[Router.scala 129:24]
  wire  switch_io_in_0_0_bits_flit_flow_egress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_0_0_bits_out_virt_channel; // @[Router.scala 129:24]
  wire  switch_io_out_0_0_valid; // @[Router.scala 129:24]
  wire  switch_io_out_0_0_bits_head; // @[Router.scala 129:24]
  wire  switch_io_out_0_0_bits_tail; // @[Router.scala 129:24]
  wire [63:0] switch_io_out_0_0_bits_payload; // @[Router.scala 129:24]
  wire  switch_io_out_0_0_bits_flow_ingress_node; // @[Router.scala 129:24]
  wire  switch_io_out_0_0_bits_flow_egress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_out_0_0_bits_virt_channel_id; // @[Router.scala 129:24]
  wire  switch_io_sel_0_0_0_0; // @[Router.scala 129:24]
  wire  switch_allocator_clock; // @[Router.scala 130:34]
  wire  switch_allocator_reset; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_ready; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_valid; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_0_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_0_1; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_0_2; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_tail; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_0_0_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_0_1_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_0_2_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_0_0_0_0; // @[Router.scala 130:34]
  wire  vc_allocator_clock; // @[Router.scala 131:30]
  wire  vc_allocator_reset; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_ready; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_valid; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_0_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_0_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_0_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_0_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_0_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_0_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_0_0_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_0_1_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_0_2_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_0_0_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_0_1_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_0_2_alloc; // @[Router.scala 131:30]
  wire [19:0] plusarg_reader_out; // @[PlusArg.scala 80:11]
  reg  switch_io_sel_REG_0_0_0_0; // @[Router.scala 176:14]
  reg [63:0] debug_tsc; // @[Router.scala 193:28]
  wire [63:0] _debug_tsc_T_1 = debug_tsc + 64'h1; // @[Router.scala 194:28]
  reg [63:0] debug_sample; // @[Router.scala 195:31]
  wire [63:0] _debug_sample_T_1 = debug_sample + 64'h1; // @[Router.scala 196:34]
  wire [19:0] _T_1 = plusarg_reader_out - 20'h1; // @[Router.scala 198:40]
  wire [63:0] _GEN_2 = {{44'd0}, _T_1}; // @[Router.scala 198:24]
  wire  _T_2 = debug_sample == _GEN_2; // @[Router.scala 198:24]
  wire  bundleIn_0_flit_ready = ingress_unit_0_from_0_io_in_ready; // @[Nodes.scala 1215:84 Router.scala 142:68]
  wire  _T_3 = bundleIn_0_flit_ready & auto_ingress_nodes_in_flit_valid; // @[Decoupled.scala 51:35]
  reg [63:0] util_ctr; // @[Router.scala 201:29]
  reg  fired; // @[Router.scala 202:26]
  wire [63:0] _GEN_3 = {{63'd0}, _T_3}; // @[Router.scala 203:28]
  wire [63:0] _util_ctr_T_1 = util_ctr + _GEN_3; // @[Router.scala 203:28]
  wire  _T_9 = plusarg_reader_out != 20'h0 & _T_2 & fired; // @[Router.scala 205:71]
  wire  fires_count = vc_allocator_io_req_0_ready & vc_allocator_io_req_0_valid; // @[Decoupled.scala 51:35]
  IngressUnit ingress_unit_0_from_0 ( // @[Router.scala 116:13]
    .clock(ingress_unit_0_from_0_clock),
    .reset(ingress_unit_0_from_0_reset),
    .io_router_req_valid(ingress_unit_0_from_0_io_router_req_valid),
    .io_vcalloc_req_ready(ingress_unit_0_from_0_io_vcalloc_req_ready),
    .io_vcalloc_req_valid(ingress_unit_0_from_0_io_vcalloc_req_valid),
    .io_vcalloc_req_bits_vc_sel_0_0(ingress_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_0),
    .io_vcalloc_req_bits_vc_sel_0_1(ingress_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_1),
    .io_vcalloc_req_bits_vc_sel_0_2(ingress_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_2),
    .io_vcalloc_resp_vc_sel_0_0(ingress_unit_0_from_0_io_vcalloc_resp_vc_sel_0_0),
    .io_vcalloc_resp_vc_sel_0_1(ingress_unit_0_from_0_io_vcalloc_resp_vc_sel_0_1),
    .io_vcalloc_resp_vc_sel_0_2(ingress_unit_0_from_0_io_vcalloc_resp_vc_sel_0_2),
    .io_out_credit_available_0_0(ingress_unit_0_from_0_io_out_credit_available_0_0),
    .io_out_credit_available_0_1(ingress_unit_0_from_0_io_out_credit_available_0_1),
    .io_out_credit_available_0_2(ingress_unit_0_from_0_io_out_credit_available_0_2),
    .io_salloc_req_0_ready(ingress_unit_0_from_0_io_salloc_req_0_ready),
    .io_salloc_req_0_valid(ingress_unit_0_from_0_io_salloc_req_0_valid),
    .io_salloc_req_0_bits_vc_sel_0_0(ingress_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_0),
    .io_salloc_req_0_bits_vc_sel_0_1(ingress_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_1),
    .io_salloc_req_0_bits_vc_sel_0_2(ingress_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_2),
    .io_salloc_req_0_bits_tail(ingress_unit_0_from_0_io_salloc_req_0_bits_tail),
    .io_out_0_valid(ingress_unit_0_from_0_io_out_0_valid),
    .io_out_0_bits_flit_head(ingress_unit_0_from_0_io_out_0_bits_flit_head),
    .io_out_0_bits_flit_tail(ingress_unit_0_from_0_io_out_0_bits_flit_tail),
    .io_out_0_bits_flit_payload(ingress_unit_0_from_0_io_out_0_bits_flit_payload),
    .io_out_0_bits_flit_flow_ingress_node(ingress_unit_0_from_0_io_out_0_bits_flit_flow_ingress_node),
    .io_out_0_bits_flit_flow_egress_node(ingress_unit_0_from_0_io_out_0_bits_flit_flow_egress_node),
    .io_out_0_bits_out_virt_channel(ingress_unit_0_from_0_io_out_0_bits_out_virt_channel),
    .io_in_ready(ingress_unit_0_from_0_io_in_ready),
    .io_in_valid(ingress_unit_0_from_0_io_in_valid),
    .io_in_bits_head(ingress_unit_0_from_0_io_in_bits_head),
    .io_in_bits_tail(ingress_unit_0_from_0_io_in_bits_tail),
    .io_in_bits_payload(ingress_unit_0_from_0_io_in_bits_payload),
    .io_in_bits_egress_id(ingress_unit_0_from_0_io_in_bits_egress_id)
  );
  OutputUnit output_unit_0_to_1 ( // @[Router.scala 122:13]
    .clock(output_unit_0_to_1_clock),
    .reset(output_unit_0_to_1_reset),
    .io_in_0_valid(output_unit_0_to_1_io_in_0_valid),
    .io_in_0_bits_head(output_unit_0_to_1_io_in_0_bits_head),
    .io_in_0_bits_tail(output_unit_0_to_1_io_in_0_bits_tail),
    .io_in_0_bits_payload(output_unit_0_to_1_io_in_0_bits_payload),
    .io_in_0_bits_flow_ingress_node(output_unit_0_to_1_io_in_0_bits_flow_ingress_node),
    .io_in_0_bits_flow_egress_node(output_unit_0_to_1_io_in_0_bits_flow_egress_node),
    .io_in_0_bits_virt_channel_id(output_unit_0_to_1_io_in_0_bits_virt_channel_id),
    .io_credit_available_0(output_unit_0_to_1_io_credit_available_0),
    .io_credit_available_1(output_unit_0_to_1_io_credit_available_1),
    .io_credit_available_2(output_unit_0_to_1_io_credit_available_2),
    .io_channel_status_0_occupied(output_unit_0_to_1_io_channel_status_0_occupied),
    .io_channel_status_1_occupied(output_unit_0_to_1_io_channel_status_1_occupied),
    .io_channel_status_2_occupied(output_unit_0_to_1_io_channel_status_2_occupied),
    .io_allocs_0_alloc(output_unit_0_to_1_io_allocs_0_alloc),
    .io_allocs_1_alloc(output_unit_0_to_1_io_allocs_1_alloc),
    .io_allocs_2_alloc(output_unit_0_to_1_io_allocs_2_alloc),
    .io_credit_alloc_0_alloc(output_unit_0_to_1_io_credit_alloc_0_alloc),
    .io_credit_alloc_1_alloc(output_unit_0_to_1_io_credit_alloc_1_alloc),
    .io_credit_alloc_2_alloc(output_unit_0_to_1_io_credit_alloc_2_alloc),
    .io_out_flit_0_valid(output_unit_0_to_1_io_out_flit_0_valid),
    .io_out_flit_0_bits_head(output_unit_0_to_1_io_out_flit_0_bits_head),
    .io_out_flit_0_bits_tail(output_unit_0_to_1_io_out_flit_0_bits_tail),
    .io_out_flit_0_bits_payload(output_unit_0_to_1_io_out_flit_0_bits_payload),
    .io_out_flit_0_bits_flow_ingress_node(output_unit_0_to_1_io_out_flit_0_bits_flow_ingress_node),
    .io_out_flit_0_bits_flow_egress_node(output_unit_0_to_1_io_out_flit_0_bits_flow_egress_node),
    .io_out_flit_0_bits_virt_channel_id(output_unit_0_to_1_io_out_flit_0_bits_virt_channel_id),
    .io_out_credit_return(output_unit_0_to_1_io_out_credit_return),
    .io_out_vc_free(output_unit_0_to_1_io_out_vc_free)
  );
  Switch switch ( // @[Router.scala 129:24]
    .clock(switch_clock),
    .reset(switch_reset),
    .io_in_0_0_valid(switch_io_in_0_0_valid),
    .io_in_0_0_bits_flit_head(switch_io_in_0_0_bits_flit_head),
    .io_in_0_0_bits_flit_tail(switch_io_in_0_0_bits_flit_tail),
    .io_in_0_0_bits_flit_payload(switch_io_in_0_0_bits_flit_payload),
    .io_in_0_0_bits_flit_flow_ingress_node(switch_io_in_0_0_bits_flit_flow_ingress_node),
    .io_in_0_0_bits_flit_flow_egress_node(switch_io_in_0_0_bits_flit_flow_egress_node),
    .io_in_0_0_bits_out_virt_channel(switch_io_in_0_0_bits_out_virt_channel),
    .io_out_0_0_valid(switch_io_out_0_0_valid),
    .io_out_0_0_bits_head(switch_io_out_0_0_bits_head),
    .io_out_0_0_bits_tail(switch_io_out_0_0_bits_tail),
    .io_out_0_0_bits_payload(switch_io_out_0_0_bits_payload),
    .io_out_0_0_bits_flow_ingress_node(switch_io_out_0_0_bits_flow_ingress_node),
    .io_out_0_0_bits_flow_egress_node(switch_io_out_0_0_bits_flow_egress_node),
    .io_out_0_0_bits_virt_channel_id(switch_io_out_0_0_bits_virt_channel_id),
    .io_sel_0_0_0_0(switch_io_sel_0_0_0_0)
  );
  SwitchAllocator switch_allocator ( // @[Router.scala 130:34]
    .clock(switch_allocator_clock),
    .reset(switch_allocator_reset),
    .io_req_0_0_ready(switch_allocator_io_req_0_0_ready),
    .io_req_0_0_valid(switch_allocator_io_req_0_0_valid),
    .io_req_0_0_bits_vc_sel_0_0(switch_allocator_io_req_0_0_bits_vc_sel_0_0),
    .io_req_0_0_bits_vc_sel_0_1(switch_allocator_io_req_0_0_bits_vc_sel_0_1),
    .io_req_0_0_bits_vc_sel_0_2(switch_allocator_io_req_0_0_bits_vc_sel_0_2),
    .io_req_0_0_bits_tail(switch_allocator_io_req_0_0_bits_tail),
    .io_credit_alloc_0_0_alloc(switch_allocator_io_credit_alloc_0_0_alloc),
    .io_credit_alloc_0_1_alloc(switch_allocator_io_credit_alloc_0_1_alloc),
    .io_credit_alloc_0_2_alloc(switch_allocator_io_credit_alloc_0_2_alloc),
    .io_switch_sel_0_0_0_0(switch_allocator_io_switch_sel_0_0_0_0)
  );
  RotatingSingleVCAllocator vc_allocator ( // @[Router.scala 131:30]
    .clock(vc_allocator_clock),
    .reset(vc_allocator_reset),
    .io_req_0_ready(vc_allocator_io_req_0_ready),
    .io_req_0_valid(vc_allocator_io_req_0_valid),
    .io_req_0_bits_vc_sel_0_0(vc_allocator_io_req_0_bits_vc_sel_0_0),
    .io_req_0_bits_vc_sel_0_1(vc_allocator_io_req_0_bits_vc_sel_0_1),
    .io_req_0_bits_vc_sel_0_2(vc_allocator_io_req_0_bits_vc_sel_0_2),
    .io_resp_0_vc_sel_0_0(vc_allocator_io_resp_0_vc_sel_0_0),
    .io_resp_0_vc_sel_0_1(vc_allocator_io_resp_0_vc_sel_0_1),
    .io_resp_0_vc_sel_0_2(vc_allocator_io_resp_0_vc_sel_0_2),
    .io_channel_status_0_0_occupied(vc_allocator_io_channel_status_0_0_occupied),
    .io_channel_status_0_1_occupied(vc_allocator_io_channel_status_0_1_occupied),
    .io_channel_status_0_2_occupied(vc_allocator_io_channel_status_0_2_occupied),
    .io_out_allocs_0_0_alloc(vc_allocator_io_out_allocs_0_0_alloc),
    .io_out_allocs_0_1_alloc(vc_allocator_io_out_allocs_0_1_alloc),
    .io_out_allocs_0_2_alloc(vc_allocator_io_out_allocs_0_2_alloc)
  );
  plusarg_reader #(.FORMAT("noc_util_sample_rate=%d"), .DEFAULT(0), .WIDTH(20)) plusarg_reader ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_out)
  );
  assign auto_ingress_nodes_in_flit_ready = ingress_unit_0_from_0_io_in_ready; // @[Nodes.scala 1215:84 Router.scala 142:68]
  assign auto_source_nodes_out_flit_0_valid = output_unit_0_to_1_io_out_flit_0_valid; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_flit_0_bits_head = output_unit_0_to_1_io_out_flit_0_bits_head; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_flit_0_bits_tail = output_unit_0_to_1_io_out_flit_0_bits_tail; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_flit_0_bits_payload = output_unit_0_to_1_io_out_flit_0_bits_payload; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_flit_0_bits_flow_ingress_node = output_unit_0_to_1_io_out_flit_0_bits_flow_ingress_node; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_flit_0_bits_flow_egress_node = output_unit_0_to_1_io_out_flit_0_bits_flow_egress_node; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_flit_0_bits_virt_channel_id = output_unit_0_to_1_io_out_flit_0_bits_virt_channel_id; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign ingress_unit_0_from_0_clock = clock;
  assign ingress_unit_0_from_0_reset = reset;
  assign ingress_unit_0_from_0_io_vcalloc_req_ready = vc_allocator_io_req_0_ready; // @[Router.scala 151:23]
  assign ingress_unit_0_from_0_io_vcalloc_resp_vc_sel_0_0 = vc_allocator_io_resp_0_vc_sel_0_0; // @[Router.scala 153:39]
  assign ingress_unit_0_from_0_io_vcalloc_resp_vc_sel_0_1 = vc_allocator_io_resp_0_vc_sel_0_1; // @[Router.scala 153:39]
  assign ingress_unit_0_from_0_io_vcalloc_resp_vc_sel_0_2 = vc_allocator_io_resp_0_vc_sel_0_2; // @[Router.scala 153:39]
  assign ingress_unit_0_from_0_io_out_credit_available_0_0 = output_unit_0_to_1_io_credit_available_0; // @[Router.scala 162:42]
  assign ingress_unit_0_from_0_io_out_credit_available_0_1 = output_unit_0_to_1_io_credit_available_1; // @[Router.scala 162:42]
  assign ingress_unit_0_from_0_io_out_credit_available_0_2 = output_unit_0_to_1_io_credit_available_2; // @[Router.scala 162:42]
  assign ingress_unit_0_from_0_io_salloc_req_0_ready = switch_allocator_io_req_0_0_ready; // @[Router.scala 165:23]
  assign ingress_unit_0_from_0_io_in_valid = auto_ingress_nodes_in_flit_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign ingress_unit_0_from_0_io_in_bits_head = auto_ingress_nodes_in_flit_bits_head; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign ingress_unit_0_from_0_io_in_bits_tail = auto_ingress_nodes_in_flit_bits_tail; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign ingress_unit_0_from_0_io_in_bits_payload = auto_ingress_nodes_in_flit_bits_payload; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign ingress_unit_0_from_0_io_in_bits_egress_id = auto_ingress_nodes_in_flit_bits_egress_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign output_unit_0_to_1_clock = clock;
  assign output_unit_0_to_1_reset = reset;
  assign output_unit_0_to_1_io_in_0_valid = switch_io_out_0_0_valid; // @[Router.scala 172:29]
  assign output_unit_0_to_1_io_in_0_bits_head = switch_io_out_0_0_bits_head; // @[Router.scala 172:29]
  assign output_unit_0_to_1_io_in_0_bits_tail = switch_io_out_0_0_bits_tail; // @[Router.scala 172:29]
  assign output_unit_0_to_1_io_in_0_bits_payload = switch_io_out_0_0_bits_payload; // @[Router.scala 172:29]
  assign output_unit_0_to_1_io_in_0_bits_flow_ingress_node = switch_io_out_0_0_bits_flow_ingress_node; // @[Router.scala 172:29]
  assign output_unit_0_to_1_io_in_0_bits_flow_egress_node = switch_io_out_0_0_bits_flow_egress_node; // @[Router.scala 172:29]
  assign output_unit_0_to_1_io_in_0_bits_virt_channel_id = switch_io_out_0_0_bits_virt_channel_id; // @[Router.scala 172:29]
  assign output_unit_0_to_1_io_allocs_0_alloc = vc_allocator_io_out_allocs_0_0_alloc; // @[Router.scala 157:33]
  assign output_unit_0_to_1_io_allocs_1_alloc = vc_allocator_io_out_allocs_0_1_alloc; // @[Router.scala 157:33]
  assign output_unit_0_to_1_io_allocs_2_alloc = vc_allocator_io_out_allocs_0_2_alloc; // @[Router.scala 157:33]
  assign output_unit_0_to_1_io_credit_alloc_0_alloc = switch_allocator_io_credit_alloc_0_0_alloc; // @[Router.scala 167:39]
  assign output_unit_0_to_1_io_credit_alloc_1_alloc = switch_allocator_io_credit_alloc_0_1_alloc; // @[Router.scala 167:39]
  assign output_unit_0_to_1_io_credit_alloc_2_alloc = switch_allocator_io_credit_alloc_0_2_alloc; // @[Router.scala 167:39]
  assign output_unit_0_to_1_io_out_credit_return = auto_source_nodes_out_credit_return; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign output_unit_0_to_1_io_out_vc_free = auto_source_nodes_out_vc_free; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign switch_clock = clock;
  assign switch_reset = reset;
  assign switch_io_in_0_0_valid = ingress_unit_0_from_0_io_out_0_valid; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_head = ingress_unit_0_from_0_io_out_0_bits_flit_head; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_tail = ingress_unit_0_from_0_io_out_0_bits_flit_tail; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_payload = ingress_unit_0_from_0_io_out_0_bits_flit_payload; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_flow_ingress_node = ingress_unit_0_from_0_io_out_0_bits_flit_flow_ingress_node; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_flow_egress_node = ingress_unit_0_from_0_io_out_0_bits_flit_flow_egress_node; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_out_virt_channel = ingress_unit_0_from_0_io_out_0_bits_out_virt_channel; // @[Router.scala 170:23]
  assign switch_io_sel_0_0_0_0 = switch_io_sel_REG_0_0_0_0; // @[Router.scala 173:19]
  assign switch_allocator_clock = clock;
  assign switch_allocator_reset = reset;
  assign switch_allocator_io_req_0_0_valid = ingress_unit_0_from_0_io_salloc_req_0_valid; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_0_0 = ingress_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_0_1 = ingress_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_1; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_0_2 = ingress_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_2; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_tail = ingress_unit_0_from_0_io_salloc_req_0_bits_tail; // @[Router.scala 165:23]
  assign vc_allocator_clock = clock;
  assign vc_allocator_reset = reset;
  assign vc_allocator_io_req_0_valid = ingress_unit_0_from_0_io_vcalloc_req_valid; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_0_0 = ingress_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_0_1 = ingress_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_1; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_0_2 = ingress_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_2; // @[Router.scala 151:23]
  assign vc_allocator_io_channel_status_0_0_occupied = output_unit_0_to_1_io_channel_status_0_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_0_1_occupied = output_unit_0_to_1_io_channel_status_1_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_0_2_occupied = output_unit_0_to_1_io_channel_status_2_occupied; // @[Router.scala 159:23]
  always @(posedge clock) begin
    switch_io_sel_REG_0_0_0_0 <= switch_allocator_io_switch_sel_0_0_0_0; // @[Router.scala 176:14]
    if (reset) begin // @[Router.scala 193:28]
      debug_tsc <= 64'h0; // @[Router.scala 193:28]
    end else begin
      debug_tsc <= _debug_tsc_T_1; // @[Router.scala 194:15]
    end
    if (reset) begin // @[Router.scala 195:31]
      debug_sample <= 64'h0; // @[Router.scala 195:31]
    end else if (debug_sample == _GEN_2) begin // @[Router.scala 198:47]
      debug_sample <= 64'h0; // @[Router.scala 198:62]
    end else begin
      debug_sample <= _debug_sample_T_1; // @[Router.scala 196:18]
    end
    if (reset) begin // @[Router.scala 201:29]
      util_ctr <= 64'h0; // @[Router.scala 201:29]
    end else begin
      util_ctr <= _util_ctr_T_1; // @[Router.scala 203:16]
    end
    if (reset) begin // @[Router.scala 202:26]
      fired <= 1'h0; // @[Router.scala 202:26]
    end else if (plusarg_reader_out != 20'h0 & _T_2 & fired) begin // @[Router.scala 205:81]
      fired <= _T_3; // @[Router.scala 208:15]
    end else begin
      fired <= fired | _T_3; // @[Router.scala 204:13]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9 & ~reset) begin
          $fwrite(32'h80000002,"nocsample %d i0 0 %d\n",debug_tsc,util_ctr); // @[Router.scala 207:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  switch_io_sel_REG_0_0_0_0 = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  debug_tsc = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  debug_sample = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  util_ctr = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  fired = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ClockSinkDomain(
  output        auto_routers_ingress_nodes_in_flit_ready,
  input         auto_routers_ingress_nodes_in_flit_valid,
  input         auto_routers_ingress_nodes_in_flit_bits_head,
  input         auto_routers_ingress_nodes_in_flit_bits_tail,
  input  [63:0] auto_routers_ingress_nodes_in_flit_bits_payload,
  input         auto_routers_ingress_nodes_in_flit_bits_egress_id,
  output        auto_routers_source_nodes_out_flit_0_valid,
  output        auto_routers_source_nodes_out_flit_0_bits_head,
  output        auto_routers_source_nodes_out_flit_0_bits_tail,
  output [63:0] auto_routers_source_nodes_out_flit_0_bits_payload,
  output        auto_routers_source_nodes_out_flit_0_bits_flow_ingress_node,
  output        auto_routers_source_nodes_out_flit_0_bits_flow_egress_node,
  output [1:0]  auto_routers_source_nodes_out_flit_0_bits_virt_channel_id,
  input  [2:0]  auto_routers_source_nodes_out_credit_return,
  input  [2:0]  auto_routers_source_nodes_out_vc_free,
  input         auto_clock_in_clock,
  input         auto_clock_in_reset
);
  wire  routers_clock; // @[NoC.scala 64:22]
  wire  routers_reset; // @[NoC.scala 64:22]
  wire  routers_auto_ingress_nodes_in_flit_ready; // @[NoC.scala 64:22]
  wire  routers_auto_ingress_nodes_in_flit_valid; // @[NoC.scala 64:22]
  wire  routers_auto_ingress_nodes_in_flit_bits_head; // @[NoC.scala 64:22]
  wire  routers_auto_ingress_nodes_in_flit_bits_tail; // @[NoC.scala 64:22]
  wire [63:0] routers_auto_ingress_nodes_in_flit_bits_payload; // @[NoC.scala 64:22]
  wire  routers_auto_ingress_nodes_in_flit_bits_egress_id; // @[NoC.scala 64:22]
  wire  routers_auto_source_nodes_out_flit_0_valid; // @[NoC.scala 64:22]
  wire  routers_auto_source_nodes_out_flit_0_bits_head; // @[NoC.scala 64:22]
  wire  routers_auto_source_nodes_out_flit_0_bits_tail; // @[NoC.scala 64:22]
  wire [63:0] routers_auto_source_nodes_out_flit_0_bits_payload; // @[NoC.scala 64:22]
  wire  routers_auto_source_nodes_out_flit_0_bits_flow_ingress_node; // @[NoC.scala 64:22]
  wire  routers_auto_source_nodes_out_flit_0_bits_flow_egress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_source_nodes_out_flit_0_bits_virt_channel_id; // @[NoC.scala 64:22]
  wire [2:0] routers_auto_source_nodes_out_credit_return; // @[NoC.scala 64:22]
  wire [2:0] routers_auto_source_nodes_out_vc_free; // @[NoC.scala 64:22]
  Router routers ( // @[NoC.scala 64:22]
    .clock(routers_clock),
    .reset(routers_reset),
    .auto_ingress_nodes_in_flit_ready(routers_auto_ingress_nodes_in_flit_ready),
    .auto_ingress_nodes_in_flit_valid(routers_auto_ingress_nodes_in_flit_valid),
    .auto_ingress_nodes_in_flit_bits_head(routers_auto_ingress_nodes_in_flit_bits_head),
    .auto_ingress_nodes_in_flit_bits_tail(routers_auto_ingress_nodes_in_flit_bits_tail),
    .auto_ingress_nodes_in_flit_bits_payload(routers_auto_ingress_nodes_in_flit_bits_payload),
    .auto_ingress_nodes_in_flit_bits_egress_id(routers_auto_ingress_nodes_in_flit_bits_egress_id),
    .auto_source_nodes_out_flit_0_valid(routers_auto_source_nodes_out_flit_0_valid),
    .auto_source_nodes_out_flit_0_bits_head(routers_auto_source_nodes_out_flit_0_bits_head),
    .auto_source_nodes_out_flit_0_bits_tail(routers_auto_source_nodes_out_flit_0_bits_tail),
    .auto_source_nodes_out_flit_0_bits_payload(routers_auto_source_nodes_out_flit_0_bits_payload),
    .auto_source_nodes_out_flit_0_bits_flow_ingress_node(routers_auto_source_nodes_out_flit_0_bits_flow_ingress_node),
    .auto_source_nodes_out_flit_0_bits_flow_egress_node(routers_auto_source_nodes_out_flit_0_bits_flow_egress_node),
    .auto_source_nodes_out_flit_0_bits_virt_channel_id(routers_auto_source_nodes_out_flit_0_bits_virt_channel_id),
    .auto_source_nodes_out_credit_return(routers_auto_source_nodes_out_credit_return),
    .auto_source_nodes_out_vc_free(routers_auto_source_nodes_out_vc_free)
  );
  assign auto_routers_ingress_nodes_in_flit_ready = routers_auto_ingress_nodes_in_flit_ready; // @[LazyModule.scala 366:16]
  assign auto_routers_source_nodes_out_flit_0_valid = routers_auto_source_nodes_out_flit_0_valid; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_flit_0_bits_head = routers_auto_source_nodes_out_flit_0_bits_head; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_flit_0_bits_tail = routers_auto_source_nodes_out_flit_0_bits_tail; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_flit_0_bits_payload = routers_auto_source_nodes_out_flit_0_bits_payload; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_flit_0_bits_flow_ingress_node =
    routers_auto_source_nodes_out_flit_0_bits_flow_ingress_node; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_flit_0_bits_flow_egress_node =
    routers_auto_source_nodes_out_flit_0_bits_flow_egress_node; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_flit_0_bits_virt_channel_id =
    routers_auto_source_nodes_out_flit_0_bits_virt_channel_id; // @[LazyModule.scala 368:12]
  assign routers_clock = auto_clock_in_clock; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign routers_reset = auto_clock_in_reset; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign routers_auto_ingress_nodes_in_flit_valid = auto_routers_ingress_nodes_in_flit_valid; // @[LazyModule.scala 366:16]
  assign routers_auto_ingress_nodes_in_flit_bits_head = auto_routers_ingress_nodes_in_flit_bits_head; // @[LazyModule.scala 366:16]
  assign routers_auto_ingress_nodes_in_flit_bits_tail = auto_routers_ingress_nodes_in_flit_bits_tail; // @[LazyModule.scala 366:16]
  assign routers_auto_ingress_nodes_in_flit_bits_payload = auto_routers_ingress_nodes_in_flit_bits_payload; // @[LazyModule.scala 366:16]
  assign routers_auto_ingress_nodes_in_flit_bits_egress_id = auto_routers_ingress_nodes_in_flit_bits_egress_id; // @[LazyModule.scala 366:16]
  assign routers_auto_source_nodes_out_credit_return = auto_routers_source_nodes_out_credit_return; // @[LazyModule.scala 368:12]
  assign routers_auto_source_nodes_out_vc_free = auto_routers_source_nodes_out_vc_free; // @[LazyModule.scala 368:12]
endmodule
module NoCMonitor(
  input        clock,
  input        reset,
  input        io_in_flit_0_valid,
  input        io_in_flit_0_bits_head,
  input        io_in_flit_0_bits_tail,
  input        io_in_flit_0_bits_flow_ingress_node,
  input        io_in_flit_0_bits_flow_egress_node,
  input  [1:0] io_in_flit_0_bits_virt_channel_id
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg  in_flight_0; // @[Monitor.scala 16:26]
  reg  in_flight_1; // @[Monitor.scala 16:26]
  reg  in_flight_2; // @[Monitor.scala 16:26]
  wire  _GEN_0 = 2'h0 == io_in_flit_0_bits_virt_channel_id | in_flight_0; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_1 = 2'h1 == io_in_flit_0_bits_virt_channel_id | in_flight_1; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_2 = 2'h2 == io_in_flit_0_bits_virt_channel_id | in_flight_2; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_4 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? in_flight_1 : in_flight_0; // @[Monitor.scala 22:{17,17}]
  wire  _GEN_5 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? in_flight_2 : _GEN_4; // @[Monitor.scala 22:{17,17}]
  wire  _T_2 = ~reset; // @[Monitor.scala 22:16]
  wire  _GEN_6 = io_in_flit_0_bits_head ? _GEN_0 : in_flight_0; // @[Monitor.scala 16:26 20:29]
  wire  _GEN_7 = io_in_flit_0_bits_head ? _GEN_1 : in_flight_1; // @[Monitor.scala 16:26 20:29]
  wire  _GEN_8 = io_in_flit_0_bits_head ? _GEN_2 : in_flight_2; // @[Monitor.scala 16:26 20:29]
  wire  _T_4 = io_in_flit_0_valid & io_in_flit_0_bits_head; // @[Monitor.scala 29:22]
  wire  _T_8 = ~io_in_flit_0_bits_flow_ingress_node & io_in_flit_0_bits_flow_egress_node; // @[Types.scala 53:39]
  wire  _GEN_22 = _T_4 & ~reset; // @[Monitor.scala 22:16]
  always @(posedge clock) begin
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_0 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h0 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_0 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_0 <= _GEN_6;
        end
      end else begin
        in_flight_0 <= _GEN_6;
      end
    end
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_1 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h1 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_1 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_1 <= _GEN_7;
        end
      end else begin
        in_flight_1 <= _GEN_7;
      end
    end
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_2 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h2 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_2 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_2 <= _GEN_8;
        end
      end else begin
        in_flight_2 <= _GEN_8;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4 & ~reset & ~(~_GEN_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed: Flit head/tail sequencing is broken\n    at Monitor.scala:22 assert (!in_flight(flit.bits.virt_channel_id), \"Flit head/tail sequencing is broken\")\n"
            ); // @[Monitor.scala 22:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_22 & ~(io_in_flit_0_bits_virt_channel_id != 2'h0 | _T_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_22 & ~(io_in_flit_0_bits_virt_channel_id != 2'h1 | _T_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_22 & ~(io_in_flit_0_bits_virt_channel_id != 2'h2 | _T_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  in_flight_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  in_flight_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  in_flight_2 = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (_T_4 & ~reset) begin
      assert(~_GEN_5); // @[Monitor.scala 22:16]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h0 | _T_8); // @[Monitor.scala 32:17]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h1 | _T_8); // @[Monitor.scala 32:17]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h2 | _T_8); // @[Monitor.scala 32:17]
    end
  end
endmodule
module Queue_4(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_head,
  input         io_enq_bits_tail,
  input  [63:0] io_enq_bits_payload,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_head,
  output        io_deq_bits_tail,
  output [63:0] io_deq_bits_payload
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg  ram_head [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_head_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_head_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_head_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_tail [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_tail_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_tail_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_tail_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_en; // @[Decoupled.scala 273:95]
  reg [63:0] ram_payload [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_payload_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_payload_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [63:0] ram_payload_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [63:0] ram_payload_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_payload_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_payload_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_payload_MPORT_en; // @[Decoupled.scala 273:95]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 278:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  assign ram_head_io_deq_bits_MPORT_en = 1'h1;
  assign ram_head_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_head_io_deq_bits_MPORT_data = ram_head[ram_head_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_head_MPORT_data = io_enq_bits_head;
  assign ram_head_MPORT_addr = 1'h0;
  assign ram_head_MPORT_mask = 1'h1;
  assign ram_head_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tail_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tail_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tail_io_deq_bits_MPORT_data = ram_tail[ram_tail_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_tail_MPORT_data = io_enq_bits_tail;
  assign ram_tail_MPORT_addr = 1'h0;
  assign ram_tail_MPORT_mask = 1'h1;
  assign ram_tail_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_payload_io_deq_bits_MPORT_en = 1'h1;
  assign ram_payload_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_payload_io_deq_bits_MPORT_data = ram_payload[ram_payload_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_payload_MPORT_data = io_enq_bits_payload;
  assign ram_payload_MPORT_addr = 1'h0;
  assign ram_payload_MPORT_mask = 1'h1;
  assign ram_payload_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = io_deq_ready | empty; // @[Decoupled.scala 303:16 323:{24,39}]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_head = ram_head_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_tail = ram_tail_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_payload = ram_payload_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  always @(posedge clock) begin
    if (ram_head_MPORT_en & ram_head_MPORT_mask) begin
      ram_head[ram_head_MPORT_addr] <= ram_head_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_tail_MPORT_en & ram_tail_MPORT_mask) begin
      ram_tail[ram_tail_MPORT_addr] <= ram_tail_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_payload_MPORT_en & ram_payload_MPORT_mask) begin
      ram_payload[ram_payload_MPORT_addr] <= ram_payload_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_head[initvar] = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tail[initvar] = _RAND_1[0:0];
  _RAND_2 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload[initvar] = _RAND_2[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module InputBuffer(
  input         clock,
  input         reset,
  input         io_enq_0_valid,
  input         io_enq_0_bits_head,
  input         io_enq_0_bits_tail,
  input  [63:0] io_enq_0_bits_payload,
  input  [1:0]  io_enq_0_bits_virt_channel_id,
  input         io_deq_0_ready,
  output        io_deq_0_valid,
  output        io_deq_0_bits_head,
  output        io_deq_0_bits_tail,
  output [63:0] io_deq_0_bits_payload,
  input         io_deq_1_ready,
  output        io_deq_1_valid,
  output        io_deq_1_bits_head,
  output        io_deq_1_bits_tail,
  output [63:0] io_deq_1_bits_payload,
  input         io_deq_2_ready,
  output        io_deq_2_valid,
  output        io_deq_2_bits_head,
  output        io_deq_2_bits_tail,
  output [63:0] io_deq_2_bits_payload
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_8;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  reg  mem_head [0:8]; // @[InputUnit.scala 85:18]
  wire  mem_head_qs_0_io_enq_bits_MPORT_en; // @[InputUnit.scala 85:18]
  wire [3:0] mem_head_qs_0_io_enq_bits_MPORT_addr; // @[InputUnit.scala 85:18]
  wire  mem_head_qs_0_io_enq_bits_MPORT_data; // @[InputUnit.scala 85:18]
  wire  mem_head_qs_1_io_enq_bits_MPORT_en; // @[InputUnit.scala 85:18]
  wire [3:0] mem_head_qs_1_io_enq_bits_MPORT_addr; // @[InputUnit.scala 85:18]
  wire  mem_head_qs_1_io_enq_bits_MPORT_data; // @[InputUnit.scala 85:18]
  wire  mem_head_qs_2_io_enq_bits_MPORT_en; // @[InputUnit.scala 85:18]
  wire [3:0] mem_head_qs_2_io_enq_bits_MPORT_addr; // @[InputUnit.scala 85:18]
  wire  mem_head_qs_2_io_enq_bits_MPORT_data; // @[InputUnit.scala 85:18]
  wire  mem_head_MPORT_data; // @[InputUnit.scala 85:18]
  wire [3:0] mem_head_MPORT_addr; // @[InputUnit.scala 85:18]
  wire  mem_head_MPORT_mask; // @[InputUnit.scala 85:18]
  wire  mem_head_MPORT_en; // @[InputUnit.scala 85:18]
  reg  mem_tail [0:8]; // @[InputUnit.scala 85:18]
  wire  mem_tail_qs_0_io_enq_bits_MPORT_en; // @[InputUnit.scala 85:18]
  wire [3:0] mem_tail_qs_0_io_enq_bits_MPORT_addr; // @[InputUnit.scala 85:18]
  wire  mem_tail_qs_0_io_enq_bits_MPORT_data; // @[InputUnit.scala 85:18]
  wire  mem_tail_qs_1_io_enq_bits_MPORT_en; // @[InputUnit.scala 85:18]
  wire [3:0] mem_tail_qs_1_io_enq_bits_MPORT_addr; // @[InputUnit.scala 85:18]
  wire  mem_tail_qs_1_io_enq_bits_MPORT_data; // @[InputUnit.scala 85:18]
  wire  mem_tail_qs_2_io_enq_bits_MPORT_en; // @[InputUnit.scala 85:18]
  wire [3:0] mem_tail_qs_2_io_enq_bits_MPORT_addr; // @[InputUnit.scala 85:18]
  wire  mem_tail_qs_2_io_enq_bits_MPORT_data; // @[InputUnit.scala 85:18]
  wire  mem_tail_MPORT_data; // @[InputUnit.scala 85:18]
  wire [3:0] mem_tail_MPORT_addr; // @[InputUnit.scala 85:18]
  wire  mem_tail_MPORT_mask; // @[InputUnit.scala 85:18]
  wire  mem_tail_MPORT_en; // @[InputUnit.scala 85:18]
  reg [63:0] mem_payload [0:8]; // @[InputUnit.scala 85:18]
  wire  mem_payload_qs_0_io_enq_bits_MPORT_en; // @[InputUnit.scala 85:18]
  wire [3:0] mem_payload_qs_0_io_enq_bits_MPORT_addr; // @[InputUnit.scala 85:18]
  wire [63:0] mem_payload_qs_0_io_enq_bits_MPORT_data; // @[InputUnit.scala 85:18]
  wire  mem_payload_qs_1_io_enq_bits_MPORT_en; // @[InputUnit.scala 85:18]
  wire [3:0] mem_payload_qs_1_io_enq_bits_MPORT_addr; // @[InputUnit.scala 85:18]
  wire [63:0] mem_payload_qs_1_io_enq_bits_MPORT_data; // @[InputUnit.scala 85:18]
  wire  mem_payload_qs_2_io_enq_bits_MPORT_en; // @[InputUnit.scala 85:18]
  wire [3:0] mem_payload_qs_2_io_enq_bits_MPORT_addr; // @[InputUnit.scala 85:18]
  wire [63:0] mem_payload_qs_2_io_enq_bits_MPORT_data; // @[InputUnit.scala 85:18]
  wire [63:0] mem_payload_MPORT_data; // @[InputUnit.scala 85:18]
  wire [3:0] mem_payload_MPORT_addr; // @[InputUnit.scala 85:18]
  wire  mem_payload_MPORT_mask; // @[InputUnit.scala 85:18]
  wire  mem_payload_MPORT_en; // @[InputUnit.scala 85:18]
  wire  qs_0_clock; // @[InputUnit.scala 90:49]
  wire  qs_0_reset; // @[InputUnit.scala 90:49]
  wire  qs_0_io_enq_ready; // @[InputUnit.scala 90:49]
  wire  qs_0_io_enq_valid; // @[InputUnit.scala 90:49]
  wire  qs_0_io_enq_bits_head; // @[InputUnit.scala 90:49]
  wire  qs_0_io_enq_bits_tail; // @[InputUnit.scala 90:49]
  wire [63:0] qs_0_io_enq_bits_payload; // @[InputUnit.scala 90:49]
  wire  qs_0_io_deq_ready; // @[InputUnit.scala 90:49]
  wire  qs_0_io_deq_valid; // @[InputUnit.scala 90:49]
  wire  qs_0_io_deq_bits_head; // @[InputUnit.scala 90:49]
  wire  qs_0_io_deq_bits_tail; // @[InputUnit.scala 90:49]
  wire [63:0] qs_0_io_deq_bits_payload; // @[InputUnit.scala 90:49]
  wire  qs_1_clock; // @[InputUnit.scala 90:49]
  wire  qs_1_reset; // @[InputUnit.scala 90:49]
  wire  qs_1_io_enq_ready; // @[InputUnit.scala 90:49]
  wire  qs_1_io_enq_valid; // @[InputUnit.scala 90:49]
  wire  qs_1_io_enq_bits_head; // @[InputUnit.scala 90:49]
  wire  qs_1_io_enq_bits_tail; // @[InputUnit.scala 90:49]
  wire [63:0] qs_1_io_enq_bits_payload; // @[InputUnit.scala 90:49]
  wire  qs_1_io_deq_ready; // @[InputUnit.scala 90:49]
  wire  qs_1_io_deq_valid; // @[InputUnit.scala 90:49]
  wire  qs_1_io_deq_bits_head; // @[InputUnit.scala 90:49]
  wire  qs_1_io_deq_bits_tail; // @[InputUnit.scala 90:49]
  wire [63:0] qs_1_io_deq_bits_payload; // @[InputUnit.scala 90:49]
  wire  qs_2_clock; // @[InputUnit.scala 90:49]
  wire  qs_2_reset; // @[InputUnit.scala 90:49]
  wire  qs_2_io_enq_ready; // @[InputUnit.scala 90:49]
  wire  qs_2_io_enq_valid; // @[InputUnit.scala 90:49]
  wire  qs_2_io_enq_bits_head; // @[InputUnit.scala 90:49]
  wire  qs_2_io_enq_bits_tail; // @[InputUnit.scala 90:49]
  wire [63:0] qs_2_io_enq_bits_payload; // @[InputUnit.scala 90:49]
  wire  qs_2_io_deq_ready; // @[InputUnit.scala 90:49]
  wire  qs_2_io_deq_valid; // @[InputUnit.scala 90:49]
  wire  qs_2_io_deq_bits_head; // @[InputUnit.scala 90:49]
  wire  qs_2_io_deq_bits_tail; // @[InputUnit.scala 90:49]
  wire [63:0] qs_2_io_deq_bits_payload; // @[InputUnit.scala 90:49]
  reg [3:0] heads_0; // @[InputUnit.scala 86:24]
  reg [3:0] heads_1; // @[InputUnit.scala 86:24]
  reg [3:0] heads_2; // @[InputUnit.scala 86:24]
  reg [3:0] tails_0; // @[InputUnit.scala 87:24]
  reg [3:0] tails_1; // @[InputUnit.scala 87:24]
  reg [3:0] tails_2; // @[InputUnit.scala 87:24]
  wire  empty_0 = heads_0 == tails_0; // @[InputUnit.scala 88:49]
  wire  empty_1 = heads_1 == tails_1; // @[InputUnit.scala 88:49]
  wire  empty_2 = heads_2 == tails_2; // @[InputUnit.scala 88:49]
  wire [3:0] vc_sel = 4'h1 << io_enq_0_bits_virt_channel_id; // @[OneHot.scala 57:35]
  wire  _direct_to_q_T_7 = vc_sel[0] & qs_0_io_enq_ready | vc_sel[1] & qs_1_io_enq_ready | vc_sel[2] & qs_2_io_enq_ready
    ; // @[Mux.scala 27:73]
  wire  _direct_to_q_T_15 = vc_sel[0] & empty_0 | vc_sel[1] & empty_1 | vc_sel[2] & empty_2; // @[Mux.scala 27:73]
  wire  direct_to_q = _direct_to_q_T_7 & _direct_to_q_T_15; // @[InputUnit.scala 96:62]
  wire  _T = ~direct_to_q; // @[InputUnit.scala 100:30]
  wire [3:0] _GEN_1 = 2'h1 == io_enq_0_bits_virt_channel_id ? tails_1 : tails_0; // @[]
  wire [3:0] _GEN_2 = 2'h2 == io_enq_0_bits_virt_channel_id ? tails_2 : _GEN_1; // @[]
  wire [1:0] _tails_T_3 = vc_sel[0] ? 2'h2 : 2'h0; // @[Mux.scala 27:73]
  wire [2:0] _tails_T_4 = vc_sel[1] ? 3'h5 : 3'h0; // @[Mux.scala 27:73]
  wire [3:0] _tails_T_5 = vc_sel[2] ? 4'h8 : 4'h0; // @[Mux.scala 27:73]
  wire [2:0] _GEN_100 = {{1'd0}, _tails_T_3}; // @[Mux.scala 27:73]
  wire [2:0] _tails_T_6 = _GEN_100 | _tails_T_4; // @[Mux.scala 27:73]
  wire [3:0] _GEN_101 = {{1'd0}, _tails_T_6}; // @[Mux.scala 27:73]
  wire [3:0] _tails_T_7 = _GEN_101 | _tails_T_5; // @[Mux.scala 27:73]
  wire  _tails_T_8 = _GEN_2 == _tails_T_7; // @[InputUnit.scala 104:14]
  wire [1:0] _tails_T_13 = vc_sel[1] ? 2'h3 : 2'h0; // @[Mux.scala 27:73]
  wire [2:0] _tails_T_14 = vc_sel[2] ? 3'h6 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _GEN_102 = {{1'd0}, _tails_T_13}; // @[Mux.scala 27:73]
  wire [2:0] _tails_T_16 = _GEN_102 | _tails_T_14; // @[Mux.scala 27:73]
  wire [3:0] _tails_T_18 = _GEN_2 + 4'h1; // @[InputUnit.scala 106:14]
  wire  _T_3 = io_enq_0_bits_virt_channel_id == 2'h0; // @[InputUnit.scala 109:46]
  wire  _T_4 = io_enq_0_bits_virt_channel_id == 2'h1; // @[InputUnit.scala 109:46]
  wire  _T_5 = io_enq_0_bits_virt_channel_id == 2'h2; // @[InputUnit.scala 109:46]
  wire  _GEN_18 = io_enq_0_valid & direct_to_q & _T_3; // @[InputUnit.scala 107:50 91:31]
  wire  _GEN_22 = io_enq_0_valid & direct_to_q & _T_4; // @[InputUnit.scala 107:50 91:31]
  wire  _GEN_26 = io_enq_0_valid & direct_to_q & _T_5; // @[InputUnit.scala 107:50 91:31]
  wire  _GEN_40 = io_enq_0_valid & ~direct_to_q ? 1'h0 : _GEN_18; // @[InputUnit.scala 100:44 91:31]
  wire  _GEN_44 = io_enq_0_valid & ~direct_to_q ? 1'h0 : _GEN_22; // @[InputUnit.scala 100:44 91:31]
  wire  _GEN_48 = io_enq_0_valid & ~direct_to_q ? 1'h0 : _GEN_26; // @[InputUnit.scala 100:44 91:31]
  wire  can_to_q_0 = ~empty_0 & qs_0_io_enq_ready; // @[InputUnit.scala 117:70]
  wire  can_to_q_1 = ~empty_1 & qs_1_io_enq_ready; // @[InputUnit.scala 117:70]
  wire  can_to_q_2 = ~empty_2 & qs_2_io_enq_ready; // @[InputUnit.scala 117:70]
  wire [2:0] _to_q_oh_enc_T = can_to_q_2 ? 3'h4 : 3'h0; // @[Mux.scala 47:70]
  wire [2:0] _to_q_oh_enc_T_1 = can_to_q_1 ? 3'h2 : _to_q_oh_enc_T; // @[Mux.scala 47:70]
  wire [2:0] to_q_oh_enc = can_to_q_0 ? 3'h1 : _to_q_oh_enc_T_1; // @[Mux.scala 47:70]
  wire  to_q_oh_0 = to_q_oh_enc[0]; // @[OneHot.scala 82:30]
  wire  to_q_oh_1 = to_q_oh_enc[1]; // @[OneHot.scala 82:30]
  wire  to_q_oh_2 = to_q_oh_enc[2]; // @[OneHot.scala 82:30]
  wire [2:0] _to_q_T = {to_q_oh_2,to_q_oh_1,to_q_oh_0}; // @[Cat.scala 33:92]
  wire  to_q_hi_1 = _to_q_T[2]; // @[OneHot.scala 30:18]
  wire [1:0] to_q_lo = _to_q_T[1:0]; // @[OneHot.scala 31:18]
  wire  _to_q_T_1 = |to_q_hi_1; // @[OneHot.scala 32:14]
  wire [1:0] _GEN_103 = {{1'd0}, to_q_hi_1}; // @[OneHot.scala 32:28]
  wire [1:0] _to_q_T_2 = _GEN_103 | to_q_lo; // @[OneHot.scala 32:28]
  wire [1:0] to_q = {_to_q_T_1,_to_q_T_2[1]}; // @[Cat.scala 33:92]
  wire  _T_7 = can_to_q_0 | can_to_q_1 | can_to_q_2; // @[package.scala 73:59]
  wire [3:0] _head_T = to_q_oh_0 ? heads_0 : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _head_T_1 = to_q_oh_1 ? heads_1 : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _head_T_2 = to_q_oh_2 ? heads_2 : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _head_T_3 = _head_T | _head_T_1; // @[Mux.scala 27:73]
  wire [3:0] head = _head_T_3 | _head_T_2; // @[Mux.scala 27:73]
  wire [1:0] _heads_T = to_q_oh_0 ? 2'h2 : 2'h0; // @[Mux.scala 27:73]
  wire [2:0] _heads_T_1 = to_q_oh_1 ? 3'h5 : 3'h0; // @[Mux.scala 27:73]
  wire [3:0] _heads_T_2 = to_q_oh_2 ? 4'h8 : 4'h0; // @[Mux.scala 27:73]
  wire [2:0] _GEN_104 = {{1'd0}, _heads_T}; // @[Mux.scala 27:73]
  wire [2:0] _heads_T_3 = _GEN_104 | _heads_T_1; // @[Mux.scala 27:73]
  wire [3:0] _GEN_105 = {{1'd0}, _heads_T_3}; // @[Mux.scala 27:73]
  wire [3:0] _heads_T_4 = _GEN_105 | _heads_T_2; // @[Mux.scala 27:73]
  wire  _heads_T_5 = head == _heads_T_4; // @[InputUnit.scala 123:16]
  wire [1:0] _heads_T_7 = to_q_oh_1 ? 2'h3 : 2'h0; // @[Mux.scala 27:73]
  wire [2:0] _heads_T_8 = to_q_oh_2 ? 3'h6 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _GEN_106 = {{1'd0}, _heads_T_7}; // @[Mux.scala 27:73]
  wire [2:0] _heads_T_10 = _GEN_106 | _heads_T_8; // @[Mux.scala 27:73]
  wire [3:0] _heads_T_12 = head + 4'h1; // @[InputUnit.scala 125:16]
  wire  _GEN_55 = to_q_oh_0 | _GEN_40; // @[InputUnit.scala 127:29 128:32]
  wire [63:0] _GEN_59 = to_q_oh_0 ? mem_payload_qs_0_io_enq_bits_MPORT_data : io_enq_0_bits_payload; // @[InputUnit.scala 127:29 129:31]
  wire  _GEN_60 = to_q_oh_0 ? mem_tail_qs_0_io_enq_bits_MPORT_data : io_enq_0_bits_tail; // @[InputUnit.scala 127:29 129:31]
  wire  _GEN_61 = to_q_oh_0 ? mem_head_qs_0_io_enq_bits_MPORT_data : io_enq_0_bits_head; // @[InputUnit.scala 127:29 129:31]
  wire  _GEN_62 = to_q_oh_1 | _GEN_44; // @[InputUnit.scala 127:29 128:32]
  wire [63:0] _GEN_66 = to_q_oh_1 ? mem_payload_qs_1_io_enq_bits_MPORT_data : io_enq_0_bits_payload; // @[InputUnit.scala 127:29 129:31]
  wire  _GEN_67 = to_q_oh_1 ? mem_tail_qs_1_io_enq_bits_MPORT_data : io_enq_0_bits_tail; // @[InputUnit.scala 127:29 129:31]
  wire  _GEN_68 = to_q_oh_1 ? mem_head_qs_1_io_enq_bits_MPORT_data : io_enq_0_bits_head; // @[InputUnit.scala 127:29 129:31]
  wire  _GEN_69 = to_q_oh_2 | _GEN_48; // @[InputUnit.scala 127:29 128:32]
  wire [63:0] _GEN_73 = to_q_oh_2 ? mem_payload_qs_2_io_enq_bits_MPORT_data : io_enq_0_bits_payload; // @[InputUnit.scala 127:29 129:31]
  wire  _GEN_74 = to_q_oh_2 ? mem_tail_qs_2_io_enq_bits_MPORT_data : io_enq_0_bits_tail; // @[InputUnit.scala 127:29 129:31]
  wire  _GEN_75 = to_q_oh_2 ? mem_head_qs_2_io_enq_bits_MPORT_data : io_enq_0_bits_head; // @[InputUnit.scala 127:29 129:31]
  Queue_4 qs_0 ( // @[InputUnit.scala 90:49]
    .clock(qs_0_clock),
    .reset(qs_0_reset),
    .io_enq_ready(qs_0_io_enq_ready),
    .io_enq_valid(qs_0_io_enq_valid),
    .io_enq_bits_head(qs_0_io_enq_bits_head),
    .io_enq_bits_tail(qs_0_io_enq_bits_tail),
    .io_enq_bits_payload(qs_0_io_enq_bits_payload),
    .io_deq_ready(qs_0_io_deq_ready),
    .io_deq_valid(qs_0_io_deq_valid),
    .io_deq_bits_head(qs_0_io_deq_bits_head),
    .io_deq_bits_tail(qs_0_io_deq_bits_tail),
    .io_deq_bits_payload(qs_0_io_deq_bits_payload)
  );
  Queue_4 qs_1 ( // @[InputUnit.scala 90:49]
    .clock(qs_1_clock),
    .reset(qs_1_reset),
    .io_enq_ready(qs_1_io_enq_ready),
    .io_enq_valid(qs_1_io_enq_valid),
    .io_enq_bits_head(qs_1_io_enq_bits_head),
    .io_enq_bits_tail(qs_1_io_enq_bits_tail),
    .io_enq_bits_payload(qs_1_io_enq_bits_payload),
    .io_deq_ready(qs_1_io_deq_ready),
    .io_deq_valid(qs_1_io_deq_valid),
    .io_deq_bits_head(qs_1_io_deq_bits_head),
    .io_deq_bits_tail(qs_1_io_deq_bits_tail),
    .io_deq_bits_payload(qs_1_io_deq_bits_payload)
  );
  Queue_4 qs_2 ( // @[InputUnit.scala 90:49]
    .clock(qs_2_clock),
    .reset(qs_2_reset),
    .io_enq_ready(qs_2_io_enq_ready),
    .io_enq_valid(qs_2_io_enq_valid),
    .io_enq_bits_head(qs_2_io_enq_bits_head),
    .io_enq_bits_tail(qs_2_io_enq_bits_tail),
    .io_enq_bits_payload(qs_2_io_enq_bits_payload),
    .io_deq_ready(qs_2_io_deq_ready),
    .io_deq_valid(qs_2_io_deq_valid),
    .io_deq_bits_head(qs_2_io_deq_bits_head),
    .io_deq_bits_tail(qs_2_io_deq_bits_tail),
    .io_deq_bits_payload(qs_2_io_deq_bits_payload)
  );
  assign mem_head_qs_0_io_enq_bits_MPORT_en = _T_7 & to_q_oh_0;
  assign mem_head_qs_0_io_enq_bits_MPORT_addr = _head_T_3 | _head_T_2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_head_qs_0_io_enq_bits_MPORT_data = mem_head[mem_head_qs_0_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `else
  assign mem_head_qs_0_io_enq_bits_MPORT_data = mem_head_qs_0_io_enq_bits_MPORT_addr >= 4'h9 ? _RAND_1[0:0] :
    mem_head[mem_head_qs_0_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_head_qs_1_io_enq_bits_MPORT_en = _T_7 & to_q_oh_1;
  assign mem_head_qs_1_io_enq_bits_MPORT_addr = _head_T_3 | _head_T_2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_head_qs_1_io_enq_bits_MPORT_data = mem_head[mem_head_qs_1_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `else
  assign mem_head_qs_1_io_enq_bits_MPORT_data = mem_head_qs_1_io_enq_bits_MPORT_addr >= 4'h9 ? _RAND_2[0:0] :
    mem_head[mem_head_qs_1_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_head_qs_2_io_enq_bits_MPORT_en = _T_7 & to_q_oh_2;
  assign mem_head_qs_2_io_enq_bits_MPORT_addr = _head_T_3 | _head_T_2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_head_qs_2_io_enq_bits_MPORT_data = mem_head[mem_head_qs_2_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `else
  assign mem_head_qs_2_io_enq_bits_MPORT_data = mem_head_qs_2_io_enq_bits_MPORT_addr >= 4'h9 ? _RAND_3[0:0] :
    mem_head[mem_head_qs_2_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_head_MPORT_data = io_enq_0_bits_head;
  assign mem_head_MPORT_addr = 2'h2 == io_enq_0_bits_virt_channel_id ? tails_2 : _GEN_1;
  assign mem_head_MPORT_mask = 1'h1;
  assign mem_head_MPORT_en = io_enq_0_valid & _T;
  assign mem_tail_qs_0_io_enq_bits_MPORT_en = _T_7 & to_q_oh_0;
  assign mem_tail_qs_0_io_enq_bits_MPORT_addr = _head_T_3 | _head_T_2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_tail_qs_0_io_enq_bits_MPORT_data = mem_tail[mem_tail_qs_0_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `else
  assign mem_tail_qs_0_io_enq_bits_MPORT_data = mem_tail_qs_0_io_enq_bits_MPORT_addr >= 4'h9 ? _RAND_5[0:0] :
    mem_tail[mem_tail_qs_0_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_tail_qs_1_io_enq_bits_MPORT_en = _T_7 & to_q_oh_1;
  assign mem_tail_qs_1_io_enq_bits_MPORT_addr = _head_T_3 | _head_T_2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_tail_qs_1_io_enq_bits_MPORT_data = mem_tail[mem_tail_qs_1_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `else
  assign mem_tail_qs_1_io_enq_bits_MPORT_data = mem_tail_qs_1_io_enq_bits_MPORT_addr >= 4'h9 ? _RAND_6[0:0] :
    mem_tail[mem_tail_qs_1_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_tail_qs_2_io_enq_bits_MPORT_en = _T_7 & to_q_oh_2;
  assign mem_tail_qs_2_io_enq_bits_MPORT_addr = _head_T_3 | _head_T_2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_tail_qs_2_io_enq_bits_MPORT_data = mem_tail[mem_tail_qs_2_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `else
  assign mem_tail_qs_2_io_enq_bits_MPORT_data = mem_tail_qs_2_io_enq_bits_MPORT_addr >= 4'h9 ? _RAND_7[0:0] :
    mem_tail[mem_tail_qs_2_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_tail_MPORT_data = io_enq_0_bits_tail;
  assign mem_tail_MPORT_addr = 2'h2 == io_enq_0_bits_virt_channel_id ? tails_2 : _GEN_1;
  assign mem_tail_MPORT_mask = 1'h1;
  assign mem_tail_MPORT_en = io_enq_0_valid & _T;
  assign mem_payload_qs_0_io_enq_bits_MPORT_en = _T_7 & to_q_oh_0;
  assign mem_payload_qs_0_io_enq_bits_MPORT_addr = _head_T_3 | _head_T_2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_payload_qs_0_io_enq_bits_MPORT_data = mem_payload[mem_payload_qs_0_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `else
  assign mem_payload_qs_0_io_enq_bits_MPORT_data = mem_payload_qs_0_io_enq_bits_MPORT_addr >= 4'h9 ? _RAND_9[63:0] :
    mem_payload[mem_payload_qs_0_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_payload_qs_1_io_enq_bits_MPORT_en = _T_7 & to_q_oh_1;
  assign mem_payload_qs_1_io_enq_bits_MPORT_addr = _head_T_3 | _head_T_2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_payload_qs_1_io_enq_bits_MPORT_data = mem_payload[mem_payload_qs_1_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `else
  assign mem_payload_qs_1_io_enq_bits_MPORT_data = mem_payload_qs_1_io_enq_bits_MPORT_addr >= 4'h9 ? _RAND_10[63:0] :
    mem_payload[mem_payload_qs_1_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_payload_qs_2_io_enq_bits_MPORT_en = _T_7 & to_q_oh_2;
  assign mem_payload_qs_2_io_enq_bits_MPORT_addr = _head_T_3 | _head_T_2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_payload_qs_2_io_enq_bits_MPORT_data = mem_payload[mem_payload_qs_2_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `else
  assign mem_payload_qs_2_io_enq_bits_MPORT_data = mem_payload_qs_2_io_enq_bits_MPORT_addr >= 4'h9 ? _RAND_11[63:0] :
    mem_payload[mem_payload_qs_2_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_payload_MPORT_data = io_enq_0_bits_payload;
  assign mem_payload_MPORT_addr = 2'h2 == io_enq_0_bits_virt_channel_id ? tails_2 : _GEN_1;
  assign mem_payload_MPORT_mask = 1'h1;
  assign mem_payload_MPORT_en = io_enq_0_valid & _T;
  assign io_deq_0_valid = qs_0_io_deq_valid; // @[InputUnit.scala 134:19]
  assign io_deq_0_bits_head = qs_0_io_deq_bits_head; // @[InputUnit.scala 134:19]
  assign io_deq_0_bits_tail = qs_0_io_deq_bits_tail; // @[InputUnit.scala 134:19]
  assign io_deq_0_bits_payload = qs_0_io_deq_bits_payload; // @[InputUnit.scala 134:19]
  assign io_deq_1_valid = qs_1_io_deq_valid; // @[InputUnit.scala 134:19]
  assign io_deq_1_bits_head = qs_1_io_deq_bits_head; // @[InputUnit.scala 134:19]
  assign io_deq_1_bits_tail = qs_1_io_deq_bits_tail; // @[InputUnit.scala 134:19]
  assign io_deq_1_bits_payload = qs_1_io_deq_bits_payload; // @[InputUnit.scala 134:19]
  assign io_deq_2_valid = qs_2_io_deq_valid; // @[InputUnit.scala 134:19]
  assign io_deq_2_bits_head = qs_2_io_deq_bits_head; // @[InputUnit.scala 134:19]
  assign io_deq_2_bits_tail = qs_2_io_deq_bits_tail; // @[InputUnit.scala 134:19]
  assign io_deq_2_bits_payload = qs_2_io_deq_bits_payload; // @[InputUnit.scala 134:19]
  assign qs_0_clock = clock;
  assign qs_0_reset = reset;
  assign qs_0_io_enq_valid = _T_7 ? _GEN_55 : _GEN_40; // @[InputUnit.scala 120:27]
  assign qs_0_io_enq_bits_head = _T_7 ? _GEN_61 : io_enq_0_bits_head; // @[InputUnit.scala 120:27]
  assign qs_0_io_enq_bits_tail = _T_7 ? _GEN_60 : io_enq_0_bits_tail; // @[InputUnit.scala 120:27]
  assign qs_0_io_enq_bits_payload = _T_7 ? _GEN_59 : io_enq_0_bits_payload; // @[InputUnit.scala 120:27]
  assign qs_0_io_deq_ready = io_deq_0_ready; // @[InputUnit.scala 134:19]
  assign qs_1_clock = clock;
  assign qs_1_reset = reset;
  assign qs_1_io_enq_valid = _T_7 ? _GEN_62 : _GEN_44; // @[InputUnit.scala 120:27]
  assign qs_1_io_enq_bits_head = _T_7 ? _GEN_68 : io_enq_0_bits_head; // @[InputUnit.scala 120:27]
  assign qs_1_io_enq_bits_tail = _T_7 ? _GEN_67 : io_enq_0_bits_tail; // @[InputUnit.scala 120:27]
  assign qs_1_io_enq_bits_payload = _T_7 ? _GEN_66 : io_enq_0_bits_payload; // @[InputUnit.scala 120:27]
  assign qs_1_io_deq_ready = io_deq_1_ready; // @[InputUnit.scala 134:19]
  assign qs_2_clock = clock;
  assign qs_2_reset = reset;
  assign qs_2_io_enq_valid = _T_7 ? _GEN_69 : _GEN_48; // @[InputUnit.scala 120:27]
  assign qs_2_io_enq_bits_head = _T_7 ? _GEN_75 : io_enq_0_bits_head; // @[InputUnit.scala 120:27]
  assign qs_2_io_enq_bits_tail = _T_7 ? _GEN_74 : io_enq_0_bits_tail; // @[InputUnit.scala 120:27]
  assign qs_2_io_enq_bits_payload = _T_7 ? _GEN_73 : io_enq_0_bits_payload; // @[InputUnit.scala 120:27]
  assign qs_2_io_deq_ready = io_deq_2_ready; // @[InputUnit.scala 134:19]
  always @(posedge clock) begin
    if (mem_head_MPORT_en & mem_head_MPORT_mask) begin
      mem_head[mem_head_MPORT_addr] <= mem_head_MPORT_data; // @[InputUnit.scala 85:18]
    end
    if (mem_tail_MPORT_en & mem_tail_MPORT_mask) begin
      mem_tail[mem_tail_MPORT_addr] <= mem_tail_MPORT_data; // @[InputUnit.scala 85:18]
    end
    if (mem_payload_MPORT_en & mem_payload_MPORT_mask) begin
      mem_payload[mem_payload_MPORT_addr] <= mem_payload_MPORT_data; // @[InputUnit.scala 85:18]
    end
    if (reset) begin // @[InputUnit.scala 86:24]
      heads_0 <= 4'h0; // @[InputUnit.scala 86:24]
    end else if (_T_7) begin // @[InputUnit.scala 120:27]
      if (2'h0 == to_q) begin // @[InputUnit.scala 122:21]
        if (_heads_T_5) begin // @[InputUnit.scala 122:27]
          heads_0 <= {{1'd0}, _heads_T_10};
        end else begin
          heads_0 <= _heads_T_12;
        end
      end
    end
    if (reset) begin // @[InputUnit.scala 86:24]
      heads_1 <= 4'h3; // @[InputUnit.scala 86:24]
    end else if (_T_7) begin // @[InputUnit.scala 120:27]
      if (2'h1 == to_q) begin // @[InputUnit.scala 122:21]
        if (_heads_T_5) begin // @[InputUnit.scala 122:27]
          heads_1 <= {{1'd0}, _heads_T_10};
        end else begin
          heads_1 <= _heads_T_12;
        end
      end
    end
    if (reset) begin // @[InputUnit.scala 86:24]
      heads_2 <= 4'h6; // @[InputUnit.scala 86:24]
    end else if (_T_7) begin // @[InputUnit.scala 120:27]
      if (2'h2 == to_q) begin // @[InputUnit.scala 122:21]
        if (_heads_T_5) begin // @[InputUnit.scala 122:27]
          heads_2 <= {{1'd0}, _heads_T_10};
        end else begin
          heads_2 <= _heads_T_12;
        end
      end
    end
    if (reset) begin // @[InputUnit.scala 87:24]
      tails_0 <= 4'h0; // @[InputUnit.scala 87:24]
    end else if (io_enq_0_valid & ~direct_to_q) begin // @[InputUnit.scala 100:44]
      if (2'h0 == io_enq_0_bits_virt_channel_id) begin // @[InputUnit.scala 103:45]
        if (_tails_T_8) begin // @[InputUnit.scala 103:51]
          tails_0 <= {{1'd0}, _tails_T_16};
        end else begin
          tails_0 <= _tails_T_18;
        end
      end
    end
    if (reset) begin // @[InputUnit.scala 87:24]
      tails_1 <= 4'h3; // @[InputUnit.scala 87:24]
    end else if (io_enq_0_valid & ~direct_to_q) begin // @[InputUnit.scala 100:44]
      if (2'h1 == io_enq_0_bits_virt_channel_id) begin // @[InputUnit.scala 103:45]
        if (_tails_T_8) begin // @[InputUnit.scala 103:51]
          tails_1 <= {{1'd0}, _tails_T_16};
        end else begin
          tails_1 <= _tails_T_18;
        end
      end
    end
    if (reset) begin // @[InputUnit.scala 87:24]
      tails_2 <= 4'h6; // @[InputUnit.scala 87:24]
    end else if (io_enq_0_valid & ~direct_to_q) begin // @[InputUnit.scala 100:44]
      if (2'h2 == io_enq_0_bits_virt_channel_id) begin // @[InputUnit.scala 103:45]
        if (_tails_T_8) begin // @[InputUnit.scala 103:51]
          tails_2 <= {{1'd0}, _tails_T_16};
        end else begin
          tails_2 <= _tails_T_18;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {1{`RANDOM}};
  _RAND_2 = {1{`RANDOM}};
  _RAND_3 = {1{`RANDOM}};
  _RAND_5 = {1{`RANDOM}};
  _RAND_6 = {1{`RANDOM}};
  _RAND_7 = {1{`RANDOM}};
  _RAND_9 = {2{`RANDOM}};
  _RAND_10 = {2{`RANDOM}};
  _RAND_11 = {2{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 9; initvar = initvar+1)
    mem_head[initvar] = _RAND_0[0:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 9; initvar = initvar+1)
    mem_tail[initvar] = _RAND_4[0:0];
  _RAND_8 = {2{`RANDOM}};
  for (initvar = 0; initvar < 9; initvar = initvar+1)
    mem_payload[initvar] = _RAND_8[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  heads_0 = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  heads_1 = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  heads_2 = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  tails_0 = _RAND_15[3:0];
  _RAND_16 = {1{`RANDOM}};
  tails_1 = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  tails_2 = _RAND_17[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Arbiter(
  input        io_in_0_valid,
  output       io_in_1_ready,
  input        io_in_1_valid,
  output       io_in_2_ready,
  input        io_in_2_valid,
  output       io_out_valid,
  output [1:0] io_out_bits_src_virt_id
);
  wire [1:0] _GEN_0 = io_in_1_valid ? 2'h1 : 2'h2; // @[Arbiter.scala 135:13 138:26 139:17]
  wire  grant_2 = ~(io_in_0_valid | io_in_1_valid); // @[Arbiter.scala 45:78]
  assign io_in_1_ready = ~io_in_0_valid; // @[Arbiter.scala 45:78]
  assign io_in_2_ready = ~(io_in_0_valid | io_in_1_valid); // @[Arbiter.scala 45:78]
  assign io_out_valid = ~grant_2 | io_in_2_valid; // @[Arbiter.scala 147:31]
  assign io_out_bits_src_virt_id = io_in_0_valid ? 2'h0 : _GEN_0; // @[Arbiter.scala 138:26 140:19]
endmodule
module SwitchArbiter_1(
  input        clock,
  input        reset,
  output       io_in_0_ready,
  input        io_in_0_valid,
  input        io_in_0_bits_vc_sel_0_0,
  input        io_in_0_bits_tail,
  output       io_in_1_ready,
  input        io_in_1_valid,
  input        io_in_1_bits_vc_sel_0_0,
  input        io_in_1_bits_tail,
  output       io_in_2_ready,
  input        io_in_2_valid,
  input        io_in_2_bits_vc_sel_0_0,
  input        io_in_2_bits_tail,
  input        io_out_0_ready,
  output       io_out_0_valid,
  output       io_out_0_bits_vc_sel_0_0,
  output       io_out_0_bits_tail,
  output [2:0] io_chosen_oh_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] lock_0; // @[SwitchAllocator.scala 24:38]
  wire [2:0] _unassigned_T = {io_in_2_valid,io_in_1_valid,io_in_0_valid}; // @[Cat.scala 33:92]
  wire [2:0] _unassigned_T_1 = ~lock_0; // @[SwitchAllocator.scala 25:54]
  wire [2:0] unassigned = _unassigned_T & _unassigned_T_1; // @[SwitchAllocator.scala 25:52]
  reg [2:0] mask; // @[SwitchAllocator.scala 27:21]
  wire [2:0] _GEN_5 = {{2'd0}, mask == 3'h0}; // @[SwitchAllocator.scala 30:58]
  wire [2:0] _sel_T_1 = unassigned & _GEN_5; // @[SwitchAllocator.scala 30:58]
  wire [5:0] _sel_T_2 = {unassigned,_sel_T_1}; // @[Cat.scala 33:92]
  wire [5:0] _sel_T_9 = _sel_T_2[5] ? 6'h20 : 6'h0; // @[Mux.scala 47:70]
  wire [5:0] _sel_T_10 = _sel_T_2[4] ? 6'h10 : _sel_T_9; // @[Mux.scala 47:70]
  wire [5:0] _sel_T_11 = _sel_T_2[3] ? 6'h8 : _sel_T_10; // @[Mux.scala 47:70]
  wire [5:0] _sel_T_12 = _sel_T_2[2] ? 6'h4 : _sel_T_11; // @[Mux.scala 47:70]
  wire [5:0] _sel_T_13 = _sel_T_2[1] ? 6'h2 : _sel_T_12; // @[Mux.scala 47:70]
  wire [5:0] sel = _sel_T_2[0] ? 6'h1 : _sel_T_13; // @[Mux.scala 47:70]
  wire [5:0] _GEN_6 = {{3'd0}, sel[5:3]}; // @[SwitchAllocator.scala 32:23]
  wire [5:0] _choices_0_T_1 = sel | _GEN_6; // @[SwitchAllocator.scala 32:23]
  wire [2:0] choices_0 = _choices_0_T_1[2:0]; // @[SwitchAllocator.scala 28:21 32:16]
  wire [2:0] in_tails = {io_in_2_bits_tail,io_in_1_bits_tail,io_in_0_bits_tail}; // @[Cat.scala 33:92]
  wire [2:0] _chosen_T = _unassigned_T & lock_0; // @[SwitchAllocator.scala 42:33]
  wire [2:0] chosen = |_chosen_T ? lock_0 : choices_0; // @[SwitchAllocator.scala 42:21]
  wire [2:0] _io_out_0_valid_T = _unassigned_T & chosen; // @[SwitchAllocator.scala 44:35]
  wire  _T_13 = io_out_0_ready & io_out_0_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _lock_0_T = ~in_tails; // @[SwitchAllocator.scala 53:27]
  wire [2:0] _lock_0_T_1 = chosen & _lock_0_T; // @[SwitchAllocator.scala 53:25]
  wire [2:0] _GEN_7 = {{1'd0}, io_chosen_oh_0[2:1]}; // @[SwitchAllocator.scala 58:71]
  wire [2:0] _mask_T_3 = io_chosen_oh_0 | _GEN_7; // @[SwitchAllocator.scala 58:71]
  wire [2:0] _GEN_8 = {{2'd0}, io_chosen_oh_0[2]}; // @[SwitchAllocator.scala 58:71]
  wire [2:0] _mask_T_4 = _mask_T_3 | _GEN_8; // @[SwitchAllocator.scala 58:71]
  wire [2:0] _mask_T_5 = ~mask; // @[SwitchAllocator.scala 60:17]
  wire [3:0] _mask_T_7 = {mask, 1'h0}; // @[SwitchAllocator.scala 60:43]
  wire [3:0] _mask_T_8 = _mask_T_7 | 4'h1; // @[SwitchAllocator.scala 60:49]
  wire [3:0] _mask_T_9 = _mask_T_5 == 3'h0 ? 4'h0 : _mask_T_8; // @[SwitchAllocator.scala 60:16]
  wire [3:0] _GEN_4 = _T_13 ? {{1'd0}, _mask_T_4} : _mask_T_9; // @[SwitchAllocator.scala 57:27 58:10 60:10]
  wire [3:0] _GEN_9 = reset ? 4'h0 : _GEN_4; // @[SwitchAllocator.scala 27:{21,21}]
  assign io_in_0_ready = chosen[0] & io_out_0_ready; // @[SwitchAllocator.scala 47:23]
  assign io_in_1_ready = chosen[1] & io_out_0_ready; // @[SwitchAllocator.scala 47:23]
  assign io_in_2_ready = chosen[2] & io_out_0_ready; // @[SwitchAllocator.scala 47:23]
  assign io_out_0_valid = |_io_out_0_valid_T; // @[SwitchAllocator.scala 44:45]
  assign io_out_0_bits_vc_sel_0_0 = chosen[0] & io_in_0_bits_vc_sel_0_0 | chosen[1] & io_in_1_bits_vc_sel_0_0 | chosen[2
    ] & io_in_2_bits_vc_sel_0_0; // @[Mux.scala 27:73]
  assign io_out_0_bits_tail = chosen[0] & io_in_0_bits_tail | chosen[1] & io_in_1_bits_tail | chosen[2] &
    io_in_2_bits_tail; // @[Mux.scala 27:73]
  assign io_chosen_oh_0 = |_chosen_T ? lock_0 : choices_0; // @[SwitchAllocator.scala 42:21]
  always @(posedge clock) begin
    if (reset) begin // @[SwitchAllocator.scala 24:38]
      lock_0 <= 3'h0; // @[SwitchAllocator.scala 24:38]
    end else if (_T_13) begin // @[SwitchAllocator.scala 52:29]
      lock_0 <= _lock_0_T_1; // @[SwitchAllocator.scala 53:15]
    end
    mask <= _GEN_9[2:0]; // @[SwitchAllocator.scala 27:{21,21}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lock_0 = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  mask = _RAND_1[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module InputUnit(
  input         clock,
  input         reset,
  output        io_router_req_valid,
  output [1:0]  io_router_req_bits_src_virt_id,
  input         io_vcalloc_req_ready,
  output        io_vcalloc_req_valid,
  output        io_vcalloc_req_bits_vc_sel_0_0,
  input         io_vcalloc_resp_vc_sel_0_0,
  input         io_out_credit_available_0_0,
  input         io_salloc_req_0_ready,
  output        io_salloc_req_0_valid,
  output        io_salloc_req_0_bits_vc_sel_0_0,
  output        io_salloc_req_0_bits_tail,
  output        io_out_0_valid,
  output        io_out_0_bits_flit_head,
  output        io_out_0_bits_flit_tail,
  output [63:0] io_out_0_bits_flit_payload,
  output [1:0]  io_debug_va_stall,
  output [1:0]  io_debug_sa_stall,
  input         io_in_flit_0_valid,
  input         io_in_flit_0_bits_head,
  input         io_in_flit_0_bits_tail,
  input  [63:0] io_in_flit_0_bits_payload,
  input         io_in_flit_0_bits_flow_egress_node,
  input  [1:0]  io_in_flit_0_bits_virt_channel_id,
  output [2:0]  io_in_credit_return,
  output [2:0]  io_in_vc_free
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire  input_buffer_clock; // @[InputUnit.scala 180:28]
  wire  input_buffer_reset; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_enq_0_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_enq_0_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_enq_0_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_enq_0_bits_payload; // @[InputUnit.scala 180:28]
  wire [1:0] input_buffer_io_enq_0_bits_virt_channel_id; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_0_ready; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_0_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_0_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_0_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_deq_0_bits_payload; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_ready; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_deq_1_bits_payload; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_ready; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_deq_2_bits_payload; // @[InputUnit.scala 180:28]
  wire  route_arbiter_io_in_0_valid; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_1_ready; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_1_valid; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_2_ready; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_2_valid; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_out_valid; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_out_bits_src_virt_id; // @[InputUnit.scala 186:29]
  wire  salloc_arb_clock; // @[InputUnit.scala 279:26]
  wire  salloc_arb_reset; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_bits_tail; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_tail; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_tail; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_tail; // @[InputUnit.scala 279:26]
  wire [2:0] salloc_arb_io_chosen_oh_0; // @[InputUnit.scala 279:26]
  reg [2:0] states_0_g; // @[InputUnit.scala 191:19]
  reg  states_0_vc_sel_0_0; // @[InputUnit.scala 191:19]
  reg [2:0] states_1_g; // @[InputUnit.scala 191:19]
  reg  states_1_vc_sel_0_0; // @[InputUnit.scala 191:19]
  reg [2:0] states_2_g; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_0_0; // @[InputUnit.scala 191:19]
  wire  _T = io_in_flit_0_valid & io_in_flit_0_bits_head; // @[InputUnit.scala 194:32]
  wire  _T_3 = ~reset; // @[InputUnit.scala 196:13]
  wire [2:0] _GEN_1 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? states_1_g : states_0_g; // @[InputUnit.scala 197:{27,27}]
  wire [2:0] _GEN_2 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? states_2_g : _GEN_1; // @[InputUnit.scala 197:{27,27}]
  wire [2:0] _states_g_T = io_in_flit_0_bits_flow_egress_node ? 3'h2 : 3'h1; // @[InputUnit.scala 199:26]
  wire [2:0] _GEN_3 = 2'h0 == io_in_flit_0_bits_virt_channel_id ? _states_g_T : states_0_g; // @[InputUnit.scala 191:19 199:{20,20}]
  wire [2:0] _GEN_4 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? _states_g_T : states_1_g; // @[InputUnit.scala 191:19 199:{20,20}]
  wire [2:0] _GEN_5 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? _states_g_T : states_2_g; // @[InputUnit.scala 191:19 199:{20,20}]
  wire  _GEN_6 = 2'h0 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_0_vc_sel_0_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_7 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_1_vc_sel_0_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_8 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_0_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_9 = 2'h0 == io_in_flit_0_bits_virt_channel_id | _GEN_6; // @[InputUnit.scala 203:{44,44}]
  wire  _GEN_10 = 2'h1 == io_in_flit_0_bits_virt_channel_id | _GEN_7; // @[InputUnit.scala 203:{44,44}]
  wire  _GEN_11 = 2'h2 == io_in_flit_0_bits_virt_channel_id | _GEN_8; // @[InputUnit.scala 203:{44,44}]
  wire [2:0] _GEN_30 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_3 : states_0_g; // @[InputUnit.scala 191:19 194:60]
  wire [2:0] _GEN_31 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_4 : states_1_g; // @[InputUnit.scala 191:19 194:60]
  wire [2:0] _GEN_32 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_5 : states_2_g; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_33 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_9 : states_0_vc_sel_0_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_34 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_10 : states_1_vc_sel_0_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_35 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_11 : states_2_vc_sel_0_0; // @[InputUnit.scala 191:19 194:60]
  wire  _T_10 = route_arbiter_io_in_0_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_51 = _T_10 ? 3'h2 : _GEN_30; // @[InputUnit.scala 215:{23,29}]
  wire  _T_11 = route_arbiter_io_in_1_ready & route_arbiter_io_in_1_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_52 = _T_11 ? 3'h2 : _GEN_31; // @[InputUnit.scala 215:{23,29}]
  wire  _T_12 = route_arbiter_io_in_2_ready & route_arbiter_io_in_2_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_53 = _T_12 ? 3'h2 : _GEN_32; // @[InputUnit.scala 215:{23,29}]
  wire [2:0] _GEN_55 = 2'h1 == io_router_req_bits_src_virt_id ? states_1_g : states_0_g; // @[InputUnit.scala 224:{25,25}]
  wire [2:0] _GEN_56 = 2'h2 == io_router_req_bits_src_virt_id ? states_2_g : _GEN_55; // @[InputUnit.scala 224:{25,25}]
  wire [2:0] _GEN_57 = 2'h0 == io_router_req_bits_src_virt_id ? 3'h2 : _GEN_51; // @[InputUnit.scala 225:{18,18}]
  wire [2:0] _GEN_58 = 2'h1 == io_router_req_bits_src_virt_id ? 3'h2 : _GEN_52; // @[InputUnit.scala 225:{18,18}]
  wire [2:0] _GEN_59 = 2'h2 == io_router_req_bits_src_virt_id ? 3'h2 : _GEN_53; // @[InputUnit.scala 225:{18,18}]
  wire  _GEN_60 = 2'h0 == io_router_req_bits_src_virt_id ? 1'h0 : _GEN_33; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_61 = 2'h1 == io_router_req_bits_src_virt_id ? 1'h0 : _GEN_34; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_62 = 2'h2 == io_router_req_bits_src_virt_id ? 1'h0 : _GEN_35; // @[InputUnit.scala 227:25 228:26]
  wire [2:0] _GEN_63 = io_router_req_valid ? _GEN_57 : _GEN_51; // @[InputUnit.scala 222:31]
  wire [2:0] _GEN_64 = io_router_req_valid ? _GEN_58 : _GEN_52; // @[InputUnit.scala 222:31]
  wire [2:0] _GEN_65 = io_router_req_valid ? _GEN_59 : _GEN_53; // @[InputUnit.scala 222:31]
  wire  _GEN_66 = io_router_req_valid ? _GEN_60 : _GEN_33; // @[InputUnit.scala 222:31]
  wire  _GEN_67 = io_router_req_valid ? _GEN_61 : _GEN_34; // @[InputUnit.scala 222:31]
  wire  _GEN_68 = io_router_req_valid ? _GEN_62 : _GEN_35; // @[InputUnit.scala 222:31]
  reg [2:0] mask; // @[InputUnit.scala 233:21]
  wire  vcalloc_vals_2 = states_2_g == 3'h2; // @[InputUnit.scala 249:32]
  wire  vcalloc_vals_1 = states_1_g == 3'h2; // @[InputUnit.scala 249:32]
  wire  vcalloc_vals_0 = states_0_g == 3'h2; // @[InputUnit.scala 249:32]
  wire [2:0] _vcalloc_filter_T = {vcalloc_vals_2,vcalloc_vals_1,vcalloc_vals_0}; // @[InputUnit.scala 236:59]
  wire [2:0] _vcalloc_filter_T_2 = ~mask; // @[InputUnit.scala 236:89]
  wire [2:0] _vcalloc_filter_T_3 = _vcalloc_filter_T & _vcalloc_filter_T_2; // @[InputUnit.scala 236:87]
  wire [5:0] _vcalloc_filter_T_4 = {vcalloc_vals_2,vcalloc_vals_1,vcalloc_vals_0,_vcalloc_filter_T_3}; // @[Cat.scala 33:92]
  wire [5:0] _vcalloc_filter_T_11 = _vcalloc_filter_T_4[5] ? 6'h20 : 6'h0; // @[Mux.scala 47:70]
  wire [5:0] _vcalloc_filter_T_12 = _vcalloc_filter_T_4[4] ? 6'h10 : _vcalloc_filter_T_11; // @[Mux.scala 47:70]
  wire [5:0] _vcalloc_filter_T_13 = _vcalloc_filter_T_4[3] ? 6'h8 : _vcalloc_filter_T_12; // @[Mux.scala 47:70]
  wire [5:0] _vcalloc_filter_T_14 = _vcalloc_filter_T_4[2] ? 6'h4 : _vcalloc_filter_T_13; // @[Mux.scala 47:70]
  wire [5:0] _vcalloc_filter_T_15 = _vcalloc_filter_T_4[1] ? 6'h2 : _vcalloc_filter_T_14; // @[Mux.scala 47:70]
  wire [5:0] vcalloc_filter = _vcalloc_filter_T_4[0] ? 6'h1 : _vcalloc_filter_T_15; // @[Mux.scala 47:70]
  wire [2:0] vcalloc_sel = vcalloc_filter[2:0] | vcalloc_filter[5:3]; // @[InputUnit.scala 237:58]
  wire [3:0] _mask_T = 4'h1 << io_router_req_bits_src_virt_id; // @[InputUnit.scala 240:18]
  wire [3:0] _mask_T_2 = _mask_T - 4'h1; // @[InputUnit.scala 240:53]
  wire  _T_23 = vcalloc_vals_0 | vcalloc_vals_1 | vcalloc_vals_2; // @[package.scala 73:59]
  wire [1:0] _mask_T_10 = vcalloc_sel[1] ? 2'h3 : 2'h0; // @[Mux.scala 27:73]
  wire [2:0] _mask_T_11 = vcalloc_sel[2] ? 3'h7 : 3'h0; // @[Mux.scala 27:73]
  wire [1:0] _GEN_21 = {{1'd0}, vcalloc_sel[0]}; // @[Mux.scala 27:73]
  wire [1:0] _mask_T_12 = _GEN_21 | _mask_T_10; // @[Mux.scala 27:73]
  wire [2:0] _GEN_22 = {{1'd0}, _mask_T_12}; // @[Mux.scala 27:73]
  wire [2:0] _mask_T_13 = _GEN_22 | _mask_T_11; // @[Mux.scala 27:73]
  wire [2:0] _GEN_69 = _T_23 ? _mask_T_13 : mask; // @[InputUnit.scala 241:34 242:10 233:21]
  wire [3:0] _GEN_70 = io_router_req_valid ? _mask_T_2 : {{1'd0}, _GEN_69}; // @[InputUnit.scala 239:31 240:10]
  wire [2:0] _GEN_71 = vcalloc_vals_0 & vcalloc_sel[0] & io_vcalloc_req_ready ? 3'h3 : _GEN_63; // @[InputUnit.scala 253:{76,82}]
  wire [2:0] _GEN_72 = vcalloc_vals_1 & vcalloc_sel[1] & io_vcalloc_req_ready ? 3'h3 : _GEN_64; // @[InputUnit.scala 253:{76,82}]
  wire [2:0] _GEN_73 = vcalloc_vals_2 & vcalloc_sel[2] & io_vcalloc_req_ready ? 3'h3 : _GEN_65; // @[InputUnit.scala 253:{76,82}]
  wire [1:0] _io_debug_va_stall_T = vcalloc_vals_1 + vcalloc_vals_2; // @[Bitwise.scala 51:90]
  wire [1:0] _GEN_23 = {{1'd0}, vcalloc_vals_0}; // @[Bitwise.scala 51:90]
  wire [2:0] _io_debug_va_stall_T_2 = _GEN_23 + _io_debug_va_stall_T; // @[Bitwise.scala 51:90]
  wire [1:0] _GEN_27 = {{1'd0}, io_vcalloc_req_ready}; // @[InputUnit.scala 266:47]
  wire  _T_33 = io_vcalloc_req_ready & io_vcalloc_req_valid; // @[Decoupled.scala 51:35]
  wire  credit_available = states_0_vc_sel_0_0 & io_out_credit_available_0_0; // @[InputUnit.scala 287:47]
  wire  _T_49 = salloc_arb_io_in_0_ready & salloc_arb_io_in_0_valid; // @[Decoupled.scala 51:35]
  wire  credit_available_1 = states_1_vc_sel_0_0 & io_out_credit_available_0_0; // @[InputUnit.scala 287:47]
  wire  _T_51 = salloc_arb_io_in_1_ready & salloc_arb_io_in_1_valid; // @[Decoupled.scala 51:35]
  wire  credit_available_2 = states_2_vc_sel_0_0 & io_out_credit_available_0_0; // @[InputUnit.scala 287:47]
  wire  _T_53 = salloc_arb_io_in_2_ready & salloc_arb_io_in_2_valid; // @[Decoupled.scala 51:35]
  wire  _io_debug_sa_stall_T_1 = salloc_arb_io_in_0_valid & ~salloc_arb_io_in_0_ready; // @[InputUnit.scala 301:67]
  wire  _io_debug_sa_stall_T_3 = salloc_arb_io_in_1_valid & ~salloc_arb_io_in_1_ready; // @[InputUnit.scala 301:67]
  wire  _io_debug_sa_stall_T_5 = salloc_arb_io_in_2_valid & ~salloc_arb_io_in_2_ready; // @[InputUnit.scala 301:67]
  wire [1:0] _io_debug_sa_stall_T_6 = _io_debug_sa_stall_T_3 + _io_debug_sa_stall_T_5; // @[Bitwise.scala 51:90]
  wire [1:0] _GEN_28 = {{1'd0}, _io_debug_sa_stall_T_1}; // @[Bitwise.scala 51:90]
  wire [2:0] _io_debug_sa_stall_T_8 = _GEN_28 + _io_debug_sa_stall_T_6; // @[Bitwise.scala 51:90]
  reg  salloc_outs_0_valid; // @[InputUnit.scala 318:8]
  reg  salloc_outs_0_flit_head; // @[InputUnit.scala 318:8]
  reg  salloc_outs_0_flit_tail; // @[InputUnit.scala 318:8]
  reg [63:0] salloc_outs_0_flit_payload; // @[InputUnit.scala 318:8]
  wire  _io_in_credit_return_T = salloc_arb_io_out_0_ready & salloc_arb_io_out_0_valid; // @[Decoupled.scala 51:35]
  wire  _io_in_vc_free_T_8 = salloc_arb_io_chosen_oh_0[0] & input_buffer_io_deq_0_bits_tail | salloc_arb_io_chosen_oh_0[
    1] & input_buffer_io_deq_1_bits_tail | salloc_arb_io_chosen_oh_0[2] & input_buffer_io_deq_2_bits_tail; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_3 = salloc_arb_io_chosen_oh_0[0] ? input_buffer_io_deq_0_bits_payload : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_4 = salloc_arb_io_chosen_oh_0[1] ? input_buffer_io_deq_1_bits_payload : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_5 = salloc_arb_io_chosen_oh_0[2] ? input_buffer_io_deq_2_bits_payload : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_6 = _salloc_outs_0_flit_payload_T_3 | _salloc_outs_0_flit_payload_T_4; // @[Mux.scala 27:73]
  wire [3:0] _GEN_36 = reset ? 4'h0 : _GEN_70; // @[InputUnit.scala 233:{21,21}]
  wire  _GEN_37 = _T & ~reset; // @[InputUnit.scala 196:13]
  InputBuffer input_buffer ( // @[InputUnit.scala 180:28]
    .clock(input_buffer_clock),
    .reset(input_buffer_reset),
    .io_enq_0_valid(input_buffer_io_enq_0_valid),
    .io_enq_0_bits_head(input_buffer_io_enq_0_bits_head),
    .io_enq_0_bits_tail(input_buffer_io_enq_0_bits_tail),
    .io_enq_0_bits_payload(input_buffer_io_enq_0_bits_payload),
    .io_enq_0_bits_virt_channel_id(input_buffer_io_enq_0_bits_virt_channel_id),
    .io_deq_0_ready(input_buffer_io_deq_0_ready),
    .io_deq_0_valid(input_buffer_io_deq_0_valid),
    .io_deq_0_bits_head(input_buffer_io_deq_0_bits_head),
    .io_deq_0_bits_tail(input_buffer_io_deq_0_bits_tail),
    .io_deq_0_bits_payload(input_buffer_io_deq_0_bits_payload),
    .io_deq_1_ready(input_buffer_io_deq_1_ready),
    .io_deq_1_valid(input_buffer_io_deq_1_valid),
    .io_deq_1_bits_head(input_buffer_io_deq_1_bits_head),
    .io_deq_1_bits_tail(input_buffer_io_deq_1_bits_tail),
    .io_deq_1_bits_payload(input_buffer_io_deq_1_bits_payload),
    .io_deq_2_ready(input_buffer_io_deq_2_ready),
    .io_deq_2_valid(input_buffer_io_deq_2_valid),
    .io_deq_2_bits_head(input_buffer_io_deq_2_bits_head),
    .io_deq_2_bits_tail(input_buffer_io_deq_2_bits_tail),
    .io_deq_2_bits_payload(input_buffer_io_deq_2_bits_payload)
  );
  Arbiter route_arbiter ( // @[InputUnit.scala 186:29]
    .io_in_0_valid(route_arbiter_io_in_0_valid),
    .io_in_1_ready(route_arbiter_io_in_1_ready),
    .io_in_1_valid(route_arbiter_io_in_1_valid),
    .io_in_2_ready(route_arbiter_io_in_2_ready),
    .io_in_2_valid(route_arbiter_io_in_2_valid),
    .io_out_valid(route_arbiter_io_out_valid),
    .io_out_bits_src_virt_id(route_arbiter_io_out_bits_src_virt_id)
  );
  SwitchArbiter_1 salloc_arb ( // @[InputUnit.scala 279:26]
    .clock(salloc_arb_clock),
    .reset(salloc_arb_reset),
    .io_in_0_ready(salloc_arb_io_in_0_ready),
    .io_in_0_valid(salloc_arb_io_in_0_valid),
    .io_in_0_bits_vc_sel_0_0(salloc_arb_io_in_0_bits_vc_sel_0_0),
    .io_in_0_bits_tail(salloc_arb_io_in_0_bits_tail),
    .io_in_1_ready(salloc_arb_io_in_1_ready),
    .io_in_1_valid(salloc_arb_io_in_1_valid),
    .io_in_1_bits_vc_sel_0_0(salloc_arb_io_in_1_bits_vc_sel_0_0),
    .io_in_1_bits_tail(salloc_arb_io_in_1_bits_tail),
    .io_in_2_ready(salloc_arb_io_in_2_ready),
    .io_in_2_valid(salloc_arb_io_in_2_valid),
    .io_in_2_bits_vc_sel_0_0(salloc_arb_io_in_2_bits_vc_sel_0_0),
    .io_in_2_bits_tail(salloc_arb_io_in_2_bits_tail),
    .io_out_0_ready(salloc_arb_io_out_0_ready),
    .io_out_0_valid(salloc_arb_io_out_0_valid),
    .io_out_0_bits_vc_sel_0_0(salloc_arb_io_out_0_bits_vc_sel_0_0),
    .io_out_0_bits_tail(salloc_arb_io_out_0_bits_tail),
    .io_chosen_oh_0(salloc_arb_io_chosen_oh_0)
  );
  assign io_router_req_valid = route_arbiter_io_out_valid; // @[InputUnit.scala 189:17]
  assign io_router_req_bits_src_virt_id = route_arbiter_io_out_bits_src_virt_id; // @[InputUnit.scala 189:17]
  assign io_vcalloc_req_valid = vcalloc_vals_0 | vcalloc_vals_1 | vcalloc_vals_2; // @[package.scala 73:59]
  assign io_vcalloc_req_bits_vc_sel_0_0 = vcalloc_sel[0] & states_0_vc_sel_0_0 | vcalloc_sel[1] & states_1_vc_sel_0_0 |
    vcalloc_sel[2] & states_2_vc_sel_0_0; // @[Mux.scala 27:73]
  assign io_salloc_req_0_valid = salloc_arb_io_out_0_valid; // @[InputUnit.scala 302:17 303:19 305:35]
  assign io_salloc_req_0_bits_vc_sel_0_0 = salloc_arb_io_out_0_bits_vc_sel_0_0; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_tail = salloc_arb_io_out_0_bits_tail; // @[InputUnit.scala 302:17]
  assign io_out_0_valid = salloc_outs_0_valid; // @[InputUnit.scala 349:21]
  assign io_out_0_bits_flit_head = salloc_outs_0_flit_head; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_flit_tail = salloc_outs_0_flit_tail; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_flit_payload = salloc_outs_0_flit_payload; // @[InputUnit.scala 350:25]
  assign io_debug_va_stall = _io_debug_va_stall_T_2[1:0] - _GEN_27; // @[InputUnit.scala 266:47]
  assign io_debug_sa_stall = _io_debug_sa_stall_T_8[1:0]; // @[Bitwise.scala 51:90]
  assign io_in_credit_return = _io_in_credit_return_T ? salloc_arb_io_chosen_oh_0 : 3'h0; // @[InputUnit.scala 322:8]
  assign io_in_vc_free = _io_in_credit_return_T & _io_in_vc_free_T_8 ? salloc_arb_io_chosen_oh_0 : 3'h0; // @[InputUnit.scala 325:8]
  assign input_buffer_clock = clock;
  assign input_buffer_reset = reset;
  assign input_buffer_io_enq_0_valid = io_in_flit_0_valid; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_head = io_in_flit_0_bits_head; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_tail = io_in_flit_0_bits_tail; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_payload = io_in_flit_0_bits_payload; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_virt_channel_id = io_in_flit_0_bits_virt_channel_id; // @[InputUnit.scala 182:28]
  assign input_buffer_io_deq_0_ready = salloc_arb_io_in_0_ready; // @[InputUnit.scala 295:36]
  assign input_buffer_io_deq_1_ready = salloc_arb_io_in_1_ready; // @[InputUnit.scala 295:36]
  assign input_buffer_io_deq_2_ready = salloc_arb_io_in_2_ready; // @[InputUnit.scala 295:36]
  assign route_arbiter_io_in_0_valid = states_0_g == 3'h1; // @[InputUnit.scala 212:22]
  assign route_arbiter_io_in_1_valid = states_1_g == 3'h1; // @[InputUnit.scala 212:22]
  assign route_arbiter_io_in_2_valid = states_2_g == 3'h1; // @[InputUnit.scala 212:22]
  assign salloc_arb_clock = clock;
  assign salloc_arb_reset = reset;
  assign salloc_arb_io_in_0_valid = states_0_g == 3'h3 & credit_available & input_buffer_io_deq_0_valid; // @[InputUnit.scala 288:50]
  assign salloc_arb_io_in_0_bits_vc_sel_0_0 = states_0_vc_sel_0_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_0_bits_tail = input_buffer_io_deq_0_bits_tail; // @[InputUnit.scala 291:19]
  assign salloc_arb_io_in_1_valid = states_1_g == 3'h3 & credit_available_1 & input_buffer_io_deq_1_valid; // @[InputUnit.scala 288:50]
  assign salloc_arb_io_in_1_bits_vc_sel_0_0 = states_1_vc_sel_0_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_1_bits_tail = input_buffer_io_deq_1_bits_tail; // @[InputUnit.scala 291:19]
  assign salloc_arb_io_in_2_valid = states_2_g == 3'h3 & credit_available_2 & input_buffer_io_deq_2_valid; // @[InputUnit.scala 288:50]
  assign salloc_arb_io_in_2_bits_vc_sel_0_0 = states_2_vc_sel_0_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_tail = input_buffer_io_deq_2_bits_tail; // @[InputUnit.scala 291:19]
  assign salloc_arb_io_out_0_ready = io_salloc_req_0_ready; // @[InputUnit.scala 302:17 303:19 304:39]
  always @(posedge clock) begin
    if (reset) begin // @[InputUnit.scala 377:23]
      states_0_g <= 3'h0; // @[InputUnit.scala 378:24]
    end else if (_T_49 & input_buffer_io_deq_0_bits_tail) begin // @[InputUnit.scala 292:35]
      states_0_g <= 3'h0; // @[InputUnit.scala 293:13]
    end else if (_T_33) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[0]) begin // @[InputUnit.scala 270:29]
        states_0_g <= 3'h3; // @[InputUnit.scala 272:21]
      end else begin
        states_0_g <= _GEN_71;
      end
    end else begin
      states_0_g <= _GEN_71;
    end
    if (_T_33) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[0]) begin // @[InputUnit.scala 270:29]
        states_0_vc_sel_0_0 <= io_vcalloc_resp_vc_sel_0_0; // @[InputUnit.scala 271:26]
      end else begin
        states_0_vc_sel_0_0 <= _GEN_66;
      end
    end else begin
      states_0_vc_sel_0_0 <= _GEN_66;
    end
    if (reset) begin // @[InputUnit.scala 377:23]
      states_1_g <= 3'h0; // @[InputUnit.scala 378:24]
    end else if (_T_51 & input_buffer_io_deq_1_bits_tail) begin // @[InputUnit.scala 292:35]
      states_1_g <= 3'h0; // @[InputUnit.scala 293:13]
    end else if (_T_33) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_g <= 3'h3; // @[InputUnit.scala 272:21]
      end else begin
        states_1_g <= _GEN_72;
      end
    end else begin
      states_1_g <= _GEN_72;
    end
    if (_T_33) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_vc_sel_0_0 <= io_vcalloc_resp_vc_sel_0_0; // @[InputUnit.scala 271:26]
      end else begin
        states_1_vc_sel_0_0 <= _GEN_67;
      end
    end else begin
      states_1_vc_sel_0_0 <= _GEN_67;
    end
    if (reset) begin // @[InputUnit.scala 377:23]
      states_2_g <= 3'h0; // @[InputUnit.scala 378:24]
    end else if (_T_53 & input_buffer_io_deq_2_bits_tail) begin // @[InputUnit.scala 292:35]
      states_2_g <= 3'h0; // @[InputUnit.scala 293:13]
    end else if (_T_33) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_g <= 3'h3; // @[InputUnit.scala 272:21]
      end else begin
        states_2_g <= _GEN_73;
      end
    end else begin
      states_2_g <= _GEN_73;
    end
    if (_T_33) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_0_0 <= io_vcalloc_resp_vc_sel_0_0; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_0_0 <= _GEN_68;
      end
    end else begin
      states_2_vc_sel_0_0 <= _GEN_68;
    end
    mask <= _GEN_36[2:0]; // @[InputUnit.scala 233:{21,21}]
    salloc_outs_0_valid <= salloc_arb_io_out_0_ready & salloc_arb_io_out_0_valid; // @[Decoupled.scala 51:35]
    salloc_outs_0_flit_head <= salloc_arb_io_chosen_oh_0[0] & input_buffer_io_deq_0_bits_head |
      salloc_arb_io_chosen_oh_0[1] & input_buffer_io_deq_1_bits_head | salloc_arb_io_chosen_oh_0[2] &
      input_buffer_io_deq_2_bits_head; // @[Mux.scala 27:73]
    salloc_outs_0_flit_tail <= salloc_arb_io_chosen_oh_0[0] & input_buffer_io_deq_0_bits_tail |
      salloc_arb_io_chosen_oh_0[1] & input_buffer_io_deq_1_bits_tail | salloc_arb_io_chosen_oh_0[2] &
      input_buffer_io_deq_2_bits_tail; // @[Mux.scala 27:73]
    salloc_outs_0_flit_payload <= _salloc_outs_0_flit_payload_T_6 | _salloc_outs_0_flit_payload_T_5; // @[Mux.scala 27:73]
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T & ~reset & ~(io_in_flit_0_bits_virt_channel_id < 2'h3)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:196 assert(id < nVirtualChannels.U)\n"); // @[InputUnit.scala 196:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_37 & ~(_GEN_2 == 3'h0)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:197 assert(states(id).g === g_i)\n"); // @[InputUnit.scala 197:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_router_req_valid & _T_3 & ~(_GEN_56 == 3'h1)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:224 assert(states(id).g === g_r)\n"); // @[InputUnit.scala 224:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_33 & vcalloc_sel[0] & _T_3 & ~vcalloc_vals_0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:274 assert(states(i).g === g_v)\n"); // @[InputUnit.scala 274:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_33 & vcalloc_sel[1] & _T_3 & ~vcalloc_vals_1) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:274 assert(states(i).g === g_v)\n"); // @[InputUnit.scala 274:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_33 & vcalloc_sel[2] & _T_3 & ~vcalloc_vals_2) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:274 assert(states(i).g === g_v)\n"); // @[InputUnit.scala 274:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  states_0_g = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  states_0_vc_sel_0_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  states_1_g = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  states_1_vc_sel_0_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  states_2_g = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  states_2_vc_sel_0_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  mask = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  salloc_outs_0_valid = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  salloc_outs_0_flit_head = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  salloc_outs_0_flit_tail = _RAND_9[0:0];
  _RAND_10 = {2{`RANDOM}};
  salloc_outs_0_flit_payload = _RAND_10[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (_T & ~reset) begin
      assert(io_in_flit_0_bits_virt_channel_id < 2'h3); // @[InputUnit.scala 196:13]
    end
    //
    if (_T & _T_3) begin
      assert(_GEN_2 == 3'h0); // @[InputUnit.scala 197:13]
    end
    //
    if (io_router_req_valid & _T_3) begin
      assert(_GEN_56 == 3'h1); // @[InputUnit.scala 224:11]
    end
    //
    if (_T_33 & vcalloc_sel[0] & _T_3) begin
      assert(vcalloc_vals_0); // @[InputUnit.scala 274:17]
    end
    //
    if (_T_33 & vcalloc_sel[1] & _T_3) begin
      assert(vcalloc_vals_1); // @[InputUnit.scala 274:17]
    end
    //
    if (_T_33 & vcalloc_sel[2] & _T_3) begin
      assert(vcalloc_vals_2); // @[InputUnit.scala 274:17]
    end
  end
endmodule
module Queue_7(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_head,
  input         io_enq_bits_tail,
  input  [63:0] io_enq_bits_payload,
  output        io_deq_valid,
  output        io_deq_bits_head,
  output        io_deq_bits_tail,
  output [63:0] io_deq_bits_payload,
  output        io_deq_bits_ingress_id,
  output [1:0]  io_count
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg  ram_head [0:2]; // @[Decoupled.scala 273:95]
  wire  ram_head_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [1:0] ram_head_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_head_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_head_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_tail [0:2]; // @[Decoupled.scala 273:95]
  wire  ram_tail_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [1:0] ram_tail_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_tail_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_tail_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_en; // @[Decoupled.scala 273:95]
  reg [63:0] ram_payload [0:2]; // @[Decoupled.scala 273:95]
  wire  ram_payload_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [1:0] ram_payload_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [63:0] ram_payload_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [63:0] ram_payload_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_payload_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_payload_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_payload_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_ingress_id [0:2]; // @[Decoupled.scala 273:95]
  wire  ram_ingress_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [1:0] ram_ingress_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_ingress_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_ingress_id_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_ingress_id_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_ingress_id_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_ingress_id_MPORT_en; // @[Decoupled.scala 273:95]
  reg [1:0] enq_ptr_value; // @[Counter.scala 61:40]
  reg [1:0] deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  wrap = enq_ptr_value == 2'h2; // @[Counter.scala 73:24]
  wire [1:0] _value_T_1 = enq_ptr_value + 2'h1; // @[Counter.scala 77:24]
  wire  do_enq = empty ? 1'h0 : _do_enq_T; // @[Decoupled.scala 315:17 280:27]
  wire  wrap_1 = deq_ptr_value == 2'h2; // @[Counter.scala 73:24]
  wire [1:0] _value_T_3 = deq_ptr_value + 2'h1; // @[Counter.scala 77:24]
  wire  do_deq = empty ? 1'h0 : io_deq_valid; // @[Decoupled.scala 315:17 317:14 281:27]
  wire [1:0] ptr_diff = enq_ptr_value - deq_ptr_value; // @[Decoupled.scala 326:32]
  wire [1:0] _io_count_T = maybe_full ? 2'h3 : 2'h0; // @[Decoupled.scala 333:10]
  wire [1:0] _io_count_T_3 = 2'h3 + ptr_diff; // @[Decoupled.scala 334:57]
  wire [1:0] _io_count_T_4 = deq_ptr_value > enq_ptr_value ? _io_count_T_3 : ptr_diff; // @[Decoupled.scala 334:10]
  assign ram_head_io_deq_bits_MPORT_en = 1'h1;
  assign ram_head_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_head_io_deq_bits_MPORT_data = ram_head[ram_head_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  `else
  assign ram_head_io_deq_bits_MPORT_data = ram_head_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_1[0:0] :
    ram_head[ram_head_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_head_MPORT_data = io_enq_bits_head;
  assign ram_head_MPORT_addr = enq_ptr_value;
  assign ram_head_MPORT_mask = 1'h1;
  assign ram_head_MPORT_en = empty ? 1'h0 : _do_enq_T;
  assign ram_tail_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tail_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_tail_io_deq_bits_MPORT_data = ram_tail[ram_tail_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  `else
  assign ram_tail_io_deq_bits_MPORT_data = ram_tail_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_3[0:0] :
    ram_tail[ram_tail_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_tail_MPORT_data = io_enq_bits_tail;
  assign ram_tail_MPORT_addr = enq_ptr_value;
  assign ram_tail_MPORT_mask = 1'h1;
  assign ram_tail_MPORT_en = empty ? 1'h0 : _do_enq_T;
  assign ram_payload_io_deq_bits_MPORT_en = 1'h1;
  assign ram_payload_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_payload_io_deq_bits_MPORT_data = ram_payload[ram_payload_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  `else
  assign ram_payload_io_deq_bits_MPORT_data = ram_payload_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_5[63:0] :
    ram_payload[ram_payload_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_payload_MPORT_data = io_enq_bits_payload;
  assign ram_payload_MPORT_addr = enq_ptr_value;
  assign ram_payload_MPORT_mask = 1'h1;
  assign ram_payload_MPORT_en = empty ? 1'h0 : _do_enq_T;
  assign ram_ingress_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_ingress_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_ingress_id_io_deq_bits_MPORT_data = ram_ingress_id[ram_ingress_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  `else
  assign ram_ingress_id_io_deq_bits_MPORT_data = ram_ingress_id_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_7[0:0] :
    ram_ingress_id[ram_ingress_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_ingress_id_MPORT_data = 1'h0;
  assign ram_ingress_id_MPORT_addr = enq_ptr_value;
  assign ram_ingress_id_MPORT_mask = 1'h1;
  assign ram_ingress_id_MPORT_en = empty ? 1'h0 : _do_enq_T;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 302:16 314:{24,39}]
  assign io_deq_bits_head = empty ? io_enq_bits_head : ram_head_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_tail = empty ? io_enq_bits_tail : ram_tail_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_payload = empty ? io_enq_bits_payload : ram_payload_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_ingress_id = empty ? 1'h0 : ram_ingress_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_count = ptr_match ? _io_count_T : _io_count_T_4; // @[Decoupled.scala 331:20]
  always @(posedge clock) begin
    if (ram_head_MPORT_en & ram_head_MPORT_mask) begin
      ram_head[ram_head_MPORT_addr] <= ram_head_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_tail_MPORT_en & ram_tail_MPORT_mask) begin
      ram_tail[ram_tail_MPORT_addr] <= ram_tail_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_payload_MPORT_en & ram_payload_MPORT_mask) begin
      ram_payload[ram_payload_MPORT_addr] <= ram_payload_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_ingress_id_MPORT_en & ram_ingress_id_MPORT_mask) begin
      ram_ingress_id[ram_ingress_id_MPORT_addr] <= ram_ingress_id_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 2'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      if (wrap) begin // @[Counter.scala 87:20]
        enq_ptr_value <= 2'h0; // @[Counter.scala 87:28]
      end else begin
        enq_ptr_value <= _value_T_1; // @[Counter.scala 77:15]
      end
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 2'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      if (wrap_1) begin // @[Counter.scala 87:20]
        deq_ptr_value <= 2'h0; // @[Counter.scala 87:28]
      end else begin
        deq_ptr_value <= _value_T_3; // @[Counter.scala 77:15]
      end
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      if (empty) begin // @[Decoupled.scala 315:17]
        maybe_full <= 1'h0;
      end else begin
        maybe_full <= _do_enq_T; // @[Decoupled.scala 280:27]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {1{`RANDOM}};
  _RAND_3 = {1{`RANDOM}};
  _RAND_5 = {2{`RANDOM}};
  _RAND_7 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_head[initvar] = _RAND_0[0:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_tail[initvar] = _RAND_2[0:0];
  _RAND_4 = {2{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_payload[initvar] = _RAND_4[63:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_ingress_id[initvar] = _RAND_6[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  enq_ptr_value = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  deq_ptr_value = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  maybe_full = _RAND_10[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module EgressUnit(
  input         clock,
  input         reset,
  input         io_in_0_valid,
  input         io_in_0_bits_head,
  input         io_in_0_bits_tail,
  input  [63:0] io_in_0_bits_payload,
  output        io_credit_available_0,
  output        io_channel_status_0_occupied,
  input         io_allocs_0_alloc,
  input         io_credit_alloc_0_alloc,
  input         io_credit_alloc_0_tail,
  output        io_out_valid,
  output        io_out_bits_head,
  output        io_out_bits_tail,
  output [63:0] io_out_bits_payload,
  output        io_out_bits_ingress_id
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  q_clock; // @[EgressUnit.scala 22:17]
  wire  q_reset; // @[EgressUnit.scala 22:17]
  wire  q_io_enq_ready; // @[EgressUnit.scala 22:17]
  wire  q_io_enq_valid; // @[EgressUnit.scala 22:17]
  wire  q_io_enq_bits_head; // @[EgressUnit.scala 22:17]
  wire  q_io_enq_bits_tail; // @[EgressUnit.scala 22:17]
  wire [63:0] q_io_enq_bits_payload; // @[EgressUnit.scala 22:17]
  wire  q_io_deq_valid; // @[EgressUnit.scala 22:17]
  wire  q_io_deq_bits_head; // @[EgressUnit.scala 22:17]
  wire  q_io_deq_bits_tail; // @[EgressUnit.scala 22:17]
  wire [63:0] q_io_deq_bits_payload; // @[EgressUnit.scala 22:17]
  wire  q_io_deq_bits_ingress_id; // @[EgressUnit.scala 22:17]
  wire [1:0] q_io_count; // @[EgressUnit.scala 22:17]
  reg  channel_empty; // @[EgressUnit.scala 20:30]
  wire  _GEN_0 = io_credit_alloc_0_alloc & io_credit_alloc_0_tail | channel_empty; // @[EgressUnit.scala 44:62 45:19 20:30]
  wire  _GEN_1 = io_allocs_0_alloc ? 1'h0 : _GEN_0; // @[EgressUnit.scala 49:29 50:19]
  Queue_7 q ( // @[EgressUnit.scala 22:17]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_head(q_io_enq_bits_head),
    .io_enq_bits_tail(q_io_enq_bits_tail),
    .io_enq_bits_payload(q_io_enq_bits_payload),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_head(q_io_deq_bits_head),
    .io_deq_bits_tail(q_io_deq_bits_tail),
    .io_deq_bits_payload(q_io_deq_bits_payload),
    .io_deq_bits_ingress_id(q_io_deq_bits_ingress_id),
    .io_count(q_io_count)
  );
  assign io_credit_available_0 = q_io_count == 2'h0; // @[EgressUnit.scala 40:40]
  assign io_channel_status_0_occupied = ~channel_empty; // @[EgressUnit.scala 41:36]
  assign io_out_valid = q_io_deq_valid; // @[EgressUnit.scala 37:10]
  assign io_out_bits_head = q_io_deq_bits_head; // @[EgressUnit.scala 37:10]
  assign io_out_bits_tail = q_io_deq_bits_tail; // @[EgressUnit.scala 37:10]
  assign io_out_bits_payload = q_io_deq_bits_payload; // @[EgressUnit.scala 37:10]
  assign io_out_bits_ingress_id = q_io_deq_bits_ingress_id; // @[EgressUnit.scala 37:10]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_in_0_valid; // @[EgressUnit.scala 23:18]
  assign q_io_enq_bits_head = io_in_0_bits_head; // @[EgressUnit.scala 24:22]
  assign q_io_enq_bits_tail = io_in_0_bits_tail; // @[EgressUnit.scala 25:22]
  assign q_io_enq_bits_payload = io_in_0_bits_payload; // @[EgressUnit.scala 36:25]
  always @(posedge clock) begin
    channel_empty <= reset | _GEN_1; // @[EgressUnit.scala 20:{30,30}]
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~(q_io_enq_valid & ~q_io_enq_ready))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at EgressUnit.scala:38 assert(!(q.io.enq.valid && !q.io.enq.ready))\n"); // @[EgressUnit.scala 38:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  channel_empty = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(~(q_io_enq_valid & ~q_io_enq_ready)); // @[EgressUnit.scala 38:9]
    end
  end
endmodule
module Switch_1(
  input         clock,
  input         reset,
  input         io_in_0_0_valid,
  input         io_in_0_0_bits_flit_head,
  input         io_in_0_0_bits_flit_tail,
  input  [63:0] io_in_0_0_bits_flit_payload,
  output        io_out_0_0_valid,
  output        io_out_0_0_bits_head,
  output        io_out_0_0_bits_tail,
  output [63:0] io_out_0_0_bits_payload,
  input         io_sel_0_0_0_0
);
  assign io_out_0_0_valid = io_in_0_0_valid & io_sel_0_0_0_0; // @[Switch.scala 48:67]
  assign io_out_0_0_bits_head = io_in_0_0_bits_flit_head; // @[Switch.scala 36:21 40:18]
  assign io_out_0_0_bits_tail = io_in_0_0_bits_flit_tail; // @[Switch.scala 36:21 40:18]
  assign io_out_0_0_bits_payload = io_in_0_0_bits_flit_payload; // @[Switch.scala 36:21 40:18]
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(1'h1); // @[Switch.scala 47:13]
    end
  end
endmodule
module SwitchArbiter_2(
  input   clock,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input   io_in_0_bits_vc_sel_0_0,
  input   io_in_0_bits_tail,
  output  io_out_0_valid,
  output  io_out_0_bits_vc_sel_0_0,
  output  io_out_0_bits_tail,
  output  io_chosen_oh_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  lock_0; // @[SwitchAllocator.scala 24:38]
  wire  unassigned = io_in_0_valid & ~lock_0; // @[SwitchAllocator.scala 25:52]
  reg  mask; // @[SwitchAllocator.scala 27:21]
  wire  _sel_T = ~mask; // @[SwitchAllocator.scala 30:60]
  wire  _sel_T_1 = unassigned & ~mask; // @[SwitchAllocator.scala 30:58]
  wire [1:0] _sel_T_2 = {unassigned,_sel_T_1}; // @[Cat.scala 33:92]
  wire [1:0] _sel_T_5 = _sel_T_2[1] ? 2'h2 : 2'h0; // @[Mux.scala 47:70]
  wire [1:0] sel = _sel_T_2[0] ? 2'h1 : _sel_T_5; // @[Mux.scala 47:70]
  wire [1:0] _GEN_3 = {{1'd0}, sel[1]}; // @[SwitchAllocator.scala 32:23]
  wire [1:0] _choices_0_T_1 = sel | _GEN_3; // @[SwitchAllocator.scala 32:23]
  wire  choices_0 = _choices_0_T_1[0]; // @[SwitchAllocator.scala 28:21 32:16]
  wire  chosen = |(io_in_0_valid & lock_0) ? lock_0 : choices_0; // @[SwitchAllocator.scala 42:21]
  wire [1:0] _mask_T_3 = {mask, 1'h0}; // @[SwitchAllocator.scala 60:43]
  wire [1:0] _mask_T_4 = _mask_T_3 | 2'h1; // @[SwitchAllocator.scala 60:49]
  wire [1:0] _mask_T_5 = ~_sel_T ? 2'h0 : _mask_T_4; // @[SwitchAllocator.scala 60:16]
  wire [1:0] _GEN_2 = io_out_0_valid ? {{1'd0}, io_chosen_oh_0} : _mask_T_5; // @[SwitchAllocator.scala 57:27 58:10 60:10]
  wire [1:0] _GEN_4 = reset ? 2'h0 : _GEN_2; // @[SwitchAllocator.scala 27:{21,21}]
  assign io_in_0_ready = |(io_in_0_valid & lock_0) ? lock_0 : choices_0; // @[SwitchAllocator.scala 42:21]
  assign io_out_0_valid = |(io_in_0_valid & chosen); // @[SwitchAllocator.scala 44:45]
  assign io_out_0_bits_vc_sel_0_0 = io_in_0_bits_vc_sel_0_0; // @[SwitchAllocator.scala 45:20]
  assign io_out_0_bits_tail = io_in_0_bits_tail; // @[SwitchAllocator.scala 45:20]
  assign io_chosen_oh_0 = |(io_in_0_valid & lock_0) ? lock_0 : choices_0; // @[SwitchAllocator.scala 42:21]
  always @(posedge clock) begin
    if (reset) begin // @[SwitchAllocator.scala 24:38]
      lock_0 <= 1'h0; // @[SwitchAllocator.scala 24:38]
    end else if (io_out_0_valid) begin // @[SwitchAllocator.scala 52:29]
      lock_0 <= chosen & ~io_in_0_bits_tail; // @[SwitchAllocator.scala 53:15]
    end
    mask <= _GEN_4[0]; // @[SwitchAllocator.scala 27:{21,21}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lock_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  mask = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SwitchAllocator_1(
  input   clock,
  input   reset,
  output  io_req_0_0_ready,
  input   io_req_0_0_valid,
  input   io_req_0_0_bits_vc_sel_0_0,
  input   io_req_0_0_bits_tail,
  output  io_credit_alloc_0_0_alloc,
  output  io_credit_alloc_0_0_tail,
  output  io_switch_sel_0_0_0_0
);
  wire  arbs_0_clock; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_reset; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_0_ready; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_0_valid; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_0_bits_vc_sel_0_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_0_bits_tail; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_out_0_valid; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_out_0_bits_vc_sel_0_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_out_0_bits_tail; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_chosen_oh_0; // @[SwitchAllocator.scala 83:45]
  SwitchArbiter_2 arbs_0 ( // @[SwitchAllocator.scala 83:45]
    .clock(arbs_0_clock),
    .reset(arbs_0_reset),
    .io_in_0_ready(arbs_0_io_in_0_ready),
    .io_in_0_valid(arbs_0_io_in_0_valid),
    .io_in_0_bits_vc_sel_0_0(arbs_0_io_in_0_bits_vc_sel_0_0),
    .io_in_0_bits_tail(arbs_0_io_in_0_bits_tail),
    .io_out_0_valid(arbs_0_io_out_0_valid),
    .io_out_0_bits_vc_sel_0_0(arbs_0_io_out_0_bits_vc_sel_0_0),
    .io_out_0_bits_tail(arbs_0_io_out_0_bits_tail),
    .io_chosen_oh_0(arbs_0_io_chosen_oh_0)
  );
  assign io_req_0_0_ready = arbs_0_io_in_0_ready & arbs_0_io_in_0_valid; // @[Decoupled.scala 51:35]
  assign io_credit_alloc_0_0_alloc = arbs_0_io_out_0_valid & arbs_0_io_out_0_bits_vc_sel_0_0; // @[SwitchAllocator.scala 120:33]
  assign io_credit_alloc_0_0_tail = arbs_0_io_out_0_valid & arbs_0_io_out_0_bits_vc_sel_0_0 & arbs_0_io_out_0_bits_tail; // @[SwitchAllocator.scala 120:67 122:21 116:44]
  assign io_switch_sel_0_0_0_0 = arbs_0_io_in_0_valid & arbs_0_io_chosen_oh_0 & arbs_0_io_out_0_valid; // @[SwitchAllocator.scala 108:97]
  assign arbs_0_clock = clock;
  assign arbs_0_reset = reset;
  assign arbs_0_io_in_0_valid = io_req_0_0_valid & io_req_0_0_bits_vc_sel_0_0; // @[SwitchAllocator.scala 95:37]
  assign arbs_0_io_in_0_bits_vc_sel_0_0 = io_req_0_0_bits_vc_sel_0_0; // @[SwitchAllocator.scala 96:25]
  assign arbs_0_io_in_0_bits_tail = io_req_0_0_bits_tail; // @[SwitchAllocator.scala 96:25]
endmodule
module RotatingSingleVCAllocator_1(
  input   clock,
  input   reset,
  output  io_req_0_ready,
  input   io_req_0_valid,
  input   io_req_0_bits_vc_sel_0_0,
  output  io_resp_0_vc_sel_0_0,
  input   io_channel_status_0_0_occupied,
  output  io_out_allocs_0_0_alloc
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg  mask; // @[SingleVCAllocator.scala 16:21]
  wire  in_arb_reqs_0_0_0 = io_req_0_bits_vc_sel_0_0 & ~io_channel_status_0_0_occupied; // @[SingleVCAllocator.scala 28:61]
  wire  in_arb_vals_0 = io_req_0_valid & in_arb_reqs_0_0_0; // @[SingleVCAllocator.scala 32:39]
  wire  _in_arb_filter_T_1 = in_arb_vals_0 & ~mask; // @[SingleVCAllocator.scala 19:84]
  wire [1:0] _in_arb_filter_T_2 = {in_arb_vals_0,_in_arb_filter_T_1}; // @[Cat.scala 33:92]
  wire [1:0] _in_arb_filter_T_5 = _in_arb_filter_T_2[1] ? 2'h2 : 2'h0; // @[Mux.scala 47:70]
  wire [1:0] in_arb_filter = _in_arb_filter_T_2[0] ? 2'h1 : _in_arb_filter_T_5; // @[Mux.scala 47:70]
  wire  _GEN_0 = in_arb_vals_0 | mask; // @[SingleVCAllocator.scala 21:26 22:10 16:21]
  assign io_req_0_ready = in_arb_filter[0] | in_arb_filter[1]; // @[SingleVCAllocator.scala 20:57]
  assign io_resp_0_vc_sel_0_0 = in_arb_vals_0 & in_arb_reqs_0_0_0; // @[SingleVCAllocator.scala 41:18]
  assign io_out_allocs_0_0_alloc = in_arb_vals_0 & in_arb_reqs_0_0_0; // @[SingleVCAllocator.scala 41:18]
  always @(posedge clock) begin
    if (reset) begin // @[SingleVCAllocator.scala 16:21]
      mask <= 1'h0; // @[SingleVCAllocator.scala 16:21]
    end else begin
      mask <= _GEN_0;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mask = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(1'h1); // @[SingleVCAllocator.scala 53:11]
    end
  end
endmodule
module RouteComputer_1(
  input   clock,
  input   reset,
  input   io_req_0_valid
);
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~io_req_0_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RouteComputer.scala:48 assert(!req.valid)\n"); // @[RouteComputer.scala 48:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(~io_req_0_valid); // @[RouteComputer.scala 48:13]
    end
  end
endmodule
module Router_1(
  input         clock,
  input         reset,
  output [1:0]  auto_debug_out_va_stall_0,
  output [1:0]  auto_debug_out_sa_stall_0,
  output        auto_egress_nodes_out_flit_valid,
  output        auto_egress_nodes_out_flit_bits_head,
  output        auto_egress_nodes_out_flit_bits_tail,
  output [63:0] auto_egress_nodes_out_flit_bits_payload,
  output        auto_egress_nodes_out_flit_bits_ingress_id,
  input         auto_dest_nodes_in_flit_0_valid,
  input         auto_dest_nodes_in_flit_0_bits_head,
  input         auto_dest_nodes_in_flit_0_bits_tail,
  input  [63:0] auto_dest_nodes_in_flit_0_bits_payload,
  input         auto_dest_nodes_in_flit_0_bits_flow_ingress_node,
  input         auto_dest_nodes_in_flit_0_bits_flow_egress_node,
  input  [1:0]  auto_dest_nodes_in_flit_0_bits_virt_channel_id,
  output [2:0]  auto_dest_nodes_in_credit_return,
  output [2:0]  auto_dest_nodes_in_vc_free
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  monitor_clock; // @[Nodes.scala 24:25]
  wire  monitor_reset; // @[Nodes.scala 24:25]
  wire  monitor_io_in_flit_0_valid; // @[Nodes.scala 24:25]
  wire  monitor_io_in_flit_0_bits_head; // @[Nodes.scala 24:25]
  wire  monitor_io_in_flit_0_bits_tail; // @[Nodes.scala 24:25]
  wire  monitor_io_in_flit_0_bits_flow_ingress_node; // @[Nodes.scala 24:25]
  wire  monitor_io_in_flit_0_bits_flow_egress_node; // @[Nodes.scala 24:25]
  wire [1:0] monitor_io_in_flit_0_bits_virt_channel_id; // @[Nodes.scala 24:25]
  wire  input_unit_0_from_0_clock; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_reset; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_router_req_valid; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_0_io_router_req_bits_src_virt_id; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_req_ready; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_req_valid; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_resp_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_out_credit_available_0_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_salloc_req_0_ready; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_salloc_req_0_valid; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_salloc_req_0_bits_tail; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_out_0_valid; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_out_0_bits_flit_head; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_out_0_bits_flit_tail; // @[Router.scala 112:13]
  wire [63:0] input_unit_0_from_0_io_out_0_bits_flit_payload; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_0_io_debug_va_stall; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_0_io_debug_sa_stall; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_in_flit_0_valid; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_in_flit_0_bits_head; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_in_flit_0_bits_tail; // @[Router.scala 112:13]
  wire [63:0] input_unit_0_from_0_io_in_flit_0_bits_payload; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_in_flit_0_bits_flow_egress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_0_io_in_flit_0_bits_virt_channel_id; // @[Router.scala 112:13]
  wire [2:0] input_unit_0_from_0_io_in_credit_return; // @[Router.scala 112:13]
  wire [2:0] input_unit_0_from_0_io_in_vc_free; // @[Router.scala 112:13]
  wire  egress_unit_0_to_0_clock; // @[Router.scala 125:13]
  wire  egress_unit_0_to_0_reset; // @[Router.scala 125:13]
  wire  egress_unit_0_to_0_io_in_0_valid; // @[Router.scala 125:13]
  wire  egress_unit_0_to_0_io_in_0_bits_head; // @[Router.scala 125:13]
  wire  egress_unit_0_to_0_io_in_0_bits_tail; // @[Router.scala 125:13]
  wire [63:0] egress_unit_0_to_0_io_in_0_bits_payload; // @[Router.scala 125:13]
  wire  egress_unit_0_to_0_io_credit_available_0; // @[Router.scala 125:13]
  wire  egress_unit_0_to_0_io_channel_status_0_occupied; // @[Router.scala 125:13]
  wire  egress_unit_0_to_0_io_allocs_0_alloc; // @[Router.scala 125:13]
  wire  egress_unit_0_to_0_io_credit_alloc_0_alloc; // @[Router.scala 125:13]
  wire  egress_unit_0_to_0_io_credit_alloc_0_tail; // @[Router.scala 125:13]
  wire  egress_unit_0_to_0_io_out_valid; // @[Router.scala 125:13]
  wire  egress_unit_0_to_0_io_out_bits_head; // @[Router.scala 125:13]
  wire  egress_unit_0_to_0_io_out_bits_tail; // @[Router.scala 125:13]
  wire [63:0] egress_unit_0_to_0_io_out_bits_payload; // @[Router.scala 125:13]
  wire  egress_unit_0_to_0_io_out_bits_ingress_id; // @[Router.scala 125:13]
  wire  switch_clock; // @[Router.scala 129:24]
  wire  switch_reset; // @[Router.scala 129:24]
  wire  switch_io_in_0_0_valid; // @[Router.scala 129:24]
  wire  switch_io_in_0_0_bits_flit_head; // @[Router.scala 129:24]
  wire  switch_io_in_0_0_bits_flit_tail; // @[Router.scala 129:24]
  wire [63:0] switch_io_in_0_0_bits_flit_payload; // @[Router.scala 129:24]
  wire  switch_io_out_0_0_valid; // @[Router.scala 129:24]
  wire  switch_io_out_0_0_bits_head; // @[Router.scala 129:24]
  wire  switch_io_out_0_0_bits_tail; // @[Router.scala 129:24]
  wire [63:0] switch_io_out_0_0_bits_payload; // @[Router.scala 129:24]
  wire  switch_io_sel_0_0_0_0; // @[Router.scala 129:24]
  wire  switch_allocator_clock; // @[Router.scala 130:34]
  wire  switch_allocator_reset; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_ready; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_valid; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_0_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_tail; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_0_0_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_0_0_tail; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_0_0_0_0; // @[Router.scala 130:34]
  wire  vc_allocator_clock; // @[Router.scala 131:30]
  wire  vc_allocator_reset; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_ready; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_valid; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_0_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_0_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_0_0_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_0_0_alloc; // @[Router.scala 131:30]
  wire  route_computer_clock; // @[Router.scala 134:32]
  wire  route_computer_reset; // @[Router.scala 134:32]
  wire  route_computer_io_req_0_valid; // @[Router.scala 134:32]
  wire [19:0] plusarg_reader_out; // @[PlusArg.scala 80:11]
  reg  switch_io_sel_REG_0_0_0_0; // @[Router.scala 176:14]
  reg [63:0] debug_tsc; // @[Router.scala 193:28]
  wire [63:0] _debug_tsc_T_1 = debug_tsc + 64'h1; // @[Router.scala 194:28]
  reg [63:0] debug_sample; // @[Router.scala 195:31]
  wire [63:0] _debug_sample_T_1 = debug_sample + 64'h1; // @[Router.scala 196:34]
  wire [19:0] _T_1 = plusarg_reader_out - 20'h1; // @[Router.scala 198:40]
  wire [63:0] _GEN_3 = {{44'd0}, _T_1}; // @[Router.scala 198:24]
  wire  _T_2 = debug_sample == _GEN_3; // @[Router.scala 198:24]
  reg [63:0] util_ctr; // @[Router.scala 201:29]
  reg  fired; // @[Router.scala 202:26]
  wire [63:0] _GEN_4 = {{63'd0}, auto_dest_nodes_in_flit_0_valid}; // @[Router.scala 203:28]
  wire [63:0] _util_ctr_T_1 = util_ctr + _GEN_4; // @[Router.scala 203:28]
  wire  _T_8 = plusarg_reader_out != 20'h0 & _T_2 & fired; // @[Router.scala 205:71]
  wire  x1_flit_valid = egress_unit_0_to_0_io_out_valid; // @[Nodes.scala 1212:84 Router.scala 144:65]
  reg [63:0] util_ctr_1; // @[Router.scala 201:29]
  reg  fired_1; // @[Router.scala 202:26]
  wire [63:0] _GEN_6 = {{63'd0}, x1_flit_valid}; // @[Router.scala 203:28]
  wire [63:0] _util_ctr_T_3 = util_ctr_1 + _GEN_6; // @[Router.scala 203:28]
  wire  _T_17 = plusarg_reader_out != 20'h0 & _T_2 & fired_1; // @[Router.scala 205:71]
  wire  fires_count = vc_allocator_io_req_0_ready & vc_allocator_io_req_0_valid; // @[Decoupled.scala 51:35]
  NoCMonitor monitor ( // @[Nodes.scala 24:25]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_flit_0_valid(monitor_io_in_flit_0_valid),
    .io_in_flit_0_bits_head(monitor_io_in_flit_0_bits_head),
    .io_in_flit_0_bits_tail(monitor_io_in_flit_0_bits_tail),
    .io_in_flit_0_bits_flow_ingress_node(monitor_io_in_flit_0_bits_flow_ingress_node),
    .io_in_flit_0_bits_flow_egress_node(monitor_io_in_flit_0_bits_flow_egress_node),
    .io_in_flit_0_bits_virt_channel_id(monitor_io_in_flit_0_bits_virt_channel_id)
  );
  InputUnit input_unit_0_from_0 ( // @[Router.scala 112:13]
    .clock(input_unit_0_from_0_clock),
    .reset(input_unit_0_from_0_reset),
    .io_router_req_valid(input_unit_0_from_0_io_router_req_valid),
    .io_router_req_bits_src_virt_id(input_unit_0_from_0_io_router_req_bits_src_virt_id),
    .io_vcalloc_req_ready(input_unit_0_from_0_io_vcalloc_req_ready),
    .io_vcalloc_req_valid(input_unit_0_from_0_io_vcalloc_req_valid),
    .io_vcalloc_req_bits_vc_sel_0_0(input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_0),
    .io_vcalloc_resp_vc_sel_0_0(input_unit_0_from_0_io_vcalloc_resp_vc_sel_0_0),
    .io_out_credit_available_0_0(input_unit_0_from_0_io_out_credit_available_0_0),
    .io_salloc_req_0_ready(input_unit_0_from_0_io_salloc_req_0_ready),
    .io_salloc_req_0_valid(input_unit_0_from_0_io_salloc_req_0_valid),
    .io_salloc_req_0_bits_vc_sel_0_0(input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_0),
    .io_salloc_req_0_bits_tail(input_unit_0_from_0_io_salloc_req_0_bits_tail),
    .io_out_0_valid(input_unit_0_from_0_io_out_0_valid),
    .io_out_0_bits_flit_head(input_unit_0_from_0_io_out_0_bits_flit_head),
    .io_out_0_bits_flit_tail(input_unit_0_from_0_io_out_0_bits_flit_tail),
    .io_out_0_bits_flit_payload(input_unit_0_from_0_io_out_0_bits_flit_payload),
    .io_debug_va_stall(input_unit_0_from_0_io_debug_va_stall),
    .io_debug_sa_stall(input_unit_0_from_0_io_debug_sa_stall),
    .io_in_flit_0_valid(input_unit_0_from_0_io_in_flit_0_valid),
    .io_in_flit_0_bits_head(input_unit_0_from_0_io_in_flit_0_bits_head),
    .io_in_flit_0_bits_tail(input_unit_0_from_0_io_in_flit_0_bits_tail),
    .io_in_flit_0_bits_payload(input_unit_0_from_0_io_in_flit_0_bits_payload),
    .io_in_flit_0_bits_flow_egress_node(input_unit_0_from_0_io_in_flit_0_bits_flow_egress_node),
    .io_in_flit_0_bits_virt_channel_id(input_unit_0_from_0_io_in_flit_0_bits_virt_channel_id),
    .io_in_credit_return(input_unit_0_from_0_io_in_credit_return),
    .io_in_vc_free(input_unit_0_from_0_io_in_vc_free)
  );
  EgressUnit egress_unit_0_to_0 ( // @[Router.scala 125:13]
    .clock(egress_unit_0_to_0_clock),
    .reset(egress_unit_0_to_0_reset),
    .io_in_0_valid(egress_unit_0_to_0_io_in_0_valid),
    .io_in_0_bits_head(egress_unit_0_to_0_io_in_0_bits_head),
    .io_in_0_bits_tail(egress_unit_0_to_0_io_in_0_bits_tail),
    .io_in_0_bits_payload(egress_unit_0_to_0_io_in_0_bits_payload),
    .io_credit_available_0(egress_unit_0_to_0_io_credit_available_0),
    .io_channel_status_0_occupied(egress_unit_0_to_0_io_channel_status_0_occupied),
    .io_allocs_0_alloc(egress_unit_0_to_0_io_allocs_0_alloc),
    .io_credit_alloc_0_alloc(egress_unit_0_to_0_io_credit_alloc_0_alloc),
    .io_credit_alloc_0_tail(egress_unit_0_to_0_io_credit_alloc_0_tail),
    .io_out_valid(egress_unit_0_to_0_io_out_valid),
    .io_out_bits_head(egress_unit_0_to_0_io_out_bits_head),
    .io_out_bits_tail(egress_unit_0_to_0_io_out_bits_tail),
    .io_out_bits_payload(egress_unit_0_to_0_io_out_bits_payload),
    .io_out_bits_ingress_id(egress_unit_0_to_0_io_out_bits_ingress_id)
  );
  Switch_1 switch ( // @[Router.scala 129:24]
    .clock(switch_clock),
    .reset(switch_reset),
    .io_in_0_0_valid(switch_io_in_0_0_valid),
    .io_in_0_0_bits_flit_head(switch_io_in_0_0_bits_flit_head),
    .io_in_0_0_bits_flit_tail(switch_io_in_0_0_bits_flit_tail),
    .io_in_0_0_bits_flit_payload(switch_io_in_0_0_bits_flit_payload),
    .io_out_0_0_valid(switch_io_out_0_0_valid),
    .io_out_0_0_bits_head(switch_io_out_0_0_bits_head),
    .io_out_0_0_bits_tail(switch_io_out_0_0_bits_tail),
    .io_out_0_0_bits_payload(switch_io_out_0_0_bits_payload),
    .io_sel_0_0_0_0(switch_io_sel_0_0_0_0)
  );
  SwitchAllocator_1 switch_allocator ( // @[Router.scala 130:34]
    .clock(switch_allocator_clock),
    .reset(switch_allocator_reset),
    .io_req_0_0_ready(switch_allocator_io_req_0_0_ready),
    .io_req_0_0_valid(switch_allocator_io_req_0_0_valid),
    .io_req_0_0_bits_vc_sel_0_0(switch_allocator_io_req_0_0_bits_vc_sel_0_0),
    .io_req_0_0_bits_tail(switch_allocator_io_req_0_0_bits_tail),
    .io_credit_alloc_0_0_alloc(switch_allocator_io_credit_alloc_0_0_alloc),
    .io_credit_alloc_0_0_tail(switch_allocator_io_credit_alloc_0_0_tail),
    .io_switch_sel_0_0_0_0(switch_allocator_io_switch_sel_0_0_0_0)
  );
  RotatingSingleVCAllocator_1 vc_allocator ( // @[Router.scala 131:30]
    .clock(vc_allocator_clock),
    .reset(vc_allocator_reset),
    .io_req_0_ready(vc_allocator_io_req_0_ready),
    .io_req_0_valid(vc_allocator_io_req_0_valid),
    .io_req_0_bits_vc_sel_0_0(vc_allocator_io_req_0_bits_vc_sel_0_0),
    .io_resp_0_vc_sel_0_0(vc_allocator_io_resp_0_vc_sel_0_0),
    .io_channel_status_0_0_occupied(vc_allocator_io_channel_status_0_0_occupied),
    .io_out_allocs_0_0_alloc(vc_allocator_io_out_allocs_0_0_alloc)
  );
  RouteComputer_1 route_computer ( // @[Router.scala 134:32]
    .clock(route_computer_clock),
    .reset(route_computer_reset),
    .io_req_0_valid(route_computer_io_req_0_valid)
  );
  plusarg_reader #(.FORMAT("noc_util_sample_rate=%d"), .DEFAULT(0), .WIDTH(20)) plusarg_reader ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_out)
  );
  assign auto_debug_out_va_stall_0 = input_unit_0_from_0_io_debug_va_stall; // @[Nodes.scala 1212:84 Router.scala 190:92]
  assign auto_debug_out_sa_stall_0 = input_unit_0_from_0_io_debug_sa_stall; // @[Nodes.scala 1212:84 Router.scala 191:92]
  assign auto_egress_nodes_out_flit_valid = egress_unit_0_to_0_io_out_valid; // @[Nodes.scala 1212:84 Router.scala 144:65]
  assign auto_egress_nodes_out_flit_bits_head = egress_unit_0_to_0_io_out_bits_head; // @[Nodes.scala 1212:84 Router.scala 144:65]
  assign auto_egress_nodes_out_flit_bits_tail = egress_unit_0_to_0_io_out_bits_tail; // @[Nodes.scala 1212:84 Router.scala 144:65]
  assign auto_egress_nodes_out_flit_bits_payload = egress_unit_0_to_0_io_out_bits_payload; // @[Nodes.scala 1212:84 Router.scala 144:65]
  assign auto_egress_nodes_out_flit_bits_ingress_id = egress_unit_0_to_0_io_out_bits_ingress_id; // @[Nodes.scala 1212:84 Router.scala 144:65]
  assign auto_dest_nodes_in_credit_return = input_unit_0_from_0_io_in_credit_return; // @[Nodes.scala 1215:84 Router.scala 141:68]
  assign auto_dest_nodes_in_vc_free = input_unit_0_from_0_io_in_vc_free; // @[Nodes.scala 1215:84 Router.scala 141:68]
  assign monitor_clock = clock;
  assign monitor_reset = reset;
  assign monitor_io_in_flit_0_valid = auto_dest_nodes_in_flit_0_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_io_in_flit_0_bits_head = auto_dest_nodes_in_flit_0_bits_head; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_io_in_flit_0_bits_tail = auto_dest_nodes_in_flit_0_bits_tail; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_io_in_flit_0_bits_flow_ingress_node = auto_dest_nodes_in_flit_0_bits_flow_ingress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_io_in_flit_0_bits_flow_egress_node = auto_dest_nodes_in_flit_0_bits_flow_egress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_io_in_flit_0_bits_virt_channel_id = auto_dest_nodes_in_flit_0_bits_virt_channel_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_0_clock = clock;
  assign input_unit_0_from_0_reset = reset;
  assign input_unit_0_from_0_io_vcalloc_req_ready = vc_allocator_io_req_0_ready; // @[Router.scala 151:23]
  assign input_unit_0_from_0_io_vcalloc_resp_vc_sel_0_0 = vc_allocator_io_resp_0_vc_sel_0_0; // @[Router.scala 153:39]
  assign input_unit_0_from_0_io_out_credit_available_0_0 = egress_unit_0_to_0_io_credit_available_0; // @[Router.scala 162:42]
  assign input_unit_0_from_0_io_salloc_req_0_ready = switch_allocator_io_req_0_0_ready; // @[Router.scala 165:23]
  assign input_unit_0_from_0_io_in_flit_0_valid = auto_dest_nodes_in_flit_0_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_0_io_in_flit_0_bits_head = auto_dest_nodes_in_flit_0_bits_head; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_0_io_in_flit_0_bits_tail = auto_dest_nodes_in_flit_0_bits_tail; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_0_io_in_flit_0_bits_payload = auto_dest_nodes_in_flit_0_bits_payload; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_0_io_in_flit_0_bits_flow_egress_node = auto_dest_nodes_in_flit_0_bits_flow_egress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_0_io_in_flit_0_bits_virt_channel_id = auto_dest_nodes_in_flit_0_bits_virt_channel_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign egress_unit_0_to_0_clock = clock;
  assign egress_unit_0_to_0_reset = reset;
  assign egress_unit_0_to_0_io_in_0_valid = switch_io_out_0_0_valid; // @[Router.scala 172:29]
  assign egress_unit_0_to_0_io_in_0_bits_head = switch_io_out_0_0_bits_head; // @[Router.scala 172:29]
  assign egress_unit_0_to_0_io_in_0_bits_tail = switch_io_out_0_0_bits_tail; // @[Router.scala 172:29]
  assign egress_unit_0_to_0_io_in_0_bits_payload = switch_io_out_0_0_bits_payload; // @[Router.scala 172:29]
  assign egress_unit_0_to_0_io_allocs_0_alloc = vc_allocator_io_out_allocs_0_0_alloc; // @[Router.scala 157:33]
  assign egress_unit_0_to_0_io_credit_alloc_0_alloc = switch_allocator_io_credit_alloc_0_0_alloc; // @[Router.scala 167:39]
  assign egress_unit_0_to_0_io_credit_alloc_0_tail = switch_allocator_io_credit_alloc_0_0_tail; // @[Router.scala 167:39]
  assign switch_clock = clock;
  assign switch_reset = reset;
  assign switch_io_in_0_0_valid = input_unit_0_from_0_io_out_0_valid; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_head = input_unit_0_from_0_io_out_0_bits_flit_head; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_tail = input_unit_0_from_0_io_out_0_bits_flit_tail; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_payload = input_unit_0_from_0_io_out_0_bits_flit_payload; // @[Router.scala 170:23]
  assign switch_io_sel_0_0_0_0 = switch_io_sel_REG_0_0_0_0; // @[Router.scala 173:19]
  assign switch_allocator_clock = clock;
  assign switch_allocator_reset = reset;
  assign switch_allocator_io_req_0_0_valid = input_unit_0_from_0_io_salloc_req_0_valid; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_0_0 = input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_tail = input_unit_0_from_0_io_salloc_req_0_bits_tail; // @[Router.scala 165:23]
  assign vc_allocator_clock = clock;
  assign vc_allocator_reset = reset;
  assign vc_allocator_io_req_0_valid = input_unit_0_from_0_io_vcalloc_req_valid; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_0_0 = input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_0; // @[Router.scala 151:23]
  assign vc_allocator_io_channel_status_0_0_occupied = egress_unit_0_to_0_io_channel_status_0_occupied; // @[Router.scala 159:23]
  assign route_computer_clock = clock;
  assign route_computer_reset = reset;
  assign route_computer_io_req_0_valid = input_unit_0_from_0_io_router_req_valid; // @[Router.scala 146:23]
  always @(posedge clock) begin
    switch_io_sel_REG_0_0_0_0 <= switch_allocator_io_switch_sel_0_0_0_0; // @[Router.scala 176:14]
    if (reset) begin // @[Router.scala 193:28]
      debug_tsc <= 64'h0; // @[Router.scala 193:28]
    end else begin
      debug_tsc <= _debug_tsc_T_1; // @[Router.scala 194:15]
    end
    if (reset) begin // @[Router.scala 195:31]
      debug_sample <= 64'h0; // @[Router.scala 195:31]
    end else if (debug_sample == _GEN_3) begin // @[Router.scala 198:47]
      debug_sample <= 64'h0; // @[Router.scala 198:62]
    end else begin
      debug_sample <= _debug_sample_T_1; // @[Router.scala 196:18]
    end
    if (reset) begin // @[Router.scala 201:29]
      util_ctr <= 64'h0; // @[Router.scala 201:29]
    end else begin
      util_ctr <= _util_ctr_T_1; // @[Router.scala 203:16]
    end
    if (reset) begin // @[Router.scala 202:26]
      fired <= 1'h0; // @[Router.scala 202:26]
    end else if (plusarg_reader_out != 20'h0 & _T_2 & fired) begin // @[Router.scala 205:81]
      fired <= auto_dest_nodes_in_flit_0_valid; // @[Router.scala 208:15]
    end else begin
      fired <= fired | auto_dest_nodes_in_flit_0_valid; // @[Router.scala 204:13]
    end
    if (reset) begin // @[Router.scala 201:29]
      util_ctr_1 <= 64'h0; // @[Router.scala 201:29]
    end else begin
      util_ctr_1 <= _util_ctr_T_3; // @[Router.scala 203:16]
    end
    if (reset) begin // @[Router.scala 202:26]
      fired_1 <= 1'h0; // @[Router.scala 202:26]
    end else if (plusarg_reader_out != 20'h0 & _T_2 & fired_1) begin // @[Router.scala 205:81]
      fired_1 <= x1_flit_valid; // @[Router.scala 208:15]
    end else begin
      fired_1 <= fired_1 | x1_flit_valid; // @[Router.scala 204:13]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8 & ~reset) begin
          $fwrite(32'h80000002,"nocsample %d 0 1 %d\n",debug_tsc,util_ctr); // @[Router.scala 207:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_17 & ~reset) begin
          $fwrite(32'h80000002,"nocsample %d 1 e0 %d\n",debug_tsc,util_ctr_1); // @[Router.scala 207:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  switch_io_sel_REG_0_0_0_0 = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  debug_tsc = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  debug_sample = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  util_ctr = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  fired = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  util_ctr_1 = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  fired_1 = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ClockSinkDomain_1(
  output [1:0]  auto_routers_debug_out_va_stall_0,
  output [1:0]  auto_routers_debug_out_sa_stall_0,
  output        auto_routers_egress_nodes_out_flit_valid,
  output        auto_routers_egress_nodes_out_flit_bits_head,
  output        auto_routers_egress_nodes_out_flit_bits_tail,
  output [63:0] auto_routers_egress_nodes_out_flit_bits_payload,
  output        auto_routers_egress_nodes_out_flit_bits_ingress_id,
  input         auto_routers_dest_nodes_in_flit_0_valid,
  input         auto_routers_dest_nodes_in_flit_0_bits_head,
  input         auto_routers_dest_nodes_in_flit_0_bits_tail,
  input  [63:0] auto_routers_dest_nodes_in_flit_0_bits_payload,
  input         auto_routers_dest_nodes_in_flit_0_bits_flow_ingress_node,
  input         auto_routers_dest_nodes_in_flit_0_bits_flow_egress_node,
  input  [1:0]  auto_routers_dest_nodes_in_flit_0_bits_virt_channel_id,
  output [2:0]  auto_routers_dest_nodes_in_credit_return,
  output [2:0]  auto_routers_dest_nodes_in_vc_free,
  input         auto_clock_in_clock,
  input         auto_clock_in_reset
);
  wire  routers_clock; // @[NoC.scala 64:22]
  wire  routers_reset; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_debug_out_va_stall_0; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_debug_out_sa_stall_0; // @[NoC.scala 64:22]
  wire  routers_auto_egress_nodes_out_flit_valid; // @[NoC.scala 64:22]
  wire  routers_auto_egress_nodes_out_flit_bits_head; // @[NoC.scala 64:22]
  wire  routers_auto_egress_nodes_out_flit_bits_tail; // @[NoC.scala 64:22]
  wire [63:0] routers_auto_egress_nodes_out_flit_bits_payload; // @[NoC.scala 64:22]
  wire  routers_auto_egress_nodes_out_flit_bits_ingress_id; // @[NoC.scala 64:22]
  wire  routers_auto_dest_nodes_in_flit_0_valid; // @[NoC.scala 64:22]
  wire  routers_auto_dest_nodes_in_flit_0_bits_head; // @[NoC.scala 64:22]
  wire  routers_auto_dest_nodes_in_flit_0_bits_tail; // @[NoC.scala 64:22]
  wire [63:0] routers_auto_dest_nodes_in_flit_0_bits_payload; // @[NoC.scala 64:22]
  wire  routers_auto_dest_nodes_in_flit_0_bits_flow_ingress_node; // @[NoC.scala 64:22]
  wire  routers_auto_dest_nodes_in_flit_0_bits_flow_egress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_dest_nodes_in_flit_0_bits_virt_channel_id; // @[NoC.scala 64:22]
  wire [2:0] routers_auto_dest_nodes_in_credit_return; // @[NoC.scala 64:22]
  wire [2:0] routers_auto_dest_nodes_in_vc_free; // @[NoC.scala 64:22]
  Router_1 routers ( // @[NoC.scala 64:22]
    .clock(routers_clock),
    .reset(routers_reset),
    .auto_debug_out_va_stall_0(routers_auto_debug_out_va_stall_0),
    .auto_debug_out_sa_stall_0(routers_auto_debug_out_sa_stall_0),
    .auto_egress_nodes_out_flit_valid(routers_auto_egress_nodes_out_flit_valid),
    .auto_egress_nodes_out_flit_bits_head(routers_auto_egress_nodes_out_flit_bits_head),
    .auto_egress_nodes_out_flit_bits_tail(routers_auto_egress_nodes_out_flit_bits_tail),
    .auto_egress_nodes_out_flit_bits_payload(routers_auto_egress_nodes_out_flit_bits_payload),
    .auto_egress_nodes_out_flit_bits_ingress_id(routers_auto_egress_nodes_out_flit_bits_ingress_id),
    .auto_dest_nodes_in_flit_0_valid(routers_auto_dest_nodes_in_flit_0_valid),
    .auto_dest_nodes_in_flit_0_bits_head(routers_auto_dest_nodes_in_flit_0_bits_head),
    .auto_dest_nodes_in_flit_0_bits_tail(routers_auto_dest_nodes_in_flit_0_bits_tail),
    .auto_dest_nodes_in_flit_0_bits_payload(routers_auto_dest_nodes_in_flit_0_bits_payload),
    .auto_dest_nodes_in_flit_0_bits_flow_ingress_node(routers_auto_dest_nodes_in_flit_0_bits_flow_ingress_node),
    .auto_dest_nodes_in_flit_0_bits_flow_egress_node(routers_auto_dest_nodes_in_flit_0_bits_flow_egress_node),
    .auto_dest_nodes_in_flit_0_bits_virt_channel_id(routers_auto_dest_nodes_in_flit_0_bits_virt_channel_id),
    .auto_dest_nodes_in_credit_return(routers_auto_dest_nodes_in_credit_return),
    .auto_dest_nodes_in_vc_free(routers_auto_dest_nodes_in_vc_free)
  );
  assign auto_routers_debug_out_va_stall_0 = routers_auto_debug_out_va_stall_0; // @[LazyModule.scala 368:12]
  assign auto_routers_debug_out_sa_stall_0 = routers_auto_debug_out_sa_stall_0; // @[LazyModule.scala 368:12]
  assign auto_routers_egress_nodes_out_flit_valid = routers_auto_egress_nodes_out_flit_valid; // @[LazyModule.scala 368:12]
  assign auto_routers_egress_nodes_out_flit_bits_head = routers_auto_egress_nodes_out_flit_bits_head; // @[LazyModule.scala 368:12]
  assign auto_routers_egress_nodes_out_flit_bits_tail = routers_auto_egress_nodes_out_flit_bits_tail; // @[LazyModule.scala 368:12]
  assign auto_routers_egress_nodes_out_flit_bits_payload = routers_auto_egress_nodes_out_flit_bits_payload; // @[LazyModule.scala 368:12]
  assign auto_routers_egress_nodes_out_flit_bits_ingress_id = routers_auto_egress_nodes_out_flit_bits_ingress_id; // @[LazyModule.scala 368:12]
  assign auto_routers_dest_nodes_in_credit_return = routers_auto_dest_nodes_in_credit_return; // @[LazyModule.scala 366:16]
  assign auto_routers_dest_nodes_in_vc_free = routers_auto_dest_nodes_in_vc_free; // @[LazyModule.scala 366:16]
  assign routers_clock = auto_clock_in_clock; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign routers_reset = auto_clock_in_reset; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_flit_0_valid = auto_routers_dest_nodes_in_flit_0_valid; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_flit_0_bits_head = auto_routers_dest_nodes_in_flit_0_bits_head; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_flit_0_bits_tail = auto_routers_dest_nodes_in_flit_0_bits_tail; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_flit_0_bits_payload = auto_routers_dest_nodes_in_flit_0_bits_payload; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_flit_0_bits_flow_ingress_node =
    auto_routers_dest_nodes_in_flit_0_bits_flow_ingress_node; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_flit_0_bits_flow_egress_node =
    auto_routers_dest_nodes_in_flit_0_bits_flow_egress_node; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_flit_0_bits_virt_channel_id = auto_routers_dest_nodes_in_flit_0_bits_virt_channel_id
    ; // @[LazyModule.scala 366:16]
endmodule
module NoC(
  input         clock,
  input         reset,
  output        io_ingress_0_flit_ready,
  input         io_ingress_0_flit_valid,
  input         io_ingress_0_flit_bits_head,
  input         io_ingress_0_flit_bits_tail,
  input  [63:0] io_ingress_0_flit_bits_payload,
  input         io_ingress_0_flit_bits_egress_id,
  output        io_egress_0_flit_valid,
  output        io_egress_0_flit_bits_head,
  output        io_egress_0_flit_bits_tail,
  output [63:0] io_egress_0_flit_bits_payload,
  output        io_egress_0_flit_bits_ingress_id,
  input         io_router_clocks_0_clock,
  input         io_router_clocks_0_reset,
  input         io_router_clocks_1_clock,
  input         io_router_clocks_1_reset
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  router_sink_domain_auto_routers_ingress_nodes_in_flit_ready; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_routers_ingress_nodes_in_flit_valid; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_routers_ingress_nodes_in_flit_bits_head; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_routers_ingress_nodes_in_flit_bits_tail; // @[NoC.scala 38:40]
  wire [63:0] router_sink_domain_auto_routers_ingress_nodes_in_flit_bits_payload; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_routers_ingress_nodes_in_flit_bits_egress_id; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_routers_source_nodes_out_flit_0_valid; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_routers_source_nodes_out_flit_0_bits_head; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_routers_source_nodes_out_flit_0_bits_tail; // @[NoC.scala 38:40]
  wire [63:0] router_sink_domain_auto_routers_source_nodes_out_flit_0_bits_payload; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_routers_source_nodes_out_flit_0_bits_flow_ingress_node; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_routers_source_nodes_out_flit_0_bits_flow_egress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_auto_routers_source_nodes_out_flit_0_bits_virt_channel_id; // @[NoC.scala 38:40]
  wire [2:0] router_sink_domain_auto_routers_source_nodes_out_credit_return; // @[NoC.scala 38:40]
  wire [2:0] router_sink_domain_auto_routers_source_nodes_out_vc_free; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_clock_in_clock; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_clock_in_reset; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_1_auto_routers_debug_out_va_stall_0; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_1_auto_routers_debug_out_sa_stall_0; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_routers_egress_nodes_out_flit_valid; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_routers_egress_nodes_out_flit_bits_head; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_routers_egress_nodes_out_flit_bits_tail; // @[NoC.scala 38:40]
  wire [63:0] router_sink_domain_1_auto_routers_egress_nodes_out_flit_bits_payload; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_routers_egress_nodes_out_flit_bits_ingress_id; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_routers_dest_nodes_in_flit_0_valid; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_routers_dest_nodes_in_flit_0_bits_head; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_routers_dest_nodes_in_flit_0_bits_tail; // @[NoC.scala 38:40]
  wire [63:0] router_sink_domain_1_auto_routers_dest_nodes_in_flit_0_bits_payload; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_routers_dest_nodes_in_flit_0_bits_flow_ingress_node; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_routers_dest_nodes_in_flit_0_bits_flow_egress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_1_auto_routers_dest_nodes_in_flit_0_bits_virt_channel_id; // @[NoC.scala 38:40]
  wire [2:0] router_sink_domain_1_auto_routers_dest_nodes_in_credit_return; // @[NoC.scala 38:40]
  wire [2:0] router_sink_domain_1_auto_routers_dest_nodes_in_vc_free; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_clock_in_clock; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_clock_in_reset; // @[NoC.scala 38:40]
  reg [63:0] debug_va_stall_ctr; // @[NoC.scala 160:37]
  reg [63:0] debug_sa_stall_ctr; // @[NoC.scala 161:37]
  wire [63:0] debug_any_stall_ctr = debug_va_stall_ctr + debug_sa_stall_ctr; // @[NoC.scala 162:50]
  wire [1:0] bundleIn_0_2_va_stall_0 = router_sink_domain_1_auto_routers_debug_out_va_stall_0; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  wire [2:0] _debug_va_stall_ctr_T = {{1'd0}, bundleIn_0_2_va_stall_0}; // @[NoC.scala 163:104]
  wire [63:0] _GEN_0 = {{62'd0}, _debug_va_stall_ctr_T[1:0]}; // @[NoC.scala 163:46]
  wire [63:0] _debug_va_stall_ctr_T_3 = debug_va_stall_ctr + _GEN_0; // @[NoC.scala 163:46]
  wire [1:0] bundleIn_0_2_sa_stall_0 = router_sink_domain_1_auto_routers_debug_out_sa_stall_0; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  wire [2:0] _debug_sa_stall_ctr_T = {{1'd0}, bundleIn_0_2_sa_stall_0}; // @[NoC.scala 164:104]
  wire [63:0] _GEN_1 = {{62'd0}, _debug_sa_stall_ctr_T[1:0]}; // @[NoC.scala 164:46]
  wire [63:0] _debug_sa_stall_ctr_T_3 = debug_sa_stall_ctr + _GEN_1; // @[NoC.scala 164:46]
  ClockSinkDomain router_sink_domain ( // @[NoC.scala 38:40]
    .auto_routers_ingress_nodes_in_flit_ready(router_sink_domain_auto_routers_ingress_nodes_in_flit_ready),
    .auto_routers_ingress_nodes_in_flit_valid(router_sink_domain_auto_routers_ingress_nodes_in_flit_valid),
    .auto_routers_ingress_nodes_in_flit_bits_head(router_sink_domain_auto_routers_ingress_nodes_in_flit_bits_head),
    .auto_routers_ingress_nodes_in_flit_bits_tail(router_sink_domain_auto_routers_ingress_nodes_in_flit_bits_tail),
    .auto_routers_ingress_nodes_in_flit_bits_payload(router_sink_domain_auto_routers_ingress_nodes_in_flit_bits_payload)
      ,
    .auto_routers_ingress_nodes_in_flit_bits_egress_id(
      router_sink_domain_auto_routers_ingress_nodes_in_flit_bits_egress_id),
    .auto_routers_source_nodes_out_flit_0_valid(router_sink_domain_auto_routers_source_nodes_out_flit_0_valid),
    .auto_routers_source_nodes_out_flit_0_bits_head(router_sink_domain_auto_routers_source_nodes_out_flit_0_bits_head),
    .auto_routers_source_nodes_out_flit_0_bits_tail(router_sink_domain_auto_routers_source_nodes_out_flit_0_bits_tail),
    .auto_routers_source_nodes_out_flit_0_bits_payload(
      router_sink_domain_auto_routers_source_nodes_out_flit_0_bits_payload),
    .auto_routers_source_nodes_out_flit_0_bits_flow_ingress_node(
      router_sink_domain_auto_routers_source_nodes_out_flit_0_bits_flow_ingress_node),
    .auto_routers_source_nodes_out_flit_0_bits_flow_egress_node(
      router_sink_domain_auto_routers_source_nodes_out_flit_0_bits_flow_egress_node),
    .auto_routers_source_nodes_out_flit_0_bits_virt_channel_id(
      router_sink_domain_auto_routers_source_nodes_out_flit_0_bits_virt_channel_id),
    .auto_routers_source_nodes_out_credit_return(router_sink_domain_auto_routers_source_nodes_out_credit_return),
    .auto_routers_source_nodes_out_vc_free(router_sink_domain_auto_routers_source_nodes_out_vc_free),
    .auto_clock_in_clock(router_sink_domain_auto_clock_in_clock),
    .auto_clock_in_reset(router_sink_domain_auto_clock_in_reset)
  );
  ClockSinkDomain_1 router_sink_domain_1 ( // @[NoC.scala 38:40]
    .auto_routers_debug_out_va_stall_0(router_sink_domain_1_auto_routers_debug_out_va_stall_0),
    .auto_routers_debug_out_sa_stall_0(router_sink_domain_1_auto_routers_debug_out_sa_stall_0),
    .auto_routers_egress_nodes_out_flit_valid(router_sink_domain_1_auto_routers_egress_nodes_out_flit_valid),
    .auto_routers_egress_nodes_out_flit_bits_head(router_sink_domain_1_auto_routers_egress_nodes_out_flit_bits_head),
    .auto_routers_egress_nodes_out_flit_bits_tail(router_sink_domain_1_auto_routers_egress_nodes_out_flit_bits_tail),
    .auto_routers_egress_nodes_out_flit_bits_payload(
      router_sink_domain_1_auto_routers_egress_nodes_out_flit_bits_payload),
    .auto_routers_egress_nodes_out_flit_bits_ingress_id(
      router_sink_domain_1_auto_routers_egress_nodes_out_flit_bits_ingress_id),
    .auto_routers_dest_nodes_in_flit_0_valid(router_sink_domain_1_auto_routers_dest_nodes_in_flit_0_valid),
    .auto_routers_dest_nodes_in_flit_0_bits_head(router_sink_domain_1_auto_routers_dest_nodes_in_flit_0_bits_head),
    .auto_routers_dest_nodes_in_flit_0_bits_tail(router_sink_domain_1_auto_routers_dest_nodes_in_flit_0_bits_tail),
    .auto_routers_dest_nodes_in_flit_0_bits_payload(router_sink_domain_1_auto_routers_dest_nodes_in_flit_0_bits_payload)
      ,
    .auto_routers_dest_nodes_in_flit_0_bits_flow_ingress_node(
      router_sink_domain_1_auto_routers_dest_nodes_in_flit_0_bits_flow_ingress_node),
    .auto_routers_dest_nodes_in_flit_0_bits_flow_egress_node(
      router_sink_domain_1_auto_routers_dest_nodes_in_flit_0_bits_flow_egress_node),
    .auto_routers_dest_nodes_in_flit_0_bits_virt_channel_id(
      router_sink_domain_1_auto_routers_dest_nodes_in_flit_0_bits_virt_channel_id),
    .auto_routers_dest_nodes_in_credit_return(router_sink_domain_1_auto_routers_dest_nodes_in_credit_return),
    .auto_routers_dest_nodes_in_vc_free(router_sink_domain_1_auto_routers_dest_nodes_in_vc_free),
    .auto_clock_in_clock(router_sink_domain_1_auto_clock_in_clock),
    .auto_clock_in_reset(router_sink_domain_1_auto_clock_in_reset)
  );
  assign io_ingress_0_flit_ready = router_sink_domain_auto_routers_ingress_nodes_in_flit_ready; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign io_egress_0_flit_valid = router_sink_domain_1_auto_routers_egress_nodes_out_flit_valid; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign io_egress_0_flit_bits_head = router_sink_domain_1_auto_routers_egress_nodes_out_flit_bits_head; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign io_egress_0_flit_bits_tail = router_sink_domain_1_auto_routers_egress_nodes_out_flit_bits_tail; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign io_egress_0_flit_bits_payload = router_sink_domain_1_auto_routers_egress_nodes_out_flit_bits_payload; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign io_egress_0_flit_bits_ingress_id = router_sink_domain_1_auto_routers_egress_nodes_out_flit_bits_ingress_id; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign router_sink_domain_auto_routers_ingress_nodes_in_flit_valid = io_ingress_0_flit_valid; // @[Nodes.scala 1212:84 NoC.scala 145:78]
  assign router_sink_domain_auto_routers_ingress_nodes_in_flit_bits_head = io_ingress_0_flit_bits_head; // @[Nodes.scala 1212:84 NoC.scala 145:78]
  assign router_sink_domain_auto_routers_ingress_nodes_in_flit_bits_tail = io_ingress_0_flit_bits_tail; // @[Nodes.scala 1212:84 NoC.scala 145:78]
  assign router_sink_domain_auto_routers_ingress_nodes_in_flit_bits_payload = io_ingress_0_flit_bits_payload; // @[Nodes.scala 1212:84 NoC.scala 145:78]
  assign router_sink_domain_auto_routers_ingress_nodes_in_flit_bits_egress_id = io_ingress_0_flit_bits_egress_id; // @[Nodes.scala 1212:84 NoC.scala 145:78]
  assign router_sink_domain_auto_routers_source_nodes_out_credit_return =
    router_sink_domain_1_auto_routers_dest_nodes_in_credit_return; // @[LazyModule.scala 355:16]
  assign router_sink_domain_auto_routers_source_nodes_out_vc_free =
    router_sink_domain_1_auto_routers_dest_nodes_in_vc_free; // @[LazyModule.scala 355:16]
  assign router_sink_domain_auto_clock_in_clock = io_router_clocks_0_clock; // @[Nodes.scala 1212:84 NoC.scala 147:88]
  assign router_sink_domain_auto_clock_in_reset = io_router_clocks_0_reset; // @[Nodes.scala 1212:84 NoC.scala 147:88]
  assign router_sink_domain_1_auto_routers_dest_nodes_in_flit_0_valid =
    router_sink_domain_auto_routers_source_nodes_out_flit_0_valid; // @[LazyModule.scala 355:16]
  assign router_sink_domain_1_auto_routers_dest_nodes_in_flit_0_bits_head =
    router_sink_domain_auto_routers_source_nodes_out_flit_0_bits_head; // @[LazyModule.scala 355:16]
  assign router_sink_domain_1_auto_routers_dest_nodes_in_flit_0_bits_tail =
    router_sink_domain_auto_routers_source_nodes_out_flit_0_bits_tail; // @[LazyModule.scala 355:16]
  assign router_sink_domain_1_auto_routers_dest_nodes_in_flit_0_bits_payload =
    router_sink_domain_auto_routers_source_nodes_out_flit_0_bits_payload; // @[LazyModule.scala 355:16]
  assign router_sink_domain_1_auto_routers_dest_nodes_in_flit_0_bits_flow_ingress_node =
    router_sink_domain_auto_routers_source_nodes_out_flit_0_bits_flow_ingress_node; // @[LazyModule.scala 355:16]
  assign router_sink_domain_1_auto_routers_dest_nodes_in_flit_0_bits_flow_egress_node =
    router_sink_domain_auto_routers_source_nodes_out_flit_0_bits_flow_egress_node; // @[LazyModule.scala 355:16]
  assign router_sink_domain_1_auto_routers_dest_nodes_in_flit_0_bits_virt_channel_id =
    router_sink_domain_auto_routers_source_nodes_out_flit_0_bits_virt_channel_id; // @[LazyModule.scala 355:16]
  assign router_sink_domain_1_auto_clock_in_clock = io_router_clocks_1_clock; // @[Nodes.scala 1212:84 NoC.scala 147:88]
  assign router_sink_domain_1_auto_clock_in_reset = io_router_clocks_1_reset; // @[Nodes.scala 1212:84 NoC.scala 147:88]
  always @(posedge clock) begin
    if (reset) begin // @[NoC.scala 160:37]
      debug_va_stall_ctr <= 64'h0; // @[NoC.scala 160:37]
    end else begin
      debug_va_stall_ctr <= _debug_va_stall_ctr_T_3; // @[NoC.scala 163:24]
    end
    if (reset) begin // @[NoC.scala 161:37]
      debug_sa_stall_ctr <= 64'h0; // @[NoC.scala 161:37]
    end else begin
      debug_sa_stall_ctr <= _debug_sa_stall_ctr_T_3; // @[NoC.scala 164:24]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  debug_va_stall_ctr = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  debug_sa_stall_ctr = _RAND_1[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MaxPeriodFibonacciLFSR(
  input   clock,
  input   reset,
  output  io_out_0,
  output  io_out_1,
  output  io_out_2,
  output  io_out_3,
  output  io_out_4,
  output  io_out_5,
  output  io_out_6,
  output  io_out_7,
  output  io_out_8,
  output  io_out_9,
  output  io_out_10,
  output  io_out_11,
  output  io_out_12,
  output  io_out_13,
  output  io_out_14,
  output  io_out_15,
  output  io_out_16,
  output  io_out_17,
  output  io_out_18,
  output  io_out_19
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
`endif // RANDOMIZE_REG_INIT
  reg  state_0; // @[PRNG.scala 55:49]
  reg  state_1; // @[PRNG.scala 55:49]
  reg  state_2; // @[PRNG.scala 55:49]
  reg  state_3; // @[PRNG.scala 55:49]
  reg  state_4; // @[PRNG.scala 55:49]
  reg  state_5; // @[PRNG.scala 55:49]
  reg  state_6; // @[PRNG.scala 55:49]
  reg  state_7; // @[PRNG.scala 55:49]
  reg  state_8; // @[PRNG.scala 55:49]
  reg  state_9; // @[PRNG.scala 55:49]
  reg  state_10; // @[PRNG.scala 55:49]
  reg  state_11; // @[PRNG.scala 55:49]
  reg  state_12; // @[PRNG.scala 55:49]
  reg  state_13; // @[PRNG.scala 55:49]
  reg  state_14; // @[PRNG.scala 55:49]
  reg  state_15; // @[PRNG.scala 55:49]
  reg  state_16; // @[PRNG.scala 55:49]
  reg  state_17; // @[PRNG.scala 55:49]
  reg  state_18; // @[PRNG.scala 55:49]
  reg  state_19; // @[PRNG.scala 55:49]
  wire  _T = state_19 ^ state_16; // @[LFSR.scala 15:41]
  assign io_out_0 = state_0; // @[PRNG.scala 78:10]
  assign io_out_1 = state_1; // @[PRNG.scala 78:10]
  assign io_out_2 = state_2; // @[PRNG.scala 78:10]
  assign io_out_3 = state_3; // @[PRNG.scala 78:10]
  assign io_out_4 = state_4; // @[PRNG.scala 78:10]
  assign io_out_5 = state_5; // @[PRNG.scala 78:10]
  assign io_out_6 = state_6; // @[PRNG.scala 78:10]
  assign io_out_7 = state_7; // @[PRNG.scala 78:10]
  assign io_out_8 = state_8; // @[PRNG.scala 78:10]
  assign io_out_9 = state_9; // @[PRNG.scala 78:10]
  assign io_out_10 = state_10; // @[PRNG.scala 78:10]
  assign io_out_11 = state_11; // @[PRNG.scala 78:10]
  assign io_out_12 = state_12; // @[PRNG.scala 78:10]
  assign io_out_13 = state_13; // @[PRNG.scala 78:10]
  assign io_out_14 = state_14; // @[PRNG.scala 78:10]
  assign io_out_15 = state_15; // @[PRNG.scala 78:10]
  assign io_out_16 = state_16; // @[PRNG.scala 78:10]
  assign io_out_17 = state_17; // @[PRNG.scala 78:10]
  assign io_out_18 = state_18; // @[PRNG.scala 78:10]
  assign io_out_19 = state_19; // @[PRNG.scala 78:10]
  always @(posedge clock) begin
    state_0 <= reset | _T; // @[PRNG.scala 55:{49,49}]
    if (reset) begin // @[PRNG.scala 55:49]
      state_1 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_1 <= state_0;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_2 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_2 <= state_1;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_3 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_3 <= state_2;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_4 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_4 <= state_3;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_5 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_5 <= state_4;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_6 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_6 <= state_5;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_7 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_7 <= state_6;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_8 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_8 <= state_7;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_9 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_9 <= state_8;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_10 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_10 <= state_9;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_11 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_11 <= state_10;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_12 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_12 <= state_11;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_13 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_13 <= state_12;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_14 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_14 <= state_13;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_15 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_15 <= state_14;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_16 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_16 <= state_15;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_17 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_17 <= state_16;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_18 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_18 <= state_17;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_19 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_19 <= state_18;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  state_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  state_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  state_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  state_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  state_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  state_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  state_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  state_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  state_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  state_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  state_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  state_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  state_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  state_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  state_15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  state_16 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  state_17 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  state_18 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  state_19 = _RAND_19[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module InputGen(
  input         clock,
  input         reset,
  input         io_out_ready,
  output        io_out_valid,
  output        io_out_bits_head,
  output        io_out_bits_tail,
  output [63:0] io_out_bits_payload,
  input         io_rob_ready,
  input  [6:0]  io_rob_idx,
  input  [31:0] io_tsc,
  output        io_fire,
  output [3:0]  io_n_flits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  packet_remaining_prng_clock; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_reset; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_0; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_1; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_2; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_3; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_4; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_5; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_6; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_7; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_8; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_9; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_10; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_11; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_12; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_13; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_14; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_15; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_16; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_17; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_18; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_19; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_clock; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_reset; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_0; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_1; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_2; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_3; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_4; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_5; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_6; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_7; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_8; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_9; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_10; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_11; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_12; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_13; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_14; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_15; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_16; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_17; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_18; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_19; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_clock; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_reset; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_0; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_1; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_2; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_3; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_4; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_5; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_6; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_7; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_8; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_9; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_10; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_11; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_12; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_13; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_14; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_15; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_16; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_17; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_18; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_19; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_clock; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_reset; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_0; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_1; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_2; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_3; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_4; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_5; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_6; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_7; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_8; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_9; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_10; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_11; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_12; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_13; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_14; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_15; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_16; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_17; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_18; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_19; // @[PRNG.scala 91:22]
  reg [3:0] flits_left; // @[TestHarness.scala 71:27]
  reg [3:0] flits_fired; // @[TestHarness.scala 72:28]
  reg [31:0] payload_tsc; // @[TestHarness.scala 74:20]
  reg [15:0] payload_rob_idx; // @[TestHarness.scala 74:20]
  wire  can_fire = flits_left == 4'h0 & io_rob_ready; // @[TestHarness.scala 76:39]
  wire [9:0] packet_remaining_lo = {packet_remaining_prng_io_out_9,packet_remaining_prng_io_out_8,
    packet_remaining_prng_io_out_7,packet_remaining_prng_io_out_6,packet_remaining_prng_io_out_5,
    packet_remaining_prng_io_out_4,packet_remaining_prng_io_out_3,packet_remaining_prng_io_out_2,
    packet_remaining_prng_io_out_1,packet_remaining_prng_io_out_0}; // @[PRNG.scala 95:17]
  wire [9:0] packet_remaining_hi = {packet_remaining_prng_io_out_19,packet_remaining_prng_io_out_18,
    packet_remaining_prng_io_out_17,packet_remaining_prng_io_out_16,packet_remaining_prng_io_out_15,
    packet_remaining_prng_io_out_14,packet_remaining_prng_io_out_13,packet_remaining_prng_io_out_12,
    packet_remaining_prng_io_out_11,packet_remaining_prng_io_out_10}; // @[PRNG.scala 95:17]
  wire [19:0] _packet_remaining_T = {packet_remaining_hi,packet_remaining_lo}; // @[PRNG.scala 95:17]
  wire [19:0] _GEN_1 = _packet_remaining_T % 20'h8; // @[TestHarness.scala 78:89]
  wire [3:0] packet_remaining = _GEN_1[3:0]; // @[TestHarness.scala 78:89]
  wire [31:0] out_payload_tsc = flits_left != 4'h0 ? payload_tsc : io_tsc; // @[TestHarness.scala 100:29 105:17 87:19]
  wire [15:0] out_payload_rob_idx = flits_left != 4'h0 ? payload_rob_idx : {{9'd0}, io_rob_idx}; // @[TestHarness.scala 100:29 105:17 88:23]
  wire [47:0] io_out_bits_payload_hi = {out_payload_tsc,out_payload_rob_idx}; // @[TestHarness.scala 86:38]
  wire [3:0] _GEN_14 = flits_left != 4'h0 ? flits_fired : 4'h0; // @[TestHarness.scala 100:29 106:29 89:27]
  wire [15:0] out_payload_flits_fired = {{12'd0}, _GEN_14}; // @[TestHarness.scala 85:25]
  wire  _io_fire_T = io_out_ready & io_out_valid; // @[Decoupled.scala 51:35]
  wire [3:0] _GEN_0 = io_fire & ~io_out_bits_tail ? packet_remaining : flits_left; // @[TestHarness.scala 94:39 95:16 71:27]
  wire [3:0] _GEN_5 = io_fire & ~io_out_bits_tail ? 4'h1 : flits_fired; // @[TestHarness.scala 94:39 98:17 72:28]
  wire [3:0] _flits_fired_T_1 = flits_fired + 4'h1; // @[TestHarness.scala 109:34]
  wire [3:0] _flits_left_T_1 = flits_left - 4'h1; // @[TestHarness.scala 110:32]
  MaxPeriodFibonacciLFSR packet_remaining_prng ( // @[PRNG.scala 91:22]
    .clock(packet_remaining_prng_clock),
    .reset(packet_remaining_prng_reset),
    .io_out_0(packet_remaining_prng_io_out_0),
    .io_out_1(packet_remaining_prng_io_out_1),
    .io_out_2(packet_remaining_prng_io_out_2),
    .io_out_3(packet_remaining_prng_io_out_3),
    .io_out_4(packet_remaining_prng_io_out_4),
    .io_out_5(packet_remaining_prng_io_out_5),
    .io_out_6(packet_remaining_prng_io_out_6),
    .io_out_7(packet_remaining_prng_io_out_7),
    .io_out_8(packet_remaining_prng_io_out_8),
    .io_out_9(packet_remaining_prng_io_out_9),
    .io_out_10(packet_remaining_prng_io_out_10),
    .io_out_11(packet_remaining_prng_io_out_11),
    .io_out_12(packet_remaining_prng_io_out_12),
    .io_out_13(packet_remaining_prng_io_out_13),
    .io_out_14(packet_remaining_prng_io_out_14),
    .io_out_15(packet_remaining_prng_io_out_15),
    .io_out_16(packet_remaining_prng_io_out_16),
    .io_out_17(packet_remaining_prng_io_out_17),
    .io_out_18(packet_remaining_prng_io_out_18),
    .io_out_19(packet_remaining_prng_io_out_19)
  );
  MaxPeriodFibonacciLFSR random_flit_delay_prng ( // @[PRNG.scala 91:22]
    .clock(random_flit_delay_prng_clock),
    .reset(random_flit_delay_prng_reset),
    .io_out_0(random_flit_delay_prng_io_out_0),
    .io_out_1(random_flit_delay_prng_io_out_1),
    .io_out_2(random_flit_delay_prng_io_out_2),
    .io_out_3(random_flit_delay_prng_io_out_3),
    .io_out_4(random_flit_delay_prng_io_out_4),
    .io_out_5(random_flit_delay_prng_io_out_5),
    .io_out_6(random_flit_delay_prng_io_out_6),
    .io_out_7(random_flit_delay_prng_io_out_7),
    .io_out_8(random_flit_delay_prng_io_out_8),
    .io_out_9(random_flit_delay_prng_io_out_9),
    .io_out_10(random_flit_delay_prng_io_out_10),
    .io_out_11(random_flit_delay_prng_io_out_11),
    .io_out_12(random_flit_delay_prng_io_out_12),
    .io_out_13(random_flit_delay_prng_io_out_13),
    .io_out_14(random_flit_delay_prng_io_out_14),
    .io_out_15(random_flit_delay_prng_io_out_15),
    .io_out_16(random_flit_delay_prng_io_out_16),
    .io_out_17(random_flit_delay_prng_io_out_17),
    .io_out_18(random_flit_delay_prng_io_out_18),
    .io_out_19(random_flit_delay_prng_io_out_19)
  );
  MaxPeriodFibonacciLFSR random_packet_delay_prng ( // @[PRNG.scala 91:22]
    .clock(random_packet_delay_prng_clock),
    .reset(random_packet_delay_prng_reset),
    .io_out_0(random_packet_delay_prng_io_out_0),
    .io_out_1(random_packet_delay_prng_io_out_1),
    .io_out_2(random_packet_delay_prng_io_out_2),
    .io_out_3(random_packet_delay_prng_io_out_3),
    .io_out_4(random_packet_delay_prng_io_out_4),
    .io_out_5(random_packet_delay_prng_io_out_5),
    .io_out_6(random_packet_delay_prng_io_out_6),
    .io_out_7(random_packet_delay_prng_io_out_7),
    .io_out_8(random_packet_delay_prng_io_out_8),
    .io_out_9(random_packet_delay_prng_io_out_9),
    .io_out_10(random_packet_delay_prng_io_out_10),
    .io_out_11(random_packet_delay_prng_io_out_11),
    .io_out_12(random_packet_delay_prng_io_out_12),
    .io_out_13(random_packet_delay_prng_io_out_13),
    .io_out_14(random_packet_delay_prng_io_out_14),
    .io_out_15(random_packet_delay_prng_io_out_15),
    .io_out_16(random_packet_delay_prng_io_out_16),
    .io_out_17(random_packet_delay_prng_io_out_17),
    .io_out_18(random_packet_delay_prng_io_out_18),
    .io_out_19(random_packet_delay_prng_io_out_19)
  );
  MaxPeriodFibonacciLFSR io_out_bits_egress_id_prng ( // @[PRNG.scala 91:22]
    .clock(io_out_bits_egress_id_prng_clock),
    .reset(io_out_bits_egress_id_prng_reset),
    .io_out_0(io_out_bits_egress_id_prng_io_out_0),
    .io_out_1(io_out_bits_egress_id_prng_io_out_1),
    .io_out_2(io_out_bits_egress_id_prng_io_out_2),
    .io_out_3(io_out_bits_egress_id_prng_io_out_3),
    .io_out_4(io_out_bits_egress_id_prng_io_out_4),
    .io_out_5(io_out_bits_egress_id_prng_io_out_5),
    .io_out_6(io_out_bits_egress_id_prng_io_out_6),
    .io_out_7(io_out_bits_egress_id_prng_io_out_7),
    .io_out_8(io_out_bits_egress_id_prng_io_out_8),
    .io_out_9(io_out_bits_egress_id_prng_io_out_9),
    .io_out_10(io_out_bits_egress_id_prng_io_out_10),
    .io_out_11(io_out_bits_egress_id_prng_io_out_11),
    .io_out_12(io_out_bits_egress_id_prng_io_out_12),
    .io_out_13(io_out_bits_egress_id_prng_io_out_13),
    .io_out_14(io_out_bits_egress_id_prng_io_out_14),
    .io_out_15(io_out_bits_egress_id_prng_io_out_15),
    .io_out_16(io_out_bits_egress_id_prng_io_out_16),
    .io_out_17(io_out_bits_egress_id_prng_io_out_17),
    .io_out_18(io_out_bits_egress_id_prng_io_out_18),
    .io_out_19(io_out_bits_egress_id_prng_io_out_19)
  );
  assign io_out_valid = flits_left != 4'h0 | can_fire; // @[TestHarness.scala 100:29 101:18 81:16]
  assign io_out_bits_head = flits_left != 4'h0 ? 1'h0 : 1'h1; // @[TestHarness.scala 100:29 102:22 82:20]
  assign io_out_bits_tail = flits_left != 4'h0 ? flits_left == 4'h1 : packet_remaining == 4'h0; // @[TestHarness.scala 100:29 103:22 83:20]
  assign io_out_bits_payload = {io_out_bits_payload_hi,out_payload_flits_fired}; // @[TestHarness.scala 86:38]
  assign io_fire = can_fire & _io_fire_T; // @[TestHarness.scala 92:23]
  assign io_n_flits = packet_remaining + 4'h1; // @[TestHarness.scala 91:34]
  assign packet_remaining_prng_clock = clock;
  assign packet_remaining_prng_reset = reset;
  assign random_flit_delay_prng_clock = clock;
  assign random_flit_delay_prng_reset = reset;
  assign random_packet_delay_prng_clock = clock;
  assign random_packet_delay_prng_reset = reset;
  assign io_out_bits_egress_id_prng_clock = clock;
  assign io_out_bits_egress_id_prng_reset = reset;
  always @(posedge clock) begin
    if (reset) begin // @[TestHarness.scala 71:27]
      flits_left <= 4'h0; // @[TestHarness.scala 71:27]
    end else if (flits_left != 4'h0) begin // @[TestHarness.scala 100:29]
      if (_io_fire_T) begin // @[TestHarness.scala 108:26]
        flits_left <= _flits_left_T_1; // @[TestHarness.scala 110:18]
      end else begin
        flits_left <= _GEN_0;
      end
    end else begin
      flits_left <= _GEN_0;
    end
    if (reset) begin // @[TestHarness.scala 72:28]
      flits_fired <= 4'h0; // @[TestHarness.scala 72:28]
    end else if (flits_left != 4'h0) begin // @[TestHarness.scala 100:29]
      if (_io_fire_T) begin // @[TestHarness.scala 108:26]
        flits_fired <= _flits_fired_T_1; // @[TestHarness.scala 109:19]
      end else begin
        flits_fired <= _GEN_5;
      end
    end else begin
      flits_fired <= _GEN_5;
    end
    if (io_fire & ~io_out_bits_tail) begin // @[TestHarness.scala 94:39]
      if (!(flits_left != 4'h0)) begin // @[TestHarness.scala 100:29]
        payload_tsc <= io_tsc; // @[TestHarness.scala 87:19]
      end
    end
    if (io_fire & ~io_out_bits_tail) begin // @[TestHarness.scala 94:39]
      if (!(flits_left != 4'h0)) begin // @[TestHarness.scala 100:29]
        payload_rob_idx <= {{9'd0}, io_rob_idx}; // @[TestHarness.scala 88:23]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  flits_left = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  flits_fired = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  payload_tsc = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  payload_rob_idx = _RAND_3[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_8(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_head,
  input         io_enq_bits_tail,
  input  [63:0] io_enq_bits_payload,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_head,
  output        io_deq_bits_tail,
  output [63:0] io_deq_bits_payload,
  output        io_deq_bits_egress_id
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg  ram_head [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_head_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_head_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_head_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_tail [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_tail_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_tail_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_tail_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_en; // @[Decoupled.scala 273:95]
  reg [63:0] ram_payload [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_payload_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_payload_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [63:0] ram_payload_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [63:0] ram_payload_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_payload_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_payload_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_payload_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_egress_id [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_egress_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_egress_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_egress_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_egress_id_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_egress_id_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_egress_id_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_egress_id_MPORT_en; // @[Decoupled.scala 273:95]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 278:28]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  wire  _GEN_12 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 318:26 280:27 318:35]
  wire  do_enq = empty ? _GEN_12 : _do_enq_T; // @[Decoupled.scala 315:17 280:27]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 315:17 317:14 281:27]
  assign ram_head_io_deq_bits_MPORT_en = 1'h1;
  assign ram_head_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_head_io_deq_bits_MPORT_data = ram_head[ram_head_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_head_MPORT_data = io_enq_bits_head;
  assign ram_head_MPORT_addr = 1'h0;
  assign ram_head_MPORT_mask = 1'h1;
  assign ram_head_MPORT_en = empty ? _GEN_12 : _do_enq_T;
  assign ram_tail_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tail_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tail_io_deq_bits_MPORT_data = ram_tail[ram_tail_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_tail_MPORT_data = io_enq_bits_tail;
  assign ram_tail_MPORT_addr = 1'h0;
  assign ram_tail_MPORT_mask = 1'h1;
  assign ram_tail_MPORT_en = empty ? _GEN_12 : _do_enq_T;
  assign ram_payload_io_deq_bits_MPORT_en = 1'h1;
  assign ram_payload_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_payload_io_deq_bits_MPORT_data = ram_payload[ram_payload_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_payload_MPORT_data = io_enq_bits_payload;
  assign ram_payload_MPORT_addr = 1'h0;
  assign ram_payload_MPORT_mask = 1'h1;
  assign ram_payload_MPORT_en = empty ? _GEN_12 : _do_enq_T;
  assign ram_egress_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_egress_id_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_egress_id_io_deq_bits_MPORT_data = ram_egress_id[ram_egress_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_egress_id_MPORT_data = 1'h0;
  assign ram_egress_id_MPORT_addr = 1'h0;
  assign ram_egress_id_MPORT_mask = 1'h1;
  assign ram_egress_id_MPORT_en = empty ? _GEN_12 : _do_enq_T;
  assign io_enq_ready = io_deq_ready | empty; // @[Decoupled.scala 303:16 323:{24,39}]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 302:16 314:{24,39}]
  assign io_deq_bits_head = empty ? io_enq_bits_head : ram_head_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_tail = empty ? io_enq_bits_tail : ram_tail_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_payload = empty ? io_enq_bits_payload : ram_payload_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_egress_id = empty ? 1'h0 : ram_egress_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  always @(posedge clock) begin
    if (ram_head_MPORT_en & ram_head_MPORT_mask) begin
      ram_head[ram_head_MPORT_addr] <= ram_head_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_tail_MPORT_en & ram_tail_MPORT_mask) begin
      ram_tail[ram_tail_MPORT_addr] <= ram_tail_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_payload_MPORT_en & ram_payload_MPORT_mask) begin
      ram_payload[ram_payload_MPORT_addr] <= ram_payload_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_egress_id_MPORT_en & ram_egress_id_MPORT_mask) begin
      ram_egress_id[ram_egress_id_MPORT_addr] <= ram_egress_id_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      if (empty) begin // @[Decoupled.scala 315:17]
        if (io_deq_ready) begin // @[Decoupled.scala 318:26]
          maybe_full <= 1'h0; // @[Decoupled.scala 318:35]
        end else begin
          maybe_full <= _do_enq_T; // @[Decoupled.scala 280:27]
        end
      end else begin
        maybe_full <= _do_enq_T; // @[Decoupled.scala 280:27]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_head[initvar] = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tail[initvar] = _RAND_1[0:0];
  _RAND_2 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload[initvar] = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_egress_id[initvar] = _RAND_3[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  maybe_full = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module NoCTester(
  input         clock,
  input         reset,
  input         io_to_noc_0_flit_ready,
  output        io_to_noc_0_flit_valid,
  output        io_to_noc_0_flit_bits_head,
  output        io_to_noc_0_flit_bits_tail,
  output [63:0] io_to_noc_0_flit_bits_payload,
  output        io_to_noc_0_flit_bits_egress_id,
  output        io_from_noc_0_flit_ready,
  input         io_from_noc_0_flit_valid,
  input         io_from_noc_0_flit_bits_head,
  input         io_from_noc_0_flit_bits_tail,
  input  [63:0] io_from_noc_0_flit_bits_payload,
  input         io_from_noc_0_flit_bits_ingress_id,
  output        io_success
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [127:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [63:0] _RAND_645;
  reg [63:0] _RAND_646;
  reg [63:0] _RAND_647;
  reg [63:0] _RAND_648;
  reg [63:0] _RAND_649;
  reg [63:0] _RAND_650;
  reg [63:0] _RAND_651;
  reg [63:0] _RAND_652;
  reg [63:0] _RAND_653;
  reg [63:0] _RAND_654;
  reg [63:0] _RAND_655;
  reg [63:0] _RAND_656;
  reg [63:0] _RAND_657;
  reg [63:0] _RAND_658;
  reg [63:0] _RAND_659;
  reg [63:0] _RAND_660;
  reg [63:0] _RAND_661;
  reg [63:0] _RAND_662;
  reg [63:0] _RAND_663;
  reg [63:0] _RAND_664;
  reg [63:0] _RAND_665;
  reg [63:0] _RAND_666;
  reg [63:0] _RAND_667;
  reg [63:0] _RAND_668;
  reg [63:0] _RAND_669;
  reg [63:0] _RAND_670;
  reg [63:0] _RAND_671;
  reg [63:0] _RAND_672;
  reg [63:0] _RAND_673;
  reg [63:0] _RAND_674;
  reg [63:0] _RAND_675;
  reg [63:0] _RAND_676;
  reg [63:0] _RAND_677;
  reg [63:0] _RAND_678;
  reg [63:0] _RAND_679;
  reg [63:0] _RAND_680;
  reg [63:0] _RAND_681;
  reg [63:0] _RAND_682;
  reg [63:0] _RAND_683;
  reg [63:0] _RAND_684;
  reg [63:0] _RAND_685;
  reg [63:0] _RAND_686;
  reg [63:0] _RAND_687;
  reg [63:0] _RAND_688;
  reg [63:0] _RAND_689;
  reg [63:0] _RAND_690;
  reg [63:0] _RAND_691;
  reg [63:0] _RAND_692;
  reg [63:0] _RAND_693;
  reg [63:0] _RAND_694;
  reg [63:0] _RAND_695;
  reg [63:0] _RAND_696;
  reg [63:0] _RAND_697;
  reg [63:0] _RAND_698;
  reg [63:0] _RAND_699;
  reg [63:0] _RAND_700;
  reg [63:0] _RAND_701;
  reg [63:0] _RAND_702;
  reg [63:0] _RAND_703;
  reg [63:0] _RAND_704;
  reg [63:0] _RAND_705;
  reg [63:0] _RAND_706;
  reg [63:0] _RAND_707;
  reg [63:0] _RAND_708;
  reg [63:0] _RAND_709;
  reg [63:0] _RAND_710;
  reg [63:0] _RAND_711;
  reg [63:0] _RAND_712;
  reg [63:0] _RAND_713;
  reg [63:0] _RAND_714;
  reg [63:0] _RAND_715;
  reg [63:0] _RAND_716;
  reg [63:0] _RAND_717;
  reg [63:0] _RAND_718;
  reg [63:0] _RAND_719;
  reg [63:0] _RAND_720;
  reg [63:0] _RAND_721;
  reg [63:0] _RAND_722;
  reg [63:0] _RAND_723;
  reg [63:0] _RAND_724;
  reg [63:0] _RAND_725;
  reg [63:0] _RAND_726;
  reg [63:0] _RAND_727;
  reg [63:0] _RAND_728;
  reg [63:0] _RAND_729;
  reg [63:0] _RAND_730;
  reg [63:0] _RAND_731;
  reg [63:0] _RAND_732;
  reg [63:0] _RAND_733;
  reg [63:0] _RAND_734;
  reg [63:0] _RAND_735;
  reg [63:0] _RAND_736;
  reg [63:0] _RAND_737;
  reg [63:0] _RAND_738;
  reg [63:0] _RAND_739;
  reg [63:0] _RAND_740;
  reg [63:0] _RAND_741;
  reg [63:0] _RAND_742;
  reg [63:0] _RAND_743;
  reg [63:0] _RAND_744;
  reg [63:0] _RAND_745;
  reg [63:0] _RAND_746;
  reg [63:0] _RAND_747;
  reg [63:0] _RAND_748;
  reg [63:0] _RAND_749;
  reg [63:0] _RAND_750;
  reg [63:0] _RAND_751;
  reg [63:0] _RAND_752;
  reg [63:0] _RAND_753;
  reg [63:0] _RAND_754;
  reg [63:0] _RAND_755;
  reg [63:0] _RAND_756;
  reg [63:0] _RAND_757;
  reg [63:0] _RAND_758;
  reg [63:0] _RAND_759;
  reg [63:0] _RAND_760;
  reg [63:0] _RAND_761;
  reg [63:0] _RAND_762;
  reg [63:0] _RAND_763;
  reg [63:0] _RAND_764;
  reg [63:0] _RAND_765;
  reg [63:0] _RAND_766;
  reg [63:0] _RAND_767;
  reg [63:0] _RAND_768;
  reg [63:0] _RAND_769;
  reg [63:0] _RAND_770;
  reg [63:0] _RAND_771;
  reg [63:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
`endif // RANDOMIZE_REG_INIT
  wire  igen_clock; // @[TestHarness.scala 171:22]
  wire  igen_reset; // @[TestHarness.scala 171:22]
  wire  igen_io_out_ready; // @[TestHarness.scala 171:22]
  wire  igen_io_out_valid; // @[TestHarness.scala 171:22]
  wire  igen_io_out_bits_head; // @[TestHarness.scala 171:22]
  wire  igen_io_out_bits_tail; // @[TestHarness.scala 171:22]
  wire [63:0] igen_io_out_bits_payload; // @[TestHarness.scala 171:22]
  wire  igen_io_rob_ready; // @[TestHarness.scala 171:22]
  wire [6:0] igen_io_rob_idx; // @[TestHarness.scala 171:22]
  wire [31:0] igen_io_tsc; // @[TestHarness.scala 171:22]
  wire  igen_io_fire; // @[TestHarness.scala 171:22]
  wire [3:0] igen_io_n_flits; // @[TestHarness.scala 171:22]
  wire  io_to_noc_0_flit_q_clock; // @[Decoupled.scala 375:21]
  wire  io_to_noc_0_flit_q_reset; // @[Decoupled.scala 375:21]
  wire  io_to_noc_0_flit_q_io_enq_ready; // @[Decoupled.scala 375:21]
  wire  io_to_noc_0_flit_q_io_enq_valid; // @[Decoupled.scala 375:21]
  wire  io_to_noc_0_flit_q_io_enq_bits_head; // @[Decoupled.scala 375:21]
  wire  io_to_noc_0_flit_q_io_enq_bits_tail; // @[Decoupled.scala 375:21]
  wire [63:0] io_to_noc_0_flit_q_io_enq_bits_payload; // @[Decoupled.scala 375:21]
  wire  io_to_noc_0_flit_q_io_deq_ready; // @[Decoupled.scala 375:21]
  wire  io_to_noc_0_flit_q_io_deq_valid; // @[Decoupled.scala 375:21]
  wire  io_to_noc_0_flit_q_io_deq_bits_head; // @[Decoupled.scala 375:21]
  wire  io_to_noc_0_flit_q_io_deq_bits_tail; // @[Decoupled.scala 375:21]
  wire [63:0] io_to_noc_0_flit_q_io_deq_bits_payload; // @[Decoupled.scala 375:21]
  wire  io_to_noc_0_flit_q_io_deq_bits_egress_id; // @[Decoupled.scala 375:21]
  wire  plusarg_reader_out; // @[PlusArg.scala 80:11]
  wire  io_from_noc_0_flit_ready_prng_clock; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_reset; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_0; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_1; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_2; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_3; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_4; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_5; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_6; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_7; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_8; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_9; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_10; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_11; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_12; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_13; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_14; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_15; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_16; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_17; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_18; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_19; // @[PRNG.scala 91:22]
  reg [31:0] txs; // @[TestHarness.scala 136:20]
  reg [31:0] flits; // @[TestHarness.scala 137:22]
  reg [31:0] tsc; // @[TestHarness.scala 141:20]
  wire [31:0] _tsc_T_1 = tsc + 32'h1; // @[TestHarness.scala 142:14]
  reg [10:0] idle_counter; // @[TestHarness.scala 144:29]
  wire [10:0] _idle_counter_T_1 = idle_counter + 11'h1; // @[TestHarness.scala 146:46]
  reg [127:0] rob_valids; // @[TestHarness.scala 156:27]
  wire [127:0] _T_5 = ~rob_valids; // @[TestHarness.scala 161:59]
  wire [6:0] _sels_0_T_128 = _T_5[126] ? 7'h7e : 7'h7f; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_129 = _T_5[125] ? 7'h7d : _sels_0_T_128; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_130 = _T_5[124] ? 7'h7c : _sels_0_T_129; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_131 = _T_5[123] ? 7'h7b : _sels_0_T_130; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_132 = _T_5[122] ? 7'h7a : _sels_0_T_131; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_133 = _T_5[121] ? 7'h79 : _sels_0_T_132; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_134 = _T_5[120] ? 7'h78 : _sels_0_T_133; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_135 = _T_5[119] ? 7'h77 : _sels_0_T_134; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_136 = _T_5[118] ? 7'h76 : _sels_0_T_135; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_137 = _T_5[117] ? 7'h75 : _sels_0_T_136; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_138 = _T_5[116] ? 7'h74 : _sels_0_T_137; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_139 = _T_5[115] ? 7'h73 : _sels_0_T_138; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_140 = _T_5[114] ? 7'h72 : _sels_0_T_139; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_141 = _T_5[113] ? 7'h71 : _sels_0_T_140; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_142 = _T_5[112] ? 7'h70 : _sels_0_T_141; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_143 = _T_5[111] ? 7'h6f : _sels_0_T_142; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_144 = _T_5[110] ? 7'h6e : _sels_0_T_143; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_145 = _T_5[109] ? 7'h6d : _sels_0_T_144; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_146 = _T_5[108] ? 7'h6c : _sels_0_T_145; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_147 = _T_5[107] ? 7'h6b : _sels_0_T_146; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_148 = _T_5[106] ? 7'h6a : _sels_0_T_147; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_149 = _T_5[105] ? 7'h69 : _sels_0_T_148; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_150 = _T_5[104] ? 7'h68 : _sels_0_T_149; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_151 = _T_5[103] ? 7'h67 : _sels_0_T_150; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_152 = _T_5[102] ? 7'h66 : _sels_0_T_151; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_153 = _T_5[101] ? 7'h65 : _sels_0_T_152; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_154 = _T_5[100] ? 7'h64 : _sels_0_T_153; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_155 = _T_5[99] ? 7'h63 : _sels_0_T_154; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_156 = _T_5[98] ? 7'h62 : _sels_0_T_155; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_157 = _T_5[97] ? 7'h61 : _sels_0_T_156; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_158 = _T_5[96] ? 7'h60 : _sels_0_T_157; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_159 = _T_5[95] ? 7'h5f : _sels_0_T_158; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_160 = _T_5[94] ? 7'h5e : _sels_0_T_159; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_161 = _T_5[93] ? 7'h5d : _sels_0_T_160; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_162 = _T_5[92] ? 7'h5c : _sels_0_T_161; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_163 = _T_5[91] ? 7'h5b : _sels_0_T_162; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_164 = _T_5[90] ? 7'h5a : _sels_0_T_163; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_165 = _T_5[89] ? 7'h59 : _sels_0_T_164; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_166 = _T_5[88] ? 7'h58 : _sels_0_T_165; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_167 = _T_5[87] ? 7'h57 : _sels_0_T_166; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_168 = _T_5[86] ? 7'h56 : _sels_0_T_167; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_169 = _T_5[85] ? 7'h55 : _sels_0_T_168; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_170 = _T_5[84] ? 7'h54 : _sels_0_T_169; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_171 = _T_5[83] ? 7'h53 : _sels_0_T_170; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_172 = _T_5[82] ? 7'h52 : _sels_0_T_171; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_173 = _T_5[81] ? 7'h51 : _sels_0_T_172; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_174 = _T_5[80] ? 7'h50 : _sels_0_T_173; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_175 = _T_5[79] ? 7'h4f : _sels_0_T_174; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_176 = _T_5[78] ? 7'h4e : _sels_0_T_175; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_177 = _T_5[77] ? 7'h4d : _sels_0_T_176; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_178 = _T_5[76] ? 7'h4c : _sels_0_T_177; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_179 = _T_5[75] ? 7'h4b : _sels_0_T_178; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_180 = _T_5[74] ? 7'h4a : _sels_0_T_179; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_181 = _T_5[73] ? 7'h49 : _sels_0_T_180; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_182 = _T_5[72] ? 7'h48 : _sels_0_T_181; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_183 = _T_5[71] ? 7'h47 : _sels_0_T_182; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_184 = _T_5[70] ? 7'h46 : _sels_0_T_183; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_185 = _T_5[69] ? 7'h45 : _sels_0_T_184; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_186 = _T_5[68] ? 7'h44 : _sels_0_T_185; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_187 = _T_5[67] ? 7'h43 : _sels_0_T_186; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_188 = _T_5[66] ? 7'h42 : _sels_0_T_187; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_189 = _T_5[65] ? 7'h41 : _sels_0_T_188; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_190 = _T_5[64] ? 7'h40 : _sels_0_T_189; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_191 = _T_5[63] ? 7'h3f : _sels_0_T_190; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_192 = _T_5[62] ? 7'h3e : _sels_0_T_191; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_193 = _T_5[61] ? 7'h3d : _sels_0_T_192; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_194 = _T_5[60] ? 7'h3c : _sels_0_T_193; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_195 = _T_5[59] ? 7'h3b : _sels_0_T_194; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_196 = _T_5[58] ? 7'h3a : _sels_0_T_195; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_197 = _T_5[57] ? 7'h39 : _sels_0_T_196; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_198 = _T_5[56] ? 7'h38 : _sels_0_T_197; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_199 = _T_5[55] ? 7'h37 : _sels_0_T_198; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_200 = _T_5[54] ? 7'h36 : _sels_0_T_199; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_201 = _T_5[53] ? 7'h35 : _sels_0_T_200; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_202 = _T_5[52] ? 7'h34 : _sels_0_T_201; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_203 = _T_5[51] ? 7'h33 : _sels_0_T_202; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_204 = _T_5[50] ? 7'h32 : _sels_0_T_203; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_205 = _T_5[49] ? 7'h31 : _sels_0_T_204; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_206 = _T_5[48] ? 7'h30 : _sels_0_T_205; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_207 = _T_5[47] ? 7'h2f : _sels_0_T_206; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_208 = _T_5[46] ? 7'h2e : _sels_0_T_207; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_209 = _T_5[45] ? 7'h2d : _sels_0_T_208; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_210 = _T_5[44] ? 7'h2c : _sels_0_T_209; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_211 = _T_5[43] ? 7'h2b : _sels_0_T_210; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_212 = _T_5[42] ? 7'h2a : _sels_0_T_211; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_213 = _T_5[41] ? 7'h29 : _sels_0_T_212; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_214 = _T_5[40] ? 7'h28 : _sels_0_T_213; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_215 = _T_5[39] ? 7'h27 : _sels_0_T_214; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_216 = _T_5[38] ? 7'h26 : _sels_0_T_215; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_217 = _T_5[37] ? 7'h25 : _sels_0_T_216; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_218 = _T_5[36] ? 7'h24 : _sels_0_T_217; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_219 = _T_5[35] ? 7'h23 : _sels_0_T_218; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_220 = _T_5[34] ? 7'h22 : _sels_0_T_219; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_221 = _T_5[33] ? 7'h21 : _sels_0_T_220; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_222 = _T_5[32] ? 7'h20 : _sels_0_T_221; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_223 = _T_5[31] ? 7'h1f : _sels_0_T_222; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_224 = _T_5[30] ? 7'h1e : _sels_0_T_223; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_225 = _T_5[29] ? 7'h1d : _sels_0_T_224; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_226 = _T_5[28] ? 7'h1c : _sels_0_T_225; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_227 = _T_5[27] ? 7'h1b : _sels_0_T_226; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_228 = _T_5[26] ? 7'h1a : _sels_0_T_227; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_229 = _T_5[25] ? 7'h19 : _sels_0_T_228; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_230 = _T_5[24] ? 7'h18 : _sels_0_T_229; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_231 = _T_5[23] ? 7'h17 : _sels_0_T_230; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_232 = _T_5[22] ? 7'h16 : _sels_0_T_231; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_233 = _T_5[21] ? 7'h15 : _sels_0_T_232; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_234 = _T_5[20] ? 7'h14 : _sels_0_T_233; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_235 = _T_5[19] ? 7'h13 : _sels_0_T_234; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_236 = _T_5[18] ? 7'h12 : _sels_0_T_235; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_237 = _T_5[17] ? 7'h11 : _sels_0_T_236; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_238 = _T_5[16] ? 7'h10 : _sels_0_T_237; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_239 = _T_5[15] ? 7'hf : _sels_0_T_238; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_240 = _T_5[14] ? 7'he : _sels_0_T_239; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_241 = _T_5[13] ? 7'hd : _sels_0_T_240; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_242 = _T_5[12] ? 7'hc : _sels_0_T_241; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_243 = _T_5[11] ? 7'hb : _sels_0_T_242; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_244 = _T_5[10] ? 7'ha : _sels_0_T_243; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_245 = _T_5[9] ? 7'h9 : _sels_0_T_244; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_246 = _T_5[8] ? 7'h8 : _sels_0_T_245; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_247 = _T_5[7] ? 7'h7 : _sels_0_T_246; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_248 = _T_5[6] ? 7'h6 : _sels_0_T_247; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_249 = _T_5[5] ? 7'h5 : _sels_0_T_248; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_250 = _T_5[4] ? 7'h4 : _sels_0_T_249; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_251 = _T_5[3] ? 7'h3 : _sels_0_T_250; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_252 = _T_5[2] ? 7'h2 : _sels_0_T_251; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_253 = _T_5[1] ? 7'h1 : _sels_0_T_252; // @[Mux.scala 47:70]
  wire [6:0] rob_alloc_ids_0 = _T_5[0] ? 7'h0 : _sels_0_T_253; // @[Mux.scala 47:70]
  wire [127:0] _GEN_389 = {{127'd0}, igen_io_fire}; // @[TestHarness.scala 187:45]
  wire [127:0] rob_allocs = _GEN_389 << rob_alloc_ids_0; // @[TestHarness.scala 187:45]
  wire  _T_67 = io_from_noc_0_flit_ready & io_from_noc_0_flit_valid; // @[Decoupled.scala 51:35]
  wire  _T_68 = _T_67 & io_from_noc_0_flit_bits_tail; // @[TestHarness.scala 218:45]
  wire [15:0] out_payload_rob_idx = io_from_noc_0_flit_bits_payload[31:16]; // @[TestHarness.scala 194:51]
  wire [65535:0] _GEN_390 = {{65535'd0}, _T_68}; // @[TestHarness.scala 218:66]
  wire [65535:0] rob_frees = _GEN_390 << out_payload_rob_idx; // @[TestHarness.scala 218:66]
  wire  idle = rob_allocs == 128'h0 & rob_frees == 65536'h0; // @[TestHarness.scala 223:30]
  wire  _T_3 = ~reset; // @[TestHarness.scala 148:9]
  reg [31:0] rob_payload_0_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_0_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_0_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_1_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_1_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_1_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_2_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_2_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_2_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_3_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_3_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_3_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_4_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_4_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_4_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_5_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_5_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_5_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_6_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_6_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_6_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_7_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_7_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_7_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_8_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_8_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_8_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_9_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_9_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_9_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_10_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_10_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_10_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_11_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_11_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_11_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_12_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_12_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_12_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_13_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_13_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_13_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_14_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_14_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_14_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_15_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_15_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_15_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_16_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_16_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_16_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_17_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_17_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_17_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_18_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_18_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_18_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_19_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_19_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_19_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_20_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_20_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_20_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_21_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_21_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_21_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_22_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_22_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_22_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_23_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_23_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_23_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_24_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_24_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_24_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_25_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_25_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_25_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_26_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_26_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_26_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_27_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_27_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_27_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_28_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_28_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_28_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_29_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_29_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_29_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_30_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_30_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_30_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_31_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_31_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_31_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_32_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_32_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_32_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_33_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_33_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_33_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_34_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_34_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_34_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_35_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_35_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_35_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_36_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_36_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_36_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_37_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_37_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_37_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_38_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_38_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_38_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_39_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_39_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_39_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_40_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_40_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_40_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_41_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_41_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_41_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_42_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_42_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_42_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_43_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_43_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_43_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_44_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_44_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_44_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_45_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_45_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_45_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_46_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_46_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_46_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_47_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_47_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_47_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_48_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_48_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_48_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_49_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_49_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_49_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_50_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_50_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_50_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_51_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_51_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_51_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_52_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_52_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_52_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_53_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_53_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_53_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_54_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_54_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_54_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_55_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_55_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_55_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_56_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_56_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_56_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_57_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_57_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_57_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_58_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_58_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_58_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_59_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_59_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_59_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_60_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_60_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_60_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_61_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_61_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_61_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_62_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_62_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_62_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_63_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_63_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_63_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_64_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_64_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_64_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_65_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_65_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_65_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_66_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_66_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_66_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_67_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_67_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_67_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_68_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_68_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_68_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_69_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_69_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_69_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_70_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_70_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_70_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_71_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_71_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_71_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_72_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_72_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_72_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_73_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_73_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_73_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_74_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_74_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_74_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_75_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_75_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_75_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_76_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_76_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_76_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_77_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_77_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_77_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_78_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_78_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_78_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_79_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_79_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_79_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_80_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_80_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_80_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_81_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_81_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_81_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_82_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_82_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_82_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_83_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_83_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_83_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_84_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_84_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_84_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_85_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_85_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_85_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_86_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_86_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_86_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_87_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_87_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_87_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_88_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_88_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_88_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_89_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_89_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_89_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_90_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_90_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_90_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_91_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_91_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_91_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_92_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_92_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_92_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_93_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_93_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_93_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_94_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_94_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_94_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_95_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_95_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_95_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_96_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_96_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_96_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_97_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_97_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_97_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_98_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_98_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_98_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_99_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_99_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_99_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_100_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_100_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_100_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_101_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_101_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_101_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_102_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_102_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_102_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_103_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_103_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_103_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_104_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_104_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_104_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_105_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_105_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_105_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_106_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_106_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_106_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_107_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_107_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_107_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_108_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_108_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_108_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_109_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_109_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_109_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_110_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_110_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_110_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_111_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_111_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_111_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_112_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_112_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_112_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_113_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_113_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_113_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_114_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_114_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_114_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_115_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_115_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_115_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_116_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_116_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_116_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_117_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_117_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_117_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_118_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_118_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_118_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_119_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_119_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_119_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_120_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_120_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_120_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_121_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_121_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_121_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_122_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_122_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_122_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_123_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_123_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_123_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_124_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_124_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_124_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_125_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_125_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_125_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_126_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_126_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_126_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_127_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_127_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_127_flits_fired; // @[TestHarness.scala 150:24]
  reg [3:0] rob_n_flits_0; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_1; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_2; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_3; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_4; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_5; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_6; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_7; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_8; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_9; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_10; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_11; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_12; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_13; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_14; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_15; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_16; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_17; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_18; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_19; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_20; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_21; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_22; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_23; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_24; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_25; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_26; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_27; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_28; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_29; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_30; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_31; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_32; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_33; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_34; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_35; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_36; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_37; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_38; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_39; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_40; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_41; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_42; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_43; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_44; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_45; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_46; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_47; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_48; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_49; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_50; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_51; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_52; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_53; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_54; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_55; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_56; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_57; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_58; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_59; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_60; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_61; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_62; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_63; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_64; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_65; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_66; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_67; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_68; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_69; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_70; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_71; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_72; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_73; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_74; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_75; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_76; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_77; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_78; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_79; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_80; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_81; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_82; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_83; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_84; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_85; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_86; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_87; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_88; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_89; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_90; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_91; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_92; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_93; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_94; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_95; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_96; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_97; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_98; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_99; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_100; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_101; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_102; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_103; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_104; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_105; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_106; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_107; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_108; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_109; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_110; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_111; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_112; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_113; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_114; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_115; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_116; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_117; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_118; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_119; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_120; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_121; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_122; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_123; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_124; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_125; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_126; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_127; // @[TestHarness.scala 153:24]
  reg [3:0] rob_flits_returned_0; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_1; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_2; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_3; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_4; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_5; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_6; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_7; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_8; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_9; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_10; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_11; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_12; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_13; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_14; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_15; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_16; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_17; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_18; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_19; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_20; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_21; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_22; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_23; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_24; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_25; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_26; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_27; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_28; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_29; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_30; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_31; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_32; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_33; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_34; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_35; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_36; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_37; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_38; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_39; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_40; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_41; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_42; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_43; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_44; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_45; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_46; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_47; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_48; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_49; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_50; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_51; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_52; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_53; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_54; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_55; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_56; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_57; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_58; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_59; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_60; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_61; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_62; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_63; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_64; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_65; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_66; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_67; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_68; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_69; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_70; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_71; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_72; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_73; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_74; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_75; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_76; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_77; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_78; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_79; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_80; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_81; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_82; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_83; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_84; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_85; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_86; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_87; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_88; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_89; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_90; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_91; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_92; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_93; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_94; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_95; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_96; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_97; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_98; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_99; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_100; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_101; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_102; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_103; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_104; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_105; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_106; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_107; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_108; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_109; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_110; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_111; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_112; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_113; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_114; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_115; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_116; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_117; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_118; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_119; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_120; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_121; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_122; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_123; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_124; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_125; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_126; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_127; // @[TestHarness.scala 154:31]
  reg [63:0] rob_tscs_0; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_1; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_2; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_3; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_4; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_5; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_6; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_7; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_8; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_9; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_10; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_11; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_12; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_13; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_14; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_15; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_16; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_17; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_18; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_19; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_20; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_21; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_22; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_23; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_24; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_25; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_26; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_27; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_28; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_29; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_30; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_31; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_32; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_33; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_34; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_35; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_36; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_37; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_38; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_39; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_40; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_41; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_42; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_43; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_44; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_45; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_46; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_47; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_48; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_49; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_50; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_51; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_52; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_53; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_54; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_55; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_56; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_57; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_58; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_59; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_60; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_61; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_62; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_63; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_64; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_65; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_66; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_67; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_68; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_69; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_70; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_71; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_72; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_73; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_74; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_75; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_76; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_77; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_78; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_79; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_80; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_81; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_82; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_83; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_84; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_85; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_86; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_87; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_88; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_89; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_90; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_91; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_92; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_93; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_94; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_95; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_96; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_97; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_98; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_99; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_100; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_101; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_102; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_103; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_104; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_105; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_106; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_107; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_108; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_109; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_110; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_111; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_112; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_113; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_114; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_115; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_116; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_117; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_118; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_119; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_120; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_121; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_122; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_123; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_124; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_125; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_126; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_127; // @[TestHarness.scala 155:21]
  wire  rob_alloc_fires_0 = _T_5 != 128'h0; // @[TestHarness.scala 30:24]
  wire [127:0] _rob_alloc_avail_T = rob_valids >> rob_alloc_ids_0; // @[TestHarness.scala 162:61]
  wire  rob_alloc_avail_0 = ~_rob_alloc_avail_T[0]; // @[TestHarness.scala 162:50]
  wire  success = txs >= 32'hc350 & rob_valids == 128'h0; // @[TestHarness.scala 163:35]
  reg  io_success_REG; // @[TestHarness.scala 164:24]
  wire  _igen_io_rob_ready_T_1 = tsc >= 32'ha; // @[TestHarness.scala 175:11]
  wire  _igen_io_rob_ready_T_2 = rob_alloc_avail_0 & rob_alloc_fires_0 & _igen_io_rob_ready_T_1; // @[TestHarness.scala 174:72]
  wire [63:0] _rob_payload_WIRE_1 = igen_io_out_bits_payload; // @[TestHarness.scala 179:{72,72}]
  wire [15:0] _GEN_257 = 7'h0 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_0_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_258 = 7'h1 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_1_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_259 = 7'h2 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_2_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_260 = 7'h3 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_3_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_261 = 7'h4 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_4_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_262 = 7'h5 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_5_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_263 = 7'h6 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_6_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_264 = 7'h7 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_7_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_265 = 7'h8 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_8_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_266 = 7'h9 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_9_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_267 = 7'ha == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_10_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_268 = 7'hb == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_11_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_269 = 7'hc == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_12_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_270 = 7'hd == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_13_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_271 = 7'he == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_14_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_272 = 7'hf == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_15_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_273 = 7'h10 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_16_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_274 = 7'h11 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_17_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_275 = 7'h12 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_18_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_276 = 7'h13 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_19_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_277 = 7'h14 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_20_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_278 = 7'h15 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_21_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_279 = 7'h16 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_22_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_280 = 7'h17 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_23_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_281 = 7'h18 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_24_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_282 = 7'h19 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_25_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_283 = 7'h1a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_26_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_284 = 7'h1b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_27_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_285 = 7'h1c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_28_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_286 = 7'h1d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_29_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_287 = 7'h1e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_30_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_288 = 7'h1f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_31_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_289 = 7'h20 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_32_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_290 = 7'h21 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_33_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_291 = 7'h22 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_34_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_292 = 7'h23 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_35_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_293 = 7'h24 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_36_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_294 = 7'h25 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_37_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_295 = 7'h26 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_38_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_296 = 7'h27 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_39_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_297 = 7'h28 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_40_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_298 = 7'h29 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_41_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_299 = 7'h2a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_42_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_300 = 7'h2b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_43_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_301 = 7'h2c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_44_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_302 = 7'h2d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_45_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_303 = 7'h2e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_46_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_304 = 7'h2f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_47_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_305 = 7'h30 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_48_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_306 = 7'h31 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_49_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_307 = 7'h32 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_50_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_308 = 7'h33 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_51_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_309 = 7'h34 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_52_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_310 = 7'h35 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_53_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_311 = 7'h36 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_54_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_312 = 7'h37 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_55_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_313 = 7'h38 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_56_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_314 = 7'h39 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_57_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_315 = 7'h3a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_58_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_316 = 7'h3b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_59_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_317 = 7'h3c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_60_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_318 = 7'h3d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_61_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_319 = 7'h3e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_62_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_320 = 7'h3f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_63_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_321 = 7'h40 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_64_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_322 = 7'h41 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_65_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_323 = 7'h42 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_66_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_324 = 7'h43 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_67_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_325 = 7'h44 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_68_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_326 = 7'h45 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_69_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_327 = 7'h46 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_70_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_328 = 7'h47 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_71_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_329 = 7'h48 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_72_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_330 = 7'h49 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_73_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_331 = 7'h4a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_74_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_332 = 7'h4b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_75_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_333 = 7'h4c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_76_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_334 = 7'h4d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_77_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_335 = 7'h4e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_78_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_336 = 7'h4f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_79_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_337 = 7'h50 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_80_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_338 = 7'h51 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_81_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_339 = 7'h52 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_82_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_340 = 7'h53 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_83_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_341 = 7'h54 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_84_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_342 = 7'h55 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_85_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_343 = 7'h56 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_86_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_344 = 7'h57 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_87_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_345 = 7'h58 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_88_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_346 = 7'h59 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_89_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_347 = 7'h5a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_90_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_348 = 7'h5b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_91_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_349 = 7'h5c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_92_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_350 = 7'h5d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_93_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_351 = 7'h5e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_94_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_352 = 7'h5f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_95_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_353 = 7'h60 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_96_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_354 = 7'h61 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_97_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_355 = 7'h62 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_98_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_356 = 7'h63 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_99_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_357 = 7'h64 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_100_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_358 = 7'h65 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_101_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_359 = 7'h66 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_102_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_360 = 7'h67 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_103_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_361 = 7'h68 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_104_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_362 = 7'h69 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_105_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_363 = 7'h6a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_106_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_364 = 7'h6b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_107_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_365 = 7'h6c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_108_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_366 = 7'h6d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_109_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_367 = 7'h6e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_110_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_368 = 7'h6f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_111_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_369 = 7'h70 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_112_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_370 = 7'h71 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_113_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_371 = 7'h72 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_114_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_372 = 7'h73 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_115_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_373 = 7'h74 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_116_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_374 = 7'h75 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_117_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_375 = 7'h76 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_118_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_376 = 7'h77 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_119_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_377 = 7'h78 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_120_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_378 = 7'h79 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_121_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_379 = 7'h7a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_122_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_380 = 7'h7b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_123_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_381 = 7'h7c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_124_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_382 = 7'h7d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_125_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_383 = 7'h7e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_126_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_384 = 7'h7f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_127_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [3:0] _rob_n_flits_T_18 = igen_io_n_flits; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_769 = 7'h0 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_0; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_770 = 7'h1 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_1; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_771 = 7'h2 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_2; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_772 = 7'h3 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_3; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_773 = 7'h4 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_4; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_774 = 7'h5 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_5; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_775 = 7'h6 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_6; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_776 = 7'h7 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_7; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_777 = 7'h8 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_8; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_778 = 7'h9 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_9; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_779 = 7'ha == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_10; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_780 = 7'hb == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_11; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_781 = 7'hc == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_12; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_782 = 7'hd == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_13; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_783 = 7'he == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_14; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_784 = 7'hf == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_15; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_785 = 7'h10 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_16; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_786 = 7'h11 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_17; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_787 = 7'h12 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_18; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_788 = 7'h13 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_19; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_789 = 7'h14 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_20; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_790 = 7'h15 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_21; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_791 = 7'h16 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_22; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_792 = 7'h17 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_23; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_793 = 7'h18 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_24; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_794 = 7'h19 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_25; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_795 = 7'h1a == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_26; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_796 = 7'h1b == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_27; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_797 = 7'h1c == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_28; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_798 = 7'h1d == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_29; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_799 = 7'h1e == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_30; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_800 = 7'h1f == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_31; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_801 = 7'h20 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_32; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_802 = 7'h21 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_33; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_803 = 7'h22 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_34; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_804 = 7'h23 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_35; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_805 = 7'h24 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_36; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_806 = 7'h25 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_37; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_807 = 7'h26 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_38; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_808 = 7'h27 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_39; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_809 = 7'h28 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_40; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_810 = 7'h29 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_41; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_811 = 7'h2a == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_42; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_812 = 7'h2b == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_43; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_813 = 7'h2c == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_44; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_814 = 7'h2d == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_45; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_815 = 7'h2e == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_46; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_816 = 7'h2f == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_47; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_817 = 7'h30 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_48; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_818 = 7'h31 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_49; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_819 = 7'h32 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_50; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_820 = 7'h33 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_51; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_821 = 7'h34 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_52; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_822 = 7'h35 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_53; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_823 = 7'h36 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_54; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_824 = 7'h37 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_55; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_825 = 7'h38 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_56; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_826 = 7'h39 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_57; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_827 = 7'h3a == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_58; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_828 = 7'h3b == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_59; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_829 = 7'h3c == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_60; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_830 = 7'h3d == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_61; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_831 = 7'h3e == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_62; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_832 = 7'h3f == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_63; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_833 = 7'h40 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_64; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_834 = 7'h41 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_65; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_835 = 7'h42 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_66; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_836 = 7'h43 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_67; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_837 = 7'h44 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_68; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_838 = 7'h45 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_69; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_839 = 7'h46 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_70; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_840 = 7'h47 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_71; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_841 = 7'h48 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_72; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_842 = 7'h49 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_73; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_843 = 7'h4a == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_74; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_844 = 7'h4b == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_75; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_845 = 7'h4c == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_76; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_846 = 7'h4d == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_77; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_847 = 7'h4e == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_78; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_848 = 7'h4f == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_79; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_849 = 7'h50 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_80; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_850 = 7'h51 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_81; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_851 = 7'h52 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_82; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_852 = 7'h53 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_83; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_853 = 7'h54 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_84; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_854 = 7'h55 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_85; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_855 = 7'h56 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_86; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_856 = 7'h57 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_87; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_857 = 7'h58 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_88; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_858 = 7'h59 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_89; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_859 = 7'h5a == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_90; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_860 = 7'h5b == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_91; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_861 = 7'h5c == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_92; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_862 = 7'h5d == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_93; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_863 = 7'h5e == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_94; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_864 = 7'h5f == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_95; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_865 = 7'h60 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_96; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_866 = 7'h61 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_97; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_867 = 7'h62 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_98; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_868 = 7'h63 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_99; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_869 = 7'h64 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_100; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_870 = 7'h65 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_101; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_871 = 7'h66 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_102; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_872 = 7'h67 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_103; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_873 = 7'h68 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_104; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_874 = 7'h69 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_105; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_875 = 7'h6a == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_106; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_876 = 7'h6b == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_107; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_877 = 7'h6c == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_108; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_878 = 7'h6d == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_109; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_879 = 7'h6e == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_110; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_880 = 7'h6f == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_111; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_881 = 7'h70 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_112; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_882 = 7'h71 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_113; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_883 = 7'h72 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_114; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_884 = 7'h73 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_115; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_885 = 7'h74 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_116; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_886 = 7'h75 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_117; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_887 = 7'h76 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_118; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_888 = 7'h77 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_119; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_889 = 7'h78 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_120; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_890 = 7'h79 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_121; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_891 = 7'h7a == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_122; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_892 = 7'h7b == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_123; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_893 = 7'h7c == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_124; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_894 = 7'h7d == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_125; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_895 = 7'h7e == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_126; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_896 = 7'h7f == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_127; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [63:0] _rob_tscs_T_22 = {{32'd0}, tsc}; // @[TestHarness.scala 184:{36,36}]
  wire [15:0] _GEN_1281 = igen_io_fire ? _GEN_257 : rob_payload_0_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1282 = igen_io_fire ? _GEN_258 : rob_payload_1_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1283 = igen_io_fire ? _GEN_259 : rob_payload_2_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1284 = igen_io_fire ? _GEN_260 : rob_payload_3_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1285 = igen_io_fire ? _GEN_261 : rob_payload_4_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1286 = igen_io_fire ? _GEN_262 : rob_payload_5_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1287 = igen_io_fire ? _GEN_263 : rob_payload_6_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1288 = igen_io_fire ? _GEN_264 : rob_payload_7_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1289 = igen_io_fire ? _GEN_265 : rob_payload_8_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1290 = igen_io_fire ? _GEN_266 : rob_payload_9_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1291 = igen_io_fire ? _GEN_267 : rob_payload_10_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1292 = igen_io_fire ? _GEN_268 : rob_payload_11_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1293 = igen_io_fire ? _GEN_269 : rob_payload_12_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1294 = igen_io_fire ? _GEN_270 : rob_payload_13_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1295 = igen_io_fire ? _GEN_271 : rob_payload_14_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1296 = igen_io_fire ? _GEN_272 : rob_payload_15_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1297 = igen_io_fire ? _GEN_273 : rob_payload_16_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1298 = igen_io_fire ? _GEN_274 : rob_payload_17_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1299 = igen_io_fire ? _GEN_275 : rob_payload_18_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1300 = igen_io_fire ? _GEN_276 : rob_payload_19_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1301 = igen_io_fire ? _GEN_277 : rob_payload_20_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1302 = igen_io_fire ? _GEN_278 : rob_payload_21_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1303 = igen_io_fire ? _GEN_279 : rob_payload_22_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1304 = igen_io_fire ? _GEN_280 : rob_payload_23_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1305 = igen_io_fire ? _GEN_281 : rob_payload_24_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1306 = igen_io_fire ? _GEN_282 : rob_payload_25_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1307 = igen_io_fire ? _GEN_283 : rob_payload_26_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1308 = igen_io_fire ? _GEN_284 : rob_payload_27_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1309 = igen_io_fire ? _GEN_285 : rob_payload_28_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1310 = igen_io_fire ? _GEN_286 : rob_payload_29_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1311 = igen_io_fire ? _GEN_287 : rob_payload_30_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1312 = igen_io_fire ? _GEN_288 : rob_payload_31_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1313 = igen_io_fire ? _GEN_289 : rob_payload_32_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1314 = igen_io_fire ? _GEN_290 : rob_payload_33_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1315 = igen_io_fire ? _GEN_291 : rob_payload_34_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1316 = igen_io_fire ? _GEN_292 : rob_payload_35_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1317 = igen_io_fire ? _GEN_293 : rob_payload_36_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1318 = igen_io_fire ? _GEN_294 : rob_payload_37_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1319 = igen_io_fire ? _GEN_295 : rob_payload_38_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1320 = igen_io_fire ? _GEN_296 : rob_payload_39_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1321 = igen_io_fire ? _GEN_297 : rob_payload_40_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1322 = igen_io_fire ? _GEN_298 : rob_payload_41_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1323 = igen_io_fire ? _GEN_299 : rob_payload_42_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1324 = igen_io_fire ? _GEN_300 : rob_payload_43_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1325 = igen_io_fire ? _GEN_301 : rob_payload_44_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1326 = igen_io_fire ? _GEN_302 : rob_payload_45_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1327 = igen_io_fire ? _GEN_303 : rob_payload_46_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1328 = igen_io_fire ? _GEN_304 : rob_payload_47_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1329 = igen_io_fire ? _GEN_305 : rob_payload_48_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1330 = igen_io_fire ? _GEN_306 : rob_payload_49_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1331 = igen_io_fire ? _GEN_307 : rob_payload_50_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1332 = igen_io_fire ? _GEN_308 : rob_payload_51_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1333 = igen_io_fire ? _GEN_309 : rob_payload_52_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1334 = igen_io_fire ? _GEN_310 : rob_payload_53_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1335 = igen_io_fire ? _GEN_311 : rob_payload_54_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1336 = igen_io_fire ? _GEN_312 : rob_payload_55_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1337 = igen_io_fire ? _GEN_313 : rob_payload_56_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1338 = igen_io_fire ? _GEN_314 : rob_payload_57_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1339 = igen_io_fire ? _GEN_315 : rob_payload_58_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1340 = igen_io_fire ? _GEN_316 : rob_payload_59_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1341 = igen_io_fire ? _GEN_317 : rob_payload_60_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1342 = igen_io_fire ? _GEN_318 : rob_payload_61_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1343 = igen_io_fire ? _GEN_319 : rob_payload_62_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1344 = igen_io_fire ? _GEN_320 : rob_payload_63_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1345 = igen_io_fire ? _GEN_321 : rob_payload_64_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1346 = igen_io_fire ? _GEN_322 : rob_payload_65_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1347 = igen_io_fire ? _GEN_323 : rob_payload_66_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1348 = igen_io_fire ? _GEN_324 : rob_payload_67_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1349 = igen_io_fire ? _GEN_325 : rob_payload_68_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1350 = igen_io_fire ? _GEN_326 : rob_payload_69_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1351 = igen_io_fire ? _GEN_327 : rob_payload_70_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1352 = igen_io_fire ? _GEN_328 : rob_payload_71_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1353 = igen_io_fire ? _GEN_329 : rob_payload_72_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1354 = igen_io_fire ? _GEN_330 : rob_payload_73_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1355 = igen_io_fire ? _GEN_331 : rob_payload_74_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1356 = igen_io_fire ? _GEN_332 : rob_payload_75_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1357 = igen_io_fire ? _GEN_333 : rob_payload_76_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1358 = igen_io_fire ? _GEN_334 : rob_payload_77_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1359 = igen_io_fire ? _GEN_335 : rob_payload_78_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1360 = igen_io_fire ? _GEN_336 : rob_payload_79_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1361 = igen_io_fire ? _GEN_337 : rob_payload_80_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1362 = igen_io_fire ? _GEN_338 : rob_payload_81_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1363 = igen_io_fire ? _GEN_339 : rob_payload_82_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1364 = igen_io_fire ? _GEN_340 : rob_payload_83_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1365 = igen_io_fire ? _GEN_341 : rob_payload_84_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1366 = igen_io_fire ? _GEN_342 : rob_payload_85_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1367 = igen_io_fire ? _GEN_343 : rob_payload_86_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1368 = igen_io_fire ? _GEN_344 : rob_payload_87_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1369 = igen_io_fire ? _GEN_345 : rob_payload_88_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1370 = igen_io_fire ? _GEN_346 : rob_payload_89_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1371 = igen_io_fire ? _GEN_347 : rob_payload_90_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1372 = igen_io_fire ? _GEN_348 : rob_payload_91_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1373 = igen_io_fire ? _GEN_349 : rob_payload_92_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1374 = igen_io_fire ? _GEN_350 : rob_payload_93_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1375 = igen_io_fire ? _GEN_351 : rob_payload_94_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1376 = igen_io_fire ? _GEN_352 : rob_payload_95_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1377 = igen_io_fire ? _GEN_353 : rob_payload_96_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1378 = igen_io_fire ? _GEN_354 : rob_payload_97_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1379 = igen_io_fire ? _GEN_355 : rob_payload_98_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1380 = igen_io_fire ? _GEN_356 : rob_payload_99_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1381 = igen_io_fire ? _GEN_357 : rob_payload_100_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1382 = igen_io_fire ? _GEN_358 : rob_payload_101_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1383 = igen_io_fire ? _GEN_359 : rob_payload_102_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1384 = igen_io_fire ? _GEN_360 : rob_payload_103_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1385 = igen_io_fire ? _GEN_361 : rob_payload_104_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1386 = igen_io_fire ? _GEN_362 : rob_payload_105_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1387 = igen_io_fire ? _GEN_363 : rob_payload_106_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1388 = igen_io_fire ? _GEN_364 : rob_payload_107_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1389 = igen_io_fire ? _GEN_365 : rob_payload_108_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1390 = igen_io_fire ? _GEN_366 : rob_payload_109_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1391 = igen_io_fire ? _GEN_367 : rob_payload_110_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1392 = igen_io_fire ? _GEN_368 : rob_payload_111_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1393 = igen_io_fire ? _GEN_369 : rob_payload_112_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1394 = igen_io_fire ? _GEN_370 : rob_payload_113_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1395 = igen_io_fire ? _GEN_371 : rob_payload_114_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1396 = igen_io_fire ? _GEN_372 : rob_payload_115_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1397 = igen_io_fire ? _GEN_373 : rob_payload_116_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1398 = igen_io_fire ? _GEN_374 : rob_payload_117_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1399 = igen_io_fire ? _GEN_375 : rob_payload_118_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1400 = igen_io_fire ? _GEN_376 : rob_payload_119_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1401 = igen_io_fire ? _GEN_377 : rob_payload_120_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1402 = igen_io_fire ? _GEN_378 : rob_payload_121_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1403 = igen_io_fire ? _GEN_379 : rob_payload_122_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1404 = igen_io_fire ? _GEN_380 : rob_payload_123_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1405 = igen_io_fire ? _GEN_381 : rob_payload_124_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1406 = igen_io_fire ? _GEN_382 : rob_payload_125_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1407 = igen_io_fire ? _GEN_383 : rob_payload_126_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1408 = igen_io_fire ? _GEN_384 : rob_payload_127_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [3:0] _GEN_1793 = igen_io_fire ? _GEN_769 : rob_flits_returned_0; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1794 = igen_io_fire ? _GEN_770 : rob_flits_returned_1; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1795 = igen_io_fire ? _GEN_771 : rob_flits_returned_2; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1796 = igen_io_fire ? _GEN_772 : rob_flits_returned_3; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1797 = igen_io_fire ? _GEN_773 : rob_flits_returned_4; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1798 = igen_io_fire ? _GEN_774 : rob_flits_returned_5; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1799 = igen_io_fire ? _GEN_775 : rob_flits_returned_6; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1800 = igen_io_fire ? _GEN_776 : rob_flits_returned_7; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1801 = igen_io_fire ? _GEN_777 : rob_flits_returned_8; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1802 = igen_io_fire ? _GEN_778 : rob_flits_returned_9; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1803 = igen_io_fire ? _GEN_779 : rob_flits_returned_10; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1804 = igen_io_fire ? _GEN_780 : rob_flits_returned_11; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1805 = igen_io_fire ? _GEN_781 : rob_flits_returned_12; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1806 = igen_io_fire ? _GEN_782 : rob_flits_returned_13; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1807 = igen_io_fire ? _GEN_783 : rob_flits_returned_14; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1808 = igen_io_fire ? _GEN_784 : rob_flits_returned_15; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1809 = igen_io_fire ? _GEN_785 : rob_flits_returned_16; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1810 = igen_io_fire ? _GEN_786 : rob_flits_returned_17; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1811 = igen_io_fire ? _GEN_787 : rob_flits_returned_18; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1812 = igen_io_fire ? _GEN_788 : rob_flits_returned_19; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1813 = igen_io_fire ? _GEN_789 : rob_flits_returned_20; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1814 = igen_io_fire ? _GEN_790 : rob_flits_returned_21; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1815 = igen_io_fire ? _GEN_791 : rob_flits_returned_22; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1816 = igen_io_fire ? _GEN_792 : rob_flits_returned_23; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1817 = igen_io_fire ? _GEN_793 : rob_flits_returned_24; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1818 = igen_io_fire ? _GEN_794 : rob_flits_returned_25; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1819 = igen_io_fire ? _GEN_795 : rob_flits_returned_26; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1820 = igen_io_fire ? _GEN_796 : rob_flits_returned_27; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1821 = igen_io_fire ? _GEN_797 : rob_flits_returned_28; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1822 = igen_io_fire ? _GEN_798 : rob_flits_returned_29; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1823 = igen_io_fire ? _GEN_799 : rob_flits_returned_30; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1824 = igen_io_fire ? _GEN_800 : rob_flits_returned_31; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1825 = igen_io_fire ? _GEN_801 : rob_flits_returned_32; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1826 = igen_io_fire ? _GEN_802 : rob_flits_returned_33; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1827 = igen_io_fire ? _GEN_803 : rob_flits_returned_34; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1828 = igen_io_fire ? _GEN_804 : rob_flits_returned_35; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1829 = igen_io_fire ? _GEN_805 : rob_flits_returned_36; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1830 = igen_io_fire ? _GEN_806 : rob_flits_returned_37; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1831 = igen_io_fire ? _GEN_807 : rob_flits_returned_38; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1832 = igen_io_fire ? _GEN_808 : rob_flits_returned_39; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1833 = igen_io_fire ? _GEN_809 : rob_flits_returned_40; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1834 = igen_io_fire ? _GEN_810 : rob_flits_returned_41; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1835 = igen_io_fire ? _GEN_811 : rob_flits_returned_42; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1836 = igen_io_fire ? _GEN_812 : rob_flits_returned_43; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1837 = igen_io_fire ? _GEN_813 : rob_flits_returned_44; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1838 = igen_io_fire ? _GEN_814 : rob_flits_returned_45; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1839 = igen_io_fire ? _GEN_815 : rob_flits_returned_46; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1840 = igen_io_fire ? _GEN_816 : rob_flits_returned_47; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1841 = igen_io_fire ? _GEN_817 : rob_flits_returned_48; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1842 = igen_io_fire ? _GEN_818 : rob_flits_returned_49; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1843 = igen_io_fire ? _GEN_819 : rob_flits_returned_50; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1844 = igen_io_fire ? _GEN_820 : rob_flits_returned_51; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1845 = igen_io_fire ? _GEN_821 : rob_flits_returned_52; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1846 = igen_io_fire ? _GEN_822 : rob_flits_returned_53; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1847 = igen_io_fire ? _GEN_823 : rob_flits_returned_54; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1848 = igen_io_fire ? _GEN_824 : rob_flits_returned_55; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1849 = igen_io_fire ? _GEN_825 : rob_flits_returned_56; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1850 = igen_io_fire ? _GEN_826 : rob_flits_returned_57; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1851 = igen_io_fire ? _GEN_827 : rob_flits_returned_58; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1852 = igen_io_fire ? _GEN_828 : rob_flits_returned_59; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1853 = igen_io_fire ? _GEN_829 : rob_flits_returned_60; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1854 = igen_io_fire ? _GEN_830 : rob_flits_returned_61; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1855 = igen_io_fire ? _GEN_831 : rob_flits_returned_62; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1856 = igen_io_fire ? _GEN_832 : rob_flits_returned_63; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1857 = igen_io_fire ? _GEN_833 : rob_flits_returned_64; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1858 = igen_io_fire ? _GEN_834 : rob_flits_returned_65; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1859 = igen_io_fire ? _GEN_835 : rob_flits_returned_66; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1860 = igen_io_fire ? _GEN_836 : rob_flits_returned_67; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1861 = igen_io_fire ? _GEN_837 : rob_flits_returned_68; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1862 = igen_io_fire ? _GEN_838 : rob_flits_returned_69; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1863 = igen_io_fire ? _GEN_839 : rob_flits_returned_70; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1864 = igen_io_fire ? _GEN_840 : rob_flits_returned_71; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1865 = igen_io_fire ? _GEN_841 : rob_flits_returned_72; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1866 = igen_io_fire ? _GEN_842 : rob_flits_returned_73; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1867 = igen_io_fire ? _GEN_843 : rob_flits_returned_74; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1868 = igen_io_fire ? _GEN_844 : rob_flits_returned_75; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1869 = igen_io_fire ? _GEN_845 : rob_flits_returned_76; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1870 = igen_io_fire ? _GEN_846 : rob_flits_returned_77; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1871 = igen_io_fire ? _GEN_847 : rob_flits_returned_78; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1872 = igen_io_fire ? _GEN_848 : rob_flits_returned_79; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1873 = igen_io_fire ? _GEN_849 : rob_flits_returned_80; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1874 = igen_io_fire ? _GEN_850 : rob_flits_returned_81; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1875 = igen_io_fire ? _GEN_851 : rob_flits_returned_82; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1876 = igen_io_fire ? _GEN_852 : rob_flits_returned_83; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1877 = igen_io_fire ? _GEN_853 : rob_flits_returned_84; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1878 = igen_io_fire ? _GEN_854 : rob_flits_returned_85; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1879 = igen_io_fire ? _GEN_855 : rob_flits_returned_86; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1880 = igen_io_fire ? _GEN_856 : rob_flits_returned_87; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1881 = igen_io_fire ? _GEN_857 : rob_flits_returned_88; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1882 = igen_io_fire ? _GEN_858 : rob_flits_returned_89; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1883 = igen_io_fire ? _GEN_859 : rob_flits_returned_90; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1884 = igen_io_fire ? _GEN_860 : rob_flits_returned_91; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1885 = igen_io_fire ? _GEN_861 : rob_flits_returned_92; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1886 = igen_io_fire ? _GEN_862 : rob_flits_returned_93; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1887 = igen_io_fire ? _GEN_863 : rob_flits_returned_94; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1888 = igen_io_fire ? _GEN_864 : rob_flits_returned_95; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1889 = igen_io_fire ? _GEN_865 : rob_flits_returned_96; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1890 = igen_io_fire ? _GEN_866 : rob_flits_returned_97; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1891 = igen_io_fire ? _GEN_867 : rob_flits_returned_98; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1892 = igen_io_fire ? _GEN_868 : rob_flits_returned_99; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1893 = igen_io_fire ? _GEN_869 : rob_flits_returned_100; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1894 = igen_io_fire ? _GEN_870 : rob_flits_returned_101; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1895 = igen_io_fire ? _GEN_871 : rob_flits_returned_102; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1896 = igen_io_fire ? _GEN_872 : rob_flits_returned_103; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1897 = igen_io_fire ? _GEN_873 : rob_flits_returned_104; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1898 = igen_io_fire ? _GEN_874 : rob_flits_returned_105; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1899 = igen_io_fire ? _GEN_875 : rob_flits_returned_106; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1900 = igen_io_fire ? _GEN_876 : rob_flits_returned_107; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1901 = igen_io_fire ? _GEN_877 : rob_flits_returned_108; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1902 = igen_io_fire ? _GEN_878 : rob_flits_returned_109; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1903 = igen_io_fire ? _GEN_879 : rob_flits_returned_110; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1904 = igen_io_fire ? _GEN_880 : rob_flits_returned_111; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1905 = igen_io_fire ? _GEN_881 : rob_flits_returned_112; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1906 = igen_io_fire ? _GEN_882 : rob_flits_returned_113; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1907 = igen_io_fire ? _GEN_883 : rob_flits_returned_114; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1908 = igen_io_fire ? _GEN_884 : rob_flits_returned_115; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1909 = igen_io_fire ? _GEN_885 : rob_flits_returned_116; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1910 = igen_io_fire ? _GEN_886 : rob_flits_returned_117; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1911 = igen_io_fire ? _GEN_887 : rob_flits_returned_118; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1912 = igen_io_fire ? _GEN_888 : rob_flits_returned_119; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1913 = igen_io_fire ? _GEN_889 : rob_flits_returned_120; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1914 = igen_io_fire ? _GEN_890 : rob_flits_returned_121; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1915 = igen_io_fire ? _GEN_891 : rob_flits_returned_122; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1916 = igen_io_fire ? _GEN_892 : rob_flits_returned_123; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1917 = igen_io_fire ? _GEN_893 : rob_flits_returned_124; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1918 = igen_io_fire ? _GEN_894 : rob_flits_returned_125; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1919 = igen_io_fire ? _GEN_895 : rob_flits_returned_126; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1920 = igen_io_fire ? _GEN_896 : rob_flits_returned_127; // @[TestHarness.scala 178:25 154:31]
  wire  enable_print_latency = plusarg_reader_out; // @[TestHarness.scala 190:81]
  wire [31:0] out_payload_tsc = io_from_noc_0_flit_bits_payload[63:32]; // @[TestHarness.scala 194:51]
  reg  packet_valid; // @[TestHarness.scala 196:31]
  reg [6:0] packet_rob_idx; // @[TestHarness.scala 197:29]
  wire [127:0] _T_25 = rob_valids >> out_payload_rob_idx; // @[TestHarness.scala 201:24]
  wire [31:0] _GEN_2050 = 7'h1 == out_payload_rob_idx[6:0] ? rob_payload_1_tsc : rob_payload_0_tsc; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2051 = 7'h2 == out_payload_rob_idx[6:0] ? rob_payload_2_tsc : _GEN_2050; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2052 = 7'h3 == out_payload_rob_idx[6:0] ? rob_payload_3_tsc : _GEN_2051; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2053 = 7'h4 == out_payload_rob_idx[6:0] ? rob_payload_4_tsc : _GEN_2052; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2054 = 7'h5 == out_payload_rob_idx[6:0] ? rob_payload_5_tsc : _GEN_2053; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2055 = 7'h6 == out_payload_rob_idx[6:0] ? rob_payload_6_tsc : _GEN_2054; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2056 = 7'h7 == out_payload_rob_idx[6:0] ? rob_payload_7_tsc : _GEN_2055; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2057 = 7'h8 == out_payload_rob_idx[6:0] ? rob_payload_8_tsc : _GEN_2056; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2058 = 7'h9 == out_payload_rob_idx[6:0] ? rob_payload_9_tsc : _GEN_2057; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2059 = 7'ha == out_payload_rob_idx[6:0] ? rob_payload_10_tsc : _GEN_2058; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2060 = 7'hb == out_payload_rob_idx[6:0] ? rob_payload_11_tsc : _GEN_2059; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2061 = 7'hc == out_payload_rob_idx[6:0] ? rob_payload_12_tsc : _GEN_2060; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2062 = 7'hd == out_payload_rob_idx[6:0] ? rob_payload_13_tsc : _GEN_2061; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2063 = 7'he == out_payload_rob_idx[6:0] ? rob_payload_14_tsc : _GEN_2062; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2064 = 7'hf == out_payload_rob_idx[6:0] ? rob_payload_15_tsc : _GEN_2063; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2065 = 7'h10 == out_payload_rob_idx[6:0] ? rob_payload_16_tsc : _GEN_2064; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2066 = 7'h11 == out_payload_rob_idx[6:0] ? rob_payload_17_tsc : _GEN_2065; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2067 = 7'h12 == out_payload_rob_idx[6:0] ? rob_payload_18_tsc : _GEN_2066; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2068 = 7'h13 == out_payload_rob_idx[6:0] ? rob_payload_19_tsc : _GEN_2067; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2069 = 7'h14 == out_payload_rob_idx[6:0] ? rob_payload_20_tsc : _GEN_2068; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2070 = 7'h15 == out_payload_rob_idx[6:0] ? rob_payload_21_tsc : _GEN_2069; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2071 = 7'h16 == out_payload_rob_idx[6:0] ? rob_payload_22_tsc : _GEN_2070; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2072 = 7'h17 == out_payload_rob_idx[6:0] ? rob_payload_23_tsc : _GEN_2071; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2073 = 7'h18 == out_payload_rob_idx[6:0] ? rob_payload_24_tsc : _GEN_2072; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2074 = 7'h19 == out_payload_rob_idx[6:0] ? rob_payload_25_tsc : _GEN_2073; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2075 = 7'h1a == out_payload_rob_idx[6:0] ? rob_payload_26_tsc : _GEN_2074; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2076 = 7'h1b == out_payload_rob_idx[6:0] ? rob_payload_27_tsc : _GEN_2075; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2077 = 7'h1c == out_payload_rob_idx[6:0] ? rob_payload_28_tsc : _GEN_2076; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2078 = 7'h1d == out_payload_rob_idx[6:0] ? rob_payload_29_tsc : _GEN_2077; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2079 = 7'h1e == out_payload_rob_idx[6:0] ? rob_payload_30_tsc : _GEN_2078; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2080 = 7'h1f == out_payload_rob_idx[6:0] ? rob_payload_31_tsc : _GEN_2079; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2081 = 7'h20 == out_payload_rob_idx[6:0] ? rob_payload_32_tsc : _GEN_2080; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2082 = 7'h21 == out_payload_rob_idx[6:0] ? rob_payload_33_tsc : _GEN_2081; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2083 = 7'h22 == out_payload_rob_idx[6:0] ? rob_payload_34_tsc : _GEN_2082; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2084 = 7'h23 == out_payload_rob_idx[6:0] ? rob_payload_35_tsc : _GEN_2083; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2085 = 7'h24 == out_payload_rob_idx[6:0] ? rob_payload_36_tsc : _GEN_2084; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2086 = 7'h25 == out_payload_rob_idx[6:0] ? rob_payload_37_tsc : _GEN_2085; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2087 = 7'h26 == out_payload_rob_idx[6:0] ? rob_payload_38_tsc : _GEN_2086; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2088 = 7'h27 == out_payload_rob_idx[6:0] ? rob_payload_39_tsc : _GEN_2087; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2089 = 7'h28 == out_payload_rob_idx[6:0] ? rob_payload_40_tsc : _GEN_2088; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2090 = 7'h29 == out_payload_rob_idx[6:0] ? rob_payload_41_tsc : _GEN_2089; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2091 = 7'h2a == out_payload_rob_idx[6:0] ? rob_payload_42_tsc : _GEN_2090; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2092 = 7'h2b == out_payload_rob_idx[6:0] ? rob_payload_43_tsc : _GEN_2091; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2093 = 7'h2c == out_payload_rob_idx[6:0] ? rob_payload_44_tsc : _GEN_2092; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2094 = 7'h2d == out_payload_rob_idx[6:0] ? rob_payload_45_tsc : _GEN_2093; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2095 = 7'h2e == out_payload_rob_idx[6:0] ? rob_payload_46_tsc : _GEN_2094; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2096 = 7'h2f == out_payload_rob_idx[6:0] ? rob_payload_47_tsc : _GEN_2095; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2097 = 7'h30 == out_payload_rob_idx[6:0] ? rob_payload_48_tsc : _GEN_2096; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2098 = 7'h31 == out_payload_rob_idx[6:0] ? rob_payload_49_tsc : _GEN_2097; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2099 = 7'h32 == out_payload_rob_idx[6:0] ? rob_payload_50_tsc : _GEN_2098; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2100 = 7'h33 == out_payload_rob_idx[6:0] ? rob_payload_51_tsc : _GEN_2099; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2101 = 7'h34 == out_payload_rob_idx[6:0] ? rob_payload_52_tsc : _GEN_2100; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2102 = 7'h35 == out_payload_rob_idx[6:0] ? rob_payload_53_tsc : _GEN_2101; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2103 = 7'h36 == out_payload_rob_idx[6:0] ? rob_payload_54_tsc : _GEN_2102; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2104 = 7'h37 == out_payload_rob_idx[6:0] ? rob_payload_55_tsc : _GEN_2103; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2105 = 7'h38 == out_payload_rob_idx[6:0] ? rob_payload_56_tsc : _GEN_2104; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2106 = 7'h39 == out_payload_rob_idx[6:0] ? rob_payload_57_tsc : _GEN_2105; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2107 = 7'h3a == out_payload_rob_idx[6:0] ? rob_payload_58_tsc : _GEN_2106; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2108 = 7'h3b == out_payload_rob_idx[6:0] ? rob_payload_59_tsc : _GEN_2107; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2109 = 7'h3c == out_payload_rob_idx[6:0] ? rob_payload_60_tsc : _GEN_2108; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2110 = 7'h3d == out_payload_rob_idx[6:0] ? rob_payload_61_tsc : _GEN_2109; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2111 = 7'h3e == out_payload_rob_idx[6:0] ? rob_payload_62_tsc : _GEN_2110; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2112 = 7'h3f == out_payload_rob_idx[6:0] ? rob_payload_63_tsc : _GEN_2111; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2113 = 7'h40 == out_payload_rob_idx[6:0] ? rob_payload_64_tsc : _GEN_2112; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2114 = 7'h41 == out_payload_rob_idx[6:0] ? rob_payload_65_tsc : _GEN_2113; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2115 = 7'h42 == out_payload_rob_idx[6:0] ? rob_payload_66_tsc : _GEN_2114; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2116 = 7'h43 == out_payload_rob_idx[6:0] ? rob_payload_67_tsc : _GEN_2115; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2117 = 7'h44 == out_payload_rob_idx[6:0] ? rob_payload_68_tsc : _GEN_2116; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2118 = 7'h45 == out_payload_rob_idx[6:0] ? rob_payload_69_tsc : _GEN_2117; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2119 = 7'h46 == out_payload_rob_idx[6:0] ? rob_payload_70_tsc : _GEN_2118; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2120 = 7'h47 == out_payload_rob_idx[6:0] ? rob_payload_71_tsc : _GEN_2119; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2121 = 7'h48 == out_payload_rob_idx[6:0] ? rob_payload_72_tsc : _GEN_2120; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2122 = 7'h49 == out_payload_rob_idx[6:0] ? rob_payload_73_tsc : _GEN_2121; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2123 = 7'h4a == out_payload_rob_idx[6:0] ? rob_payload_74_tsc : _GEN_2122; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2124 = 7'h4b == out_payload_rob_idx[6:0] ? rob_payload_75_tsc : _GEN_2123; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2125 = 7'h4c == out_payload_rob_idx[6:0] ? rob_payload_76_tsc : _GEN_2124; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2126 = 7'h4d == out_payload_rob_idx[6:0] ? rob_payload_77_tsc : _GEN_2125; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2127 = 7'h4e == out_payload_rob_idx[6:0] ? rob_payload_78_tsc : _GEN_2126; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2128 = 7'h4f == out_payload_rob_idx[6:0] ? rob_payload_79_tsc : _GEN_2127; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2129 = 7'h50 == out_payload_rob_idx[6:0] ? rob_payload_80_tsc : _GEN_2128; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2130 = 7'h51 == out_payload_rob_idx[6:0] ? rob_payload_81_tsc : _GEN_2129; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2131 = 7'h52 == out_payload_rob_idx[6:0] ? rob_payload_82_tsc : _GEN_2130; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2132 = 7'h53 == out_payload_rob_idx[6:0] ? rob_payload_83_tsc : _GEN_2131; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2133 = 7'h54 == out_payload_rob_idx[6:0] ? rob_payload_84_tsc : _GEN_2132; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2134 = 7'h55 == out_payload_rob_idx[6:0] ? rob_payload_85_tsc : _GEN_2133; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2135 = 7'h56 == out_payload_rob_idx[6:0] ? rob_payload_86_tsc : _GEN_2134; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2136 = 7'h57 == out_payload_rob_idx[6:0] ? rob_payload_87_tsc : _GEN_2135; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2137 = 7'h58 == out_payload_rob_idx[6:0] ? rob_payload_88_tsc : _GEN_2136; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2138 = 7'h59 == out_payload_rob_idx[6:0] ? rob_payload_89_tsc : _GEN_2137; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2139 = 7'h5a == out_payload_rob_idx[6:0] ? rob_payload_90_tsc : _GEN_2138; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2140 = 7'h5b == out_payload_rob_idx[6:0] ? rob_payload_91_tsc : _GEN_2139; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2141 = 7'h5c == out_payload_rob_idx[6:0] ? rob_payload_92_tsc : _GEN_2140; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2142 = 7'h5d == out_payload_rob_idx[6:0] ? rob_payload_93_tsc : _GEN_2141; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2143 = 7'h5e == out_payload_rob_idx[6:0] ? rob_payload_94_tsc : _GEN_2142; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2144 = 7'h5f == out_payload_rob_idx[6:0] ? rob_payload_95_tsc : _GEN_2143; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2145 = 7'h60 == out_payload_rob_idx[6:0] ? rob_payload_96_tsc : _GEN_2144; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2146 = 7'h61 == out_payload_rob_idx[6:0] ? rob_payload_97_tsc : _GEN_2145; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2147 = 7'h62 == out_payload_rob_idx[6:0] ? rob_payload_98_tsc : _GEN_2146; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2148 = 7'h63 == out_payload_rob_idx[6:0] ? rob_payload_99_tsc : _GEN_2147; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2149 = 7'h64 == out_payload_rob_idx[6:0] ? rob_payload_100_tsc : _GEN_2148; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2150 = 7'h65 == out_payload_rob_idx[6:0] ? rob_payload_101_tsc : _GEN_2149; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2151 = 7'h66 == out_payload_rob_idx[6:0] ? rob_payload_102_tsc : _GEN_2150; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2152 = 7'h67 == out_payload_rob_idx[6:0] ? rob_payload_103_tsc : _GEN_2151; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2153 = 7'h68 == out_payload_rob_idx[6:0] ? rob_payload_104_tsc : _GEN_2152; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2154 = 7'h69 == out_payload_rob_idx[6:0] ? rob_payload_105_tsc : _GEN_2153; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2155 = 7'h6a == out_payload_rob_idx[6:0] ? rob_payload_106_tsc : _GEN_2154; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2156 = 7'h6b == out_payload_rob_idx[6:0] ? rob_payload_107_tsc : _GEN_2155; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2157 = 7'h6c == out_payload_rob_idx[6:0] ? rob_payload_108_tsc : _GEN_2156; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2158 = 7'h6d == out_payload_rob_idx[6:0] ? rob_payload_109_tsc : _GEN_2157; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2159 = 7'h6e == out_payload_rob_idx[6:0] ? rob_payload_110_tsc : _GEN_2158; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2160 = 7'h6f == out_payload_rob_idx[6:0] ? rob_payload_111_tsc : _GEN_2159; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2161 = 7'h70 == out_payload_rob_idx[6:0] ? rob_payload_112_tsc : _GEN_2160; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2162 = 7'h71 == out_payload_rob_idx[6:0] ? rob_payload_113_tsc : _GEN_2161; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2163 = 7'h72 == out_payload_rob_idx[6:0] ? rob_payload_114_tsc : _GEN_2162; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2164 = 7'h73 == out_payload_rob_idx[6:0] ? rob_payload_115_tsc : _GEN_2163; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2165 = 7'h74 == out_payload_rob_idx[6:0] ? rob_payload_116_tsc : _GEN_2164; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2166 = 7'h75 == out_payload_rob_idx[6:0] ? rob_payload_117_tsc : _GEN_2165; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2167 = 7'h76 == out_payload_rob_idx[6:0] ? rob_payload_118_tsc : _GEN_2166; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2168 = 7'h77 == out_payload_rob_idx[6:0] ? rob_payload_119_tsc : _GEN_2167; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2169 = 7'h78 == out_payload_rob_idx[6:0] ? rob_payload_120_tsc : _GEN_2168; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2170 = 7'h79 == out_payload_rob_idx[6:0] ? rob_payload_121_tsc : _GEN_2169; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2171 = 7'h7a == out_payload_rob_idx[6:0] ? rob_payload_122_tsc : _GEN_2170; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2172 = 7'h7b == out_payload_rob_idx[6:0] ? rob_payload_123_tsc : _GEN_2171; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2173 = 7'h7c == out_payload_rob_idx[6:0] ? rob_payload_124_tsc : _GEN_2172; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2174 = 7'h7d == out_payload_rob_idx[6:0] ? rob_payload_125_tsc : _GEN_2173; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2175 = 7'h7e == out_payload_rob_idx[6:0] ? rob_payload_126_tsc : _GEN_2174; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_2176 = 7'h7f == out_payload_rob_idx[6:0] ? rob_payload_127_tsc : _GEN_2175; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2178 = 7'h1 == out_payload_rob_idx[6:0] ? rob_payload_1_rob_idx : rob_payload_0_rob_idx; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2179 = 7'h2 == out_payload_rob_idx[6:0] ? rob_payload_2_rob_idx : _GEN_2178; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2180 = 7'h3 == out_payload_rob_idx[6:0] ? rob_payload_3_rob_idx : _GEN_2179; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2181 = 7'h4 == out_payload_rob_idx[6:0] ? rob_payload_4_rob_idx : _GEN_2180; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2182 = 7'h5 == out_payload_rob_idx[6:0] ? rob_payload_5_rob_idx : _GEN_2181; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2183 = 7'h6 == out_payload_rob_idx[6:0] ? rob_payload_6_rob_idx : _GEN_2182; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2184 = 7'h7 == out_payload_rob_idx[6:0] ? rob_payload_7_rob_idx : _GEN_2183; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2185 = 7'h8 == out_payload_rob_idx[6:0] ? rob_payload_8_rob_idx : _GEN_2184; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2186 = 7'h9 == out_payload_rob_idx[6:0] ? rob_payload_9_rob_idx : _GEN_2185; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2187 = 7'ha == out_payload_rob_idx[6:0] ? rob_payload_10_rob_idx : _GEN_2186; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2188 = 7'hb == out_payload_rob_idx[6:0] ? rob_payload_11_rob_idx : _GEN_2187; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2189 = 7'hc == out_payload_rob_idx[6:0] ? rob_payload_12_rob_idx : _GEN_2188; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2190 = 7'hd == out_payload_rob_idx[6:0] ? rob_payload_13_rob_idx : _GEN_2189; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2191 = 7'he == out_payload_rob_idx[6:0] ? rob_payload_14_rob_idx : _GEN_2190; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2192 = 7'hf == out_payload_rob_idx[6:0] ? rob_payload_15_rob_idx : _GEN_2191; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2193 = 7'h10 == out_payload_rob_idx[6:0] ? rob_payload_16_rob_idx : _GEN_2192; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2194 = 7'h11 == out_payload_rob_idx[6:0] ? rob_payload_17_rob_idx : _GEN_2193; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2195 = 7'h12 == out_payload_rob_idx[6:0] ? rob_payload_18_rob_idx : _GEN_2194; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2196 = 7'h13 == out_payload_rob_idx[6:0] ? rob_payload_19_rob_idx : _GEN_2195; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2197 = 7'h14 == out_payload_rob_idx[6:0] ? rob_payload_20_rob_idx : _GEN_2196; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2198 = 7'h15 == out_payload_rob_idx[6:0] ? rob_payload_21_rob_idx : _GEN_2197; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2199 = 7'h16 == out_payload_rob_idx[6:0] ? rob_payload_22_rob_idx : _GEN_2198; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2200 = 7'h17 == out_payload_rob_idx[6:0] ? rob_payload_23_rob_idx : _GEN_2199; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2201 = 7'h18 == out_payload_rob_idx[6:0] ? rob_payload_24_rob_idx : _GEN_2200; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2202 = 7'h19 == out_payload_rob_idx[6:0] ? rob_payload_25_rob_idx : _GEN_2201; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2203 = 7'h1a == out_payload_rob_idx[6:0] ? rob_payload_26_rob_idx : _GEN_2202; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2204 = 7'h1b == out_payload_rob_idx[6:0] ? rob_payload_27_rob_idx : _GEN_2203; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2205 = 7'h1c == out_payload_rob_idx[6:0] ? rob_payload_28_rob_idx : _GEN_2204; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2206 = 7'h1d == out_payload_rob_idx[6:0] ? rob_payload_29_rob_idx : _GEN_2205; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2207 = 7'h1e == out_payload_rob_idx[6:0] ? rob_payload_30_rob_idx : _GEN_2206; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2208 = 7'h1f == out_payload_rob_idx[6:0] ? rob_payload_31_rob_idx : _GEN_2207; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2209 = 7'h20 == out_payload_rob_idx[6:0] ? rob_payload_32_rob_idx : _GEN_2208; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2210 = 7'h21 == out_payload_rob_idx[6:0] ? rob_payload_33_rob_idx : _GEN_2209; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2211 = 7'h22 == out_payload_rob_idx[6:0] ? rob_payload_34_rob_idx : _GEN_2210; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2212 = 7'h23 == out_payload_rob_idx[6:0] ? rob_payload_35_rob_idx : _GEN_2211; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2213 = 7'h24 == out_payload_rob_idx[6:0] ? rob_payload_36_rob_idx : _GEN_2212; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2214 = 7'h25 == out_payload_rob_idx[6:0] ? rob_payload_37_rob_idx : _GEN_2213; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2215 = 7'h26 == out_payload_rob_idx[6:0] ? rob_payload_38_rob_idx : _GEN_2214; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2216 = 7'h27 == out_payload_rob_idx[6:0] ? rob_payload_39_rob_idx : _GEN_2215; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2217 = 7'h28 == out_payload_rob_idx[6:0] ? rob_payload_40_rob_idx : _GEN_2216; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2218 = 7'h29 == out_payload_rob_idx[6:0] ? rob_payload_41_rob_idx : _GEN_2217; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2219 = 7'h2a == out_payload_rob_idx[6:0] ? rob_payload_42_rob_idx : _GEN_2218; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2220 = 7'h2b == out_payload_rob_idx[6:0] ? rob_payload_43_rob_idx : _GEN_2219; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2221 = 7'h2c == out_payload_rob_idx[6:0] ? rob_payload_44_rob_idx : _GEN_2220; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2222 = 7'h2d == out_payload_rob_idx[6:0] ? rob_payload_45_rob_idx : _GEN_2221; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2223 = 7'h2e == out_payload_rob_idx[6:0] ? rob_payload_46_rob_idx : _GEN_2222; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2224 = 7'h2f == out_payload_rob_idx[6:0] ? rob_payload_47_rob_idx : _GEN_2223; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2225 = 7'h30 == out_payload_rob_idx[6:0] ? rob_payload_48_rob_idx : _GEN_2224; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2226 = 7'h31 == out_payload_rob_idx[6:0] ? rob_payload_49_rob_idx : _GEN_2225; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2227 = 7'h32 == out_payload_rob_idx[6:0] ? rob_payload_50_rob_idx : _GEN_2226; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2228 = 7'h33 == out_payload_rob_idx[6:0] ? rob_payload_51_rob_idx : _GEN_2227; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2229 = 7'h34 == out_payload_rob_idx[6:0] ? rob_payload_52_rob_idx : _GEN_2228; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2230 = 7'h35 == out_payload_rob_idx[6:0] ? rob_payload_53_rob_idx : _GEN_2229; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2231 = 7'h36 == out_payload_rob_idx[6:0] ? rob_payload_54_rob_idx : _GEN_2230; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2232 = 7'h37 == out_payload_rob_idx[6:0] ? rob_payload_55_rob_idx : _GEN_2231; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2233 = 7'h38 == out_payload_rob_idx[6:0] ? rob_payload_56_rob_idx : _GEN_2232; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2234 = 7'h39 == out_payload_rob_idx[6:0] ? rob_payload_57_rob_idx : _GEN_2233; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2235 = 7'h3a == out_payload_rob_idx[6:0] ? rob_payload_58_rob_idx : _GEN_2234; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2236 = 7'h3b == out_payload_rob_idx[6:0] ? rob_payload_59_rob_idx : _GEN_2235; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2237 = 7'h3c == out_payload_rob_idx[6:0] ? rob_payload_60_rob_idx : _GEN_2236; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2238 = 7'h3d == out_payload_rob_idx[6:0] ? rob_payload_61_rob_idx : _GEN_2237; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2239 = 7'h3e == out_payload_rob_idx[6:0] ? rob_payload_62_rob_idx : _GEN_2238; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2240 = 7'h3f == out_payload_rob_idx[6:0] ? rob_payload_63_rob_idx : _GEN_2239; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2241 = 7'h40 == out_payload_rob_idx[6:0] ? rob_payload_64_rob_idx : _GEN_2240; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2242 = 7'h41 == out_payload_rob_idx[6:0] ? rob_payload_65_rob_idx : _GEN_2241; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2243 = 7'h42 == out_payload_rob_idx[6:0] ? rob_payload_66_rob_idx : _GEN_2242; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2244 = 7'h43 == out_payload_rob_idx[6:0] ? rob_payload_67_rob_idx : _GEN_2243; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2245 = 7'h44 == out_payload_rob_idx[6:0] ? rob_payload_68_rob_idx : _GEN_2244; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2246 = 7'h45 == out_payload_rob_idx[6:0] ? rob_payload_69_rob_idx : _GEN_2245; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2247 = 7'h46 == out_payload_rob_idx[6:0] ? rob_payload_70_rob_idx : _GEN_2246; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2248 = 7'h47 == out_payload_rob_idx[6:0] ? rob_payload_71_rob_idx : _GEN_2247; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2249 = 7'h48 == out_payload_rob_idx[6:0] ? rob_payload_72_rob_idx : _GEN_2248; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2250 = 7'h49 == out_payload_rob_idx[6:0] ? rob_payload_73_rob_idx : _GEN_2249; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2251 = 7'h4a == out_payload_rob_idx[6:0] ? rob_payload_74_rob_idx : _GEN_2250; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2252 = 7'h4b == out_payload_rob_idx[6:0] ? rob_payload_75_rob_idx : _GEN_2251; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2253 = 7'h4c == out_payload_rob_idx[6:0] ? rob_payload_76_rob_idx : _GEN_2252; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2254 = 7'h4d == out_payload_rob_idx[6:0] ? rob_payload_77_rob_idx : _GEN_2253; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2255 = 7'h4e == out_payload_rob_idx[6:0] ? rob_payload_78_rob_idx : _GEN_2254; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2256 = 7'h4f == out_payload_rob_idx[6:0] ? rob_payload_79_rob_idx : _GEN_2255; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2257 = 7'h50 == out_payload_rob_idx[6:0] ? rob_payload_80_rob_idx : _GEN_2256; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2258 = 7'h51 == out_payload_rob_idx[6:0] ? rob_payload_81_rob_idx : _GEN_2257; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2259 = 7'h52 == out_payload_rob_idx[6:0] ? rob_payload_82_rob_idx : _GEN_2258; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2260 = 7'h53 == out_payload_rob_idx[6:0] ? rob_payload_83_rob_idx : _GEN_2259; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2261 = 7'h54 == out_payload_rob_idx[6:0] ? rob_payload_84_rob_idx : _GEN_2260; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2262 = 7'h55 == out_payload_rob_idx[6:0] ? rob_payload_85_rob_idx : _GEN_2261; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2263 = 7'h56 == out_payload_rob_idx[6:0] ? rob_payload_86_rob_idx : _GEN_2262; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2264 = 7'h57 == out_payload_rob_idx[6:0] ? rob_payload_87_rob_idx : _GEN_2263; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2265 = 7'h58 == out_payload_rob_idx[6:0] ? rob_payload_88_rob_idx : _GEN_2264; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2266 = 7'h59 == out_payload_rob_idx[6:0] ? rob_payload_89_rob_idx : _GEN_2265; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2267 = 7'h5a == out_payload_rob_idx[6:0] ? rob_payload_90_rob_idx : _GEN_2266; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2268 = 7'h5b == out_payload_rob_idx[6:0] ? rob_payload_91_rob_idx : _GEN_2267; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2269 = 7'h5c == out_payload_rob_idx[6:0] ? rob_payload_92_rob_idx : _GEN_2268; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2270 = 7'h5d == out_payload_rob_idx[6:0] ? rob_payload_93_rob_idx : _GEN_2269; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2271 = 7'h5e == out_payload_rob_idx[6:0] ? rob_payload_94_rob_idx : _GEN_2270; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2272 = 7'h5f == out_payload_rob_idx[6:0] ? rob_payload_95_rob_idx : _GEN_2271; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2273 = 7'h60 == out_payload_rob_idx[6:0] ? rob_payload_96_rob_idx : _GEN_2272; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2274 = 7'h61 == out_payload_rob_idx[6:0] ? rob_payload_97_rob_idx : _GEN_2273; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2275 = 7'h62 == out_payload_rob_idx[6:0] ? rob_payload_98_rob_idx : _GEN_2274; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2276 = 7'h63 == out_payload_rob_idx[6:0] ? rob_payload_99_rob_idx : _GEN_2275; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2277 = 7'h64 == out_payload_rob_idx[6:0] ? rob_payload_100_rob_idx : _GEN_2276; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2278 = 7'h65 == out_payload_rob_idx[6:0] ? rob_payload_101_rob_idx : _GEN_2277; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2279 = 7'h66 == out_payload_rob_idx[6:0] ? rob_payload_102_rob_idx : _GEN_2278; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2280 = 7'h67 == out_payload_rob_idx[6:0] ? rob_payload_103_rob_idx : _GEN_2279; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2281 = 7'h68 == out_payload_rob_idx[6:0] ? rob_payload_104_rob_idx : _GEN_2280; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2282 = 7'h69 == out_payload_rob_idx[6:0] ? rob_payload_105_rob_idx : _GEN_2281; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2283 = 7'h6a == out_payload_rob_idx[6:0] ? rob_payload_106_rob_idx : _GEN_2282; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2284 = 7'h6b == out_payload_rob_idx[6:0] ? rob_payload_107_rob_idx : _GEN_2283; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2285 = 7'h6c == out_payload_rob_idx[6:0] ? rob_payload_108_rob_idx : _GEN_2284; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2286 = 7'h6d == out_payload_rob_idx[6:0] ? rob_payload_109_rob_idx : _GEN_2285; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2287 = 7'h6e == out_payload_rob_idx[6:0] ? rob_payload_110_rob_idx : _GEN_2286; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2288 = 7'h6f == out_payload_rob_idx[6:0] ? rob_payload_111_rob_idx : _GEN_2287; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2289 = 7'h70 == out_payload_rob_idx[6:0] ? rob_payload_112_rob_idx : _GEN_2288; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2290 = 7'h71 == out_payload_rob_idx[6:0] ? rob_payload_113_rob_idx : _GEN_2289; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2291 = 7'h72 == out_payload_rob_idx[6:0] ? rob_payload_114_rob_idx : _GEN_2290; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2292 = 7'h73 == out_payload_rob_idx[6:0] ? rob_payload_115_rob_idx : _GEN_2291; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2293 = 7'h74 == out_payload_rob_idx[6:0] ? rob_payload_116_rob_idx : _GEN_2292; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2294 = 7'h75 == out_payload_rob_idx[6:0] ? rob_payload_117_rob_idx : _GEN_2293; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2295 = 7'h76 == out_payload_rob_idx[6:0] ? rob_payload_118_rob_idx : _GEN_2294; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2296 = 7'h77 == out_payload_rob_idx[6:0] ? rob_payload_119_rob_idx : _GEN_2295; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2297 = 7'h78 == out_payload_rob_idx[6:0] ? rob_payload_120_rob_idx : _GEN_2296; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2298 = 7'h79 == out_payload_rob_idx[6:0] ? rob_payload_121_rob_idx : _GEN_2297; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2299 = 7'h7a == out_payload_rob_idx[6:0] ? rob_payload_122_rob_idx : _GEN_2298; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2300 = 7'h7b == out_payload_rob_idx[6:0] ? rob_payload_123_rob_idx : _GEN_2299; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2301 = 7'h7c == out_payload_rob_idx[6:0] ? rob_payload_124_rob_idx : _GEN_2300; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2302 = 7'h7d == out_payload_rob_idx[6:0] ? rob_payload_125_rob_idx : _GEN_2301; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2303 = 7'h7e == out_payload_rob_idx[6:0] ? rob_payload_126_rob_idx : _GEN_2302; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2304 = 7'h7f == out_payload_rob_idx[6:0] ? rob_payload_127_rob_idx : _GEN_2303; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2306 = 7'h1 == out_payload_rob_idx[6:0] ? rob_payload_1_flits_fired : rob_payload_0_flits_fired; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2307 = 7'h2 == out_payload_rob_idx[6:0] ? rob_payload_2_flits_fired : _GEN_2306; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2308 = 7'h3 == out_payload_rob_idx[6:0] ? rob_payload_3_flits_fired : _GEN_2307; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2309 = 7'h4 == out_payload_rob_idx[6:0] ? rob_payload_4_flits_fired : _GEN_2308; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2310 = 7'h5 == out_payload_rob_idx[6:0] ? rob_payload_5_flits_fired : _GEN_2309; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2311 = 7'h6 == out_payload_rob_idx[6:0] ? rob_payload_6_flits_fired : _GEN_2310; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2312 = 7'h7 == out_payload_rob_idx[6:0] ? rob_payload_7_flits_fired : _GEN_2311; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2313 = 7'h8 == out_payload_rob_idx[6:0] ? rob_payload_8_flits_fired : _GEN_2312; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2314 = 7'h9 == out_payload_rob_idx[6:0] ? rob_payload_9_flits_fired : _GEN_2313; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2315 = 7'ha == out_payload_rob_idx[6:0] ? rob_payload_10_flits_fired : _GEN_2314; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2316 = 7'hb == out_payload_rob_idx[6:0] ? rob_payload_11_flits_fired : _GEN_2315; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2317 = 7'hc == out_payload_rob_idx[6:0] ? rob_payload_12_flits_fired : _GEN_2316; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2318 = 7'hd == out_payload_rob_idx[6:0] ? rob_payload_13_flits_fired : _GEN_2317; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2319 = 7'he == out_payload_rob_idx[6:0] ? rob_payload_14_flits_fired : _GEN_2318; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2320 = 7'hf == out_payload_rob_idx[6:0] ? rob_payload_15_flits_fired : _GEN_2319; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2321 = 7'h10 == out_payload_rob_idx[6:0] ? rob_payload_16_flits_fired : _GEN_2320; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2322 = 7'h11 == out_payload_rob_idx[6:0] ? rob_payload_17_flits_fired : _GEN_2321; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2323 = 7'h12 == out_payload_rob_idx[6:0] ? rob_payload_18_flits_fired : _GEN_2322; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2324 = 7'h13 == out_payload_rob_idx[6:0] ? rob_payload_19_flits_fired : _GEN_2323; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2325 = 7'h14 == out_payload_rob_idx[6:0] ? rob_payload_20_flits_fired : _GEN_2324; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2326 = 7'h15 == out_payload_rob_idx[6:0] ? rob_payload_21_flits_fired : _GEN_2325; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2327 = 7'h16 == out_payload_rob_idx[6:0] ? rob_payload_22_flits_fired : _GEN_2326; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2328 = 7'h17 == out_payload_rob_idx[6:0] ? rob_payload_23_flits_fired : _GEN_2327; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2329 = 7'h18 == out_payload_rob_idx[6:0] ? rob_payload_24_flits_fired : _GEN_2328; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2330 = 7'h19 == out_payload_rob_idx[6:0] ? rob_payload_25_flits_fired : _GEN_2329; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2331 = 7'h1a == out_payload_rob_idx[6:0] ? rob_payload_26_flits_fired : _GEN_2330; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2332 = 7'h1b == out_payload_rob_idx[6:0] ? rob_payload_27_flits_fired : _GEN_2331; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2333 = 7'h1c == out_payload_rob_idx[6:0] ? rob_payload_28_flits_fired : _GEN_2332; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2334 = 7'h1d == out_payload_rob_idx[6:0] ? rob_payload_29_flits_fired : _GEN_2333; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2335 = 7'h1e == out_payload_rob_idx[6:0] ? rob_payload_30_flits_fired : _GEN_2334; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2336 = 7'h1f == out_payload_rob_idx[6:0] ? rob_payload_31_flits_fired : _GEN_2335; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2337 = 7'h20 == out_payload_rob_idx[6:0] ? rob_payload_32_flits_fired : _GEN_2336; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2338 = 7'h21 == out_payload_rob_idx[6:0] ? rob_payload_33_flits_fired : _GEN_2337; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2339 = 7'h22 == out_payload_rob_idx[6:0] ? rob_payload_34_flits_fired : _GEN_2338; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2340 = 7'h23 == out_payload_rob_idx[6:0] ? rob_payload_35_flits_fired : _GEN_2339; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2341 = 7'h24 == out_payload_rob_idx[6:0] ? rob_payload_36_flits_fired : _GEN_2340; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2342 = 7'h25 == out_payload_rob_idx[6:0] ? rob_payload_37_flits_fired : _GEN_2341; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2343 = 7'h26 == out_payload_rob_idx[6:0] ? rob_payload_38_flits_fired : _GEN_2342; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2344 = 7'h27 == out_payload_rob_idx[6:0] ? rob_payload_39_flits_fired : _GEN_2343; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2345 = 7'h28 == out_payload_rob_idx[6:0] ? rob_payload_40_flits_fired : _GEN_2344; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2346 = 7'h29 == out_payload_rob_idx[6:0] ? rob_payload_41_flits_fired : _GEN_2345; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2347 = 7'h2a == out_payload_rob_idx[6:0] ? rob_payload_42_flits_fired : _GEN_2346; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2348 = 7'h2b == out_payload_rob_idx[6:0] ? rob_payload_43_flits_fired : _GEN_2347; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2349 = 7'h2c == out_payload_rob_idx[6:0] ? rob_payload_44_flits_fired : _GEN_2348; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2350 = 7'h2d == out_payload_rob_idx[6:0] ? rob_payload_45_flits_fired : _GEN_2349; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2351 = 7'h2e == out_payload_rob_idx[6:0] ? rob_payload_46_flits_fired : _GEN_2350; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2352 = 7'h2f == out_payload_rob_idx[6:0] ? rob_payload_47_flits_fired : _GEN_2351; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2353 = 7'h30 == out_payload_rob_idx[6:0] ? rob_payload_48_flits_fired : _GEN_2352; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2354 = 7'h31 == out_payload_rob_idx[6:0] ? rob_payload_49_flits_fired : _GEN_2353; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2355 = 7'h32 == out_payload_rob_idx[6:0] ? rob_payload_50_flits_fired : _GEN_2354; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2356 = 7'h33 == out_payload_rob_idx[6:0] ? rob_payload_51_flits_fired : _GEN_2355; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2357 = 7'h34 == out_payload_rob_idx[6:0] ? rob_payload_52_flits_fired : _GEN_2356; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2358 = 7'h35 == out_payload_rob_idx[6:0] ? rob_payload_53_flits_fired : _GEN_2357; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2359 = 7'h36 == out_payload_rob_idx[6:0] ? rob_payload_54_flits_fired : _GEN_2358; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2360 = 7'h37 == out_payload_rob_idx[6:0] ? rob_payload_55_flits_fired : _GEN_2359; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2361 = 7'h38 == out_payload_rob_idx[6:0] ? rob_payload_56_flits_fired : _GEN_2360; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2362 = 7'h39 == out_payload_rob_idx[6:0] ? rob_payload_57_flits_fired : _GEN_2361; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2363 = 7'h3a == out_payload_rob_idx[6:0] ? rob_payload_58_flits_fired : _GEN_2362; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2364 = 7'h3b == out_payload_rob_idx[6:0] ? rob_payload_59_flits_fired : _GEN_2363; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2365 = 7'h3c == out_payload_rob_idx[6:0] ? rob_payload_60_flits_fired : _GEN_2364; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2366 = 7'h3d == out_payload_rob_idx[6:0] ? rob_payload_61_flits_fired : _GEN_2365; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2367 = 7'h3e == out_payload_rob_idx[6:0] ? rob_payload_62_flits_fired : _GEN_2366; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2368 = 7'h3f == out_payload_rob_idx[6:0] ? rob_payload_63_flits_fired : _GEN_2367; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2369 = 7'h40 == out_payload_rob_idx[6:0] ? rob_payload_64_flits_fired : _GEN_2368; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2370 = 7'h41 == out_payload_rob_idx[6:0] ? rob_payload_65_flits_fired : _GEN_2369; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2371 = 7'h42 == out_payload_rob_idx[6:0] ? rob_payload_66_flits_fired : _GEN_2370; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2372 = 7'h43 == out_payload_rob_idx[6:0] ? rob_payload_67_flits_fired : _GEN_2371; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2373 = 7'h44 == out_payload_rob_idx[6:0] ? rob_payload_68_flits_fired : _GEN_2372; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2374 = 7'h45 == out_payload_rob_idx[6:0] ? rob_payload_69_flits_fired : _GEN_2373; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2375 = 7'h46 == out_payload_rob_idx[6:0] ? rob_payload_70_flits_fired : _GEN_2374; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2376 = 7'h47 == out_payload_rob_idx[6:0] ? rob_payload_71_flits_fired : _GEN_2375; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2377 = 7'h48 == out_payload_rob_idx[6:0] ? rob_payload_72_flits_fired : _GEN_2376; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2378 = 7'h49 == out_payload_rob_idx[6:0] ? rob_payload_73_flits_fired : _GEN_2377; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2379 = 7'h4a == out_payload_rob_idx[6:0] ? rob_payload_74_flits_fired : _GEN_2378; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2380 = 7'h4b == out_payload_rob_idx[6:0] ? rob_payload_75_flits_fired : _GEN_2379; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2381 = 7'h4c == out_payload_rob_idx[6:0] ? rob_payload_76_flits_fired : _GEN_2380; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2382 = 7'h4d == out_payload_rob_idx[6:0] ? rob_payload_77_flits_fired : _GEN_2381; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2383 = 7'h4e == out_payload_rob_idx[6:0] ? rob_payload_78_flits_fired : _GEN_2382; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2384 = 7'h4f == out_payload_rob_idx[6:0] ? rob_payload_79_flits_fired : _GEN_2383; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2385 = 7'h50 == out_payload_rob_idx[6:0] ? rob_payload_80_flits_fired : _GEN_2384; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2386 = 7'h51 == out_payload_rob_idx[6:0] ? rob_payload_81_flits_fired : _GEN_2385; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2387 = 7'h52 == out_payload_rob_idx[6:0] ? rob_payload_82_flits_fired : _GEN_2386; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2388 = 7'h53 == out_payload_rob_idx[6:0] ? rob_payload_83_flits_fired : _GEN_2387; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2389 = 7'h54 == out_payload_rob_idx[6:0] ? rob_payload_84_flits_fired : _GEN_2388; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2390 = 7'h55 == out_payload_rob_idx[6:0] ? rob_payload_85_flits_fired : _GEN_2389; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2391 = 7'h56 == out_payload_rob_idx[6:0] ? rob_payload_86_flits_fired : _GEN_2390; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2392 = 7'h57 == out_payload_rob_idx[6:0] ? rob_payload_87_flits_fired : _GEN_2391; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2393 = 7'h58 == out_payload_rob_idx[6:0] ? rob_payload_88_flits_fired : _GEN_2392; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2394 = 7'h59 == out_payload_rob_idx[6:0] ? rob_payload_89_flits_fired : _GEN_2393; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2395 = 7'h5a == out_payload_rob_idx[6:0] ? rob_payload_90_flits_fired : _GEN_2394; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2396 = 7'h5b == out_payload_rob_idx[6:0] ? rob_payload_91_flits_fired : _GEN_2395; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2397 = 7'h5c == out_payload_rob_idx[6:0] ? rob_payload_92_flits_fired : _GEN_2396; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2398 = 7'h5d == out_payload_rob_idx[6:0] ? rob_payload_93_flits_fired : _GEN_2397; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2399 = 7'h5e == out_payload_rob_idx[6:0] ? rob_payload_94_flits_fired : _GEN_2398; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2400 = 7'h5f == out_payload_rob_idx[6:0] ? rob_payload_95_flits_fired : _GEN_2399; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2401 = 7'h60 == out_payload_rob_idx[6:0] ? rob_payload_96_flits_fired : _GEN_2400; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2402 = 7'h61 == out_payload_rob_idx[6:0] ? rob_payload_97_flits_fired : _GEN_2401; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2403 = 7'h62 == out_payload_rob_idx[6:0] ? rob_payload_98_flits_fired : _GEN_2402; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2404 = 7'h63 == out_payload_rob_idx[6:0] ? rob_payload_99_flits_fired : _GEN_2403; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2405 = 7'h64 == out_payload_rob_idx[6:0] ? rob_payload_100_flits_fired : _GEN_2404; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2406 = 7'h65 == out_payload_rob_idx[6:0] ? rob_payload_101_flits_fired : _GEN_2405; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2407 = 7'h66 == out_payload_rob_idx[6:0] ? rob_payload_102_flits_fired : _GEN_2406; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2408 = 7'h67 == out_payload_rob_idx[6:0] ? rob_payload_103_flits_fired : _GEN_2407; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2409 = 7'h68 == out_payload_rob_idx[6:0] ? rob_payload_104_flits_fired : _GEN_2408; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2410 = 7'h69 == out_payload_rob_idx[6:0] ? rob_payload_105_flits_fired : _GEN_2409; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2411 = 7'h6a == out_payload_rob_idx[6:0] ? rob_payload_106_flits_fired : _GEN_2410; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2412 = 7'h6b == out_payload_rob_idx[6:0] ? rob_payload_107_flits_fired : _GEN_2411; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2413 = 7'h6c == out_payload_rob_idx[6:0] ? rob_payload_108_flits_fired : _GEN_2412; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2414 = 7'h6d == out_payload_rob_idx[6:0] ? rob_payload_109_flits_fired : _GEN_2413; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2415 = 7'h6e == out_payload_rob_idx[6:0] ? rob_payload_110_flits_fired : _GEN_2414; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2416 = 7'h6f == out_payload_rob_idx[6:0] ? rob_payload_111_flits_fired : _GEN_2415; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2417 = 7'h70 == out_payload_rob_idx[6:0] ? rob_payload_112_flits_fired : _GEN_2416; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2418 = 7'h71 == out_payload_rob_idx[6:0] ? rob_payload_113_flits_fired : _GEN_2417; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2419 = 7'h72 == out_payload_rob_idx[6:0] ? rob_payload_114_flits_fired : _GEN_2418; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2420 = 7'h73 == out_payload_rob_idx[6:0] ? rob_payload_115_flits_fired : _GEN_2419; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2421 = 7'h74 == out_payload_rob_idx[6:0] ? rob_payload_116_flits_fired : _GEN_2420; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2422 = 7'h75 == out_payload_rob_idx[6:0] ? rob_payload_117_flits_fired : _GEN_2421; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2423 = 7'h76 == out_payload_rob_idx[6:0] ? rob_payload_118_flits_fired : _GEN_2422; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2424 = 7'h77 == out_payload_rob_idx[6:0] ? rob_payload_119_flits_fired : _GEN_2423; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2425 = 7'h78 == out_payload_rob_idx[6:0] ? rob_payload_120_flits_fired : _GEN_2424; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2426 = 7'h79 == out_payload_rob_idx[6:0] ? rob_payload_121_flits_fired : _GEN_2425; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2427 = 7'h7a == out_payload_rob_idx[6:0] ? rob_payload_122_flits_fired : _GEN_2426; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2428 = 7'h7b == out_payload_rob_idx[6:0] ? rob_payload_123_flits_fired : _GEN_2427; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2429 = 7'h7c == out_payload_rob_idx[6:0] ? rob_payload_124_flits_fired : _GEN_2428; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2430 = 7'h7d == out_payload_rob_idx[6:0] ? rob_payload_125_flits_fired : _GEN_2429; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2431 = 7'h7e == out_payload_rob_idx[6:0] ? rob_payload_126_flits_fired : _GEN_2430; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_2432 = 7'h7f == out_payload_rob_idx[6:0] ? rob_payload_127_flits_fired : _GEN_2431; // @[TestHarness.scala 202:{35,35}]
  wire [63:0] _T_31 = {_GEN_2176,_GEN_2304,_GEN_2432}; // @[TestHarness.scala 202:35]
  wire [3:0] _GEN_2690 = 7'h1 == out_payload_rob_idx[6:0] ? rob_flits_returned_1 : rob_flits_returned_0; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2691 = 7'h2 == out_payload_rob_idx[6:0] ? rob_flits_returned_2 : _GEN_2690; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2692 = 7'h3 == out_payload_rob_idx[6:0] ? rob_flits_returned_3 : _GEN_2691; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2693 = 7'h4 == out_payload_rob_idx[6:0] ? rob_flits_returned_4 : _GEN_2692; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2694 = 7'h5 == out_payload_rob_idx[6:0] ? rob_flits_returned_5 : _GEN_2693; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2695 = 7'h6 == out_payload_rob_idx[6:0] ? rob_flits_returned_6 : _GEN_2694; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2696 = 7'h7 == out_payload_rob_idx[6:0] ? rob_flits_returned_7 : _GEN_2695; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2697 = 7'h8 == out_payload_rob_idx[6:0] ? rob_flits_returned_8 : _GEN_2696; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2698 = 7'h9 == out_payload_rob_idx[6:0] ? rob_flits_returned_9 : _GEN_2697; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2699 = 7'ha == out_payload_rob_idx[6:0] ? rob_flits_returned_10 : _GEN_2698; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2700 = 7'hb == out_payload_rob_idx[6:0] ? rob_flits_returned_11 : _GEN_2699; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2701 = 7'hc == out_payload_rob_idx[6:0] ? rob_flits_returned_12 : _GEN_2700; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2702 = 7'hd == out_payload_rob_idx[6:0] ? rob_flits_returned_13 : _GEN_2701; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2703 = 7'he == out_payload_rob_idx[6:0] ? rob_flits_returned_14 : _GEN_2702; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2704 = 7'hf == out_payload_rob_idx[6:0] ? rob_flits_returned_15 : _GEN_2703; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2705 = 7'h10 == out_payload_rob_idx[6:0] ? rob_flits_returned_16 : _GEN_2704; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2706 = 7'h11 == out_payload_rob_idx[6:0] ? rob_flits_returned_17 : _GEN_2705; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2707 = 7'h12 == out_payload_rob_idx[6:0] ? rob_flits_returned_18 : _GEN_2706; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2708 = 7'h13 == out_payload_rob_idx[6:0] ? rob_flits_returned_19 : _GEN_2707; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2709 = 7'h14 == out_payload_rob_idx[6:0] ? rob_flits_returned_20 : _GEN_2708; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2710 = 7'h15 == out_payload_rob_idx[6:0] ? rob_flits_returned_21 : _GEN_2709; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2711 = 7'h16 == out_payload_rob_idx[6:0] ? rob_flits_returned_22 : _GEN_2710; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2712 = 7'h17 == out_payload_rob_idx[6:0] ? rob_flits_returned_23 : _GEN_2711; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2713 = 7'h18 == out_payload_rob_idx[6:0] ? rob_flits_returned_24 : _GEN_2712; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2714 = 7'h19 == out_payload_rob_idx[6:0] ? rob_flits_returned_25 : _GEN_2713; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2715 = 7'h1a == out_payload_rob_idx[6:0] ? rob_flits_returned_26 : _GEN_2714; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2716 = 7'h1b == out_payload_rob_idx[6:0] ? rob_flits_returned_27 : _GEN_2715; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2717 = 7'h1c == out_payload_rob_idx[6:0] ? rob_flits_returned_28 : _GEN_2716; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2718 = 7'h1d == out_payload_rob_idx[6:0] ? rob_flits_returned_29 : _GEN_2717; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2719 = 7'h1e == out_payload_rob_idx[6:0] ? rob_flits_returned_30 : _GEN_2718; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2720 = 7'h1f == out_payload_rob_idx[6:0] ? rob_flits_returned_31 : _GEN_2719; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2721 = 7'h20 == out_payload_rob_idx[6:0] ? rob_flits_returned_32 : _GEN_2720; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2722 = 7'h21 == out_payload_rob_idx[6:0] ? rob_flits_returned_33 : _GEN_2721; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2723 = 7'h22 == out_payload_rob_idx[6:0] ? rob_flits_returned_34 : _GEN_2722; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2724 = 7'h23 == out_payload_rob_idx[6:0] ? rob_flits_returned_35 : _GEN_2723; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2725 = 7'h24 == out_payload_rob_idx[6:0] ? rob_flits_returned_36 : _GEN_2724; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2726 = 7'h25 == out_payload_rob_idx[6:0] ? rob_flits_returned_37 : _GEN_2725; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2727 = 7'h26 == out_payload_rob_idx[6:0] ? rob_flits_returned_38 : _GEN_2726; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2728 = 7'h27 == out_payload_rob_idx[6:0] ? rob_flits_returned_39 : _GEN_2727; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2729 = 7'h28 == out_payload_rob_idx[6:0] ? rob_flits_returned_40 : _GEN_2728; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2730 = 7'h29 == out_payload_rob_idx[6:0] ? rob_flits_returned_41 : _GEN_2729; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2731 = 7'h2a == out_payload_rob_idx[6:0] ? rob_flits_returned_42 : _GEN_2730; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2732 = 7'h2b == out_payload_rob_idx[6:0] ? rob_flits_returned_43 : _GEN_2731; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2733 = 7'h2c == out_payload_rob_idx[6:0] ? rob_flits_returned_44 : _GEN_2732; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2734 = 7'h2d == out_payload_rob_idx[6:0] ? rob_flits_returned_45 : _GEN_2733; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2735 = 7'h2e == out_payload_rob_idx[6:0] ? rob_flits_returned_46 : _GEN_2734; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2736 = 7'h2f == out_payload_rob_idx[6:0] ? rob_flits_returned_47 : _GEN_2735; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2737 = 7'h30 == out_payload_rob_idx[6:0] ? rob_flits_returned_48 : _GEN_2736; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2738 = 7'h31 == out_payload_rob_idx[6:0] ? rob_flits_returned_49 : _GEN_2737; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2739 = 7'h32 == out_payload_rob_idx[6:0] ? rob_flits_returned_50 : _GEN_2738; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2740 = 7'h33 == out_payload_rob_idx[6:0] ? rob_flits_returned_51 : _GEN_2739; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2741 = 7'h34 == out_payload_rob_idx[6:0] ? rob_flits_returned_52 : _GEN_2740; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2742 = 7'h35 == out_payload_rob_idx[6:0] ? rob_flits_returned_53 : _GEN_2741; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2743 = 7'h36 == out_payload_rob_idx[6:0] ? rob_flits_returned_54 : _GEN_2742; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2744 = 7'h37 == out_payload_rob_idx[6:0] ? rob_flits_returned_55 : _GEN_2743; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2745 = 7'h38 == out_payload_rob_idx[6:0] ? rob_flits_returned_56 : _GEN_2744; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2746 = 7'h39 == out_payload_rob_idx[6:0] ? rob_flits_returned_57 : _GEN_2745; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2747 = 7'h3a == out_payload_rob_idx[6:0] ? rob_flits_returned_58 : _GEN_2746; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2748 = 7'h3b == out_payload_rob_idx[6:0] ? rob_flits_returned_59 : _GEN_2747; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2749 = 7'h3c == out_payload_rob_idx[6:0] ? rob_flits_returned_60 : _GEN_2748; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2750 = 7'h3d == out_payload_rob_idx[6:0] ? rob_flits_returned_61 : _GEN_2749; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2751 = 7'h3e == out_payload_rob_idx[6:0] ? rob_flits_returned_62 : _GEN_2750; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2752 = 7'h3f == out_payload_rob_idx[6:0] ? rob_flits_returned_63 : _GEN_2751; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2753 = 7'h40 == out_payload_rob_idx[6:0] ? rob_flits_returned_64 : _GEN_2752; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2754 = 7'h41 == out_payload_rob_idx[6:0] ? rob_flits_returned_65 : _GEN_2753; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2755 = 7'h42 == out_payload_rob_idx[6:0] ? rob_flits_returned_66 : _GEN_2754; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2756 = 7'h43 == out_payload_rob_idx[6:0] ? rob_flits_returned_67 : _GEN_2755; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2757 = 7'h44 == out_payload_rob_idx[6:0] ? rob_flits_returned_68 : _GEN_2756; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2758 = 7'h45 == out_payload_rob_idx[6:0] ? rob_flits_returned_69 : _GEN_2757; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2759 = 7'h46 == out_payload_rob_idx[6:0] ? rob_flits_returned_70 : _GEN_2758; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2760 = 7'h47 == out_payload_rob_idx[6:0] ? rob_flits_returned_71 : _GEN_2759; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2761 = 7'h48 == out_payload_rob_idx[6:0] ? rob_flits_returned_72 : _GEN_2760; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2762 = 7'h49 == out_payload_rob_idx[6:0] ? rob_flits_returned_73 : _GEN_2761; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2763 = 7'h4a == out_payload_rob_idx[6:0] ? rob_flits_returned_74 : _GEN_2762; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2764 = 7'h4b == out_payload_rob_idx[6:0] ? rob_flits_returned_75 : _GEN_2763; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2765 = 7'h4c == out_payload_rob_idx[6:0] ? rob_flits_returned_76 : _GEN_2764; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2766 = 7'h4d == out_payload_rob_idx[6:0] ? rob_flits_returned_77 : _GEN_2765; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2767 = 7'h4e == out_payload_rob_idx[6:0] ? rob_flits_returned_78 : _GEN_2766; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2768 = 7'h4f == out_payload_rob_idx[6:0] ? rob_flits_returned_79 : _GEN_2767; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2769 = 7'h50 == out_payload_rob_idx[6:0] ? rob_flits_returned_80 : _GEN_2768; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2770 = 7'h51 == out_payload_rob_idx[6:0] ? rob_flits_returned_81 : _GEN_2769; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2771 = 7'h52 == out_payload_rob_idx[6:0] ? rob_flits_returned_82 : _GEN_2770; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2772 = 7'h53 == out_payload_rob_idx[6:0] ? rob_flits_returned_83 : _GEN_2771; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2773 = 7'h54 == out_payload_rob_idx[6:0] ? rob_flits_returned_84 : _GEN_2772; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2774 = 7'h55 == out_payload_rob_idx[6:0] ? rob_flits_returned_85 : _GEN_2773; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2775 = 7'h56 == out_payload_rob_idx[6:0] ? rob_flits_returned_86 : _GEN_2774; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2776 = 7'h57 == out_payload_rob_idx[6:0] ? rob_flits_returned_87 : _GEN_2775; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2777 = 7'h58 == out_payload_rob_idx[6:0] ? rob_flits_returned_88 : _GEN_2776; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2778 = 7'h59 == out_payload_rob_idx[6:0] ? rob_flits_returned_89 : _GEN_2777; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2779 = 7'h5a == out_payload_rob_idx[6:0] ? rob_flits_returned_90 : _GEN_2778; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2780 = 7'h5b == out_payload_rob_idx[6:0] ? rob_flits_returned_91 : _GEN_2779; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2781 = 7'h5c == out_payload_rob_idx[6:0] ? rob_flits_returned_92 : _GEN_2780; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2782 = 7'h5d == out_payload_rob_idx[6:0] ? rob_flits_returned_93 : _GEN_2781; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2783 = 7'h5e == out_payload_rob_idx[6:0] ? rob_flits_returned_94 : _GEN_2782; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2784 = 7'h5f == out_payload_rob_idx[6:0] ? rob_flits_returned_95 : _GEN_2783; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2785 = 7'h60 == out_payload_rob_idx[6:0] ? rob_flits_returned_96 : _GEN_2784; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2786 = 7'h61 == out_payload_rob_idx[6:0] ? rob_flits_returned_97 : _GEN_2785; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2787 = 7'h62 == out_payload_rob_idx[6:0] ? rob_flits_returned_98 : _GEN_2786; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2788 = 7'h63 == out_payload_rob_idx[6:0] ? rob_flits_returned_99 : _GEN_2787; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2789 = 7'h64 == out_payload_rob_idx[6:0] ? rob_flits_returned_100 : _GEN_2788; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2790 = 7'h65 == out_payload_rob_idx[6:0] ? rob_flits_returned_101 : _GEN_2789; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2791 = 7'h66 == out_payload_rob_idx[6:0] ? rob_flits_returned_102 : _GEN_2790; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2792 = 7'h67 == out_payload_rob_idx[6:0] ? rob_flits_returned_103 : _GEN_2791; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2793 = 7'h68 == out_payload_rob_idx[6:0] ? rob_flits_returned_104 : _GEN_2792; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2794 = 7'h69 == out_payload_rob_idx[6:0] ? rob_flits_returned_105 : _GEN_2793; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2795 = 7'h6a == out_payload_rob_idx[6:0] ? rob_flits_returned_106 : _GEN_2794; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2796 = 7'h6b == out_payload_rob_idx[6:0] ? rob_flits_returned_107 : _GEN_2795; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2797 = 7'h6c == out_payload_rob_idx[6:0] ? rob_flits_returned_108 : _GEN_2796; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2798 = 7'h6d == out_payload_rob_idx[6:0] ? rob_flits_returned_109 : _GEN_2797; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2799 = 7'h6e == out_payload_rob_idx[6:0] ? rob_flits_returned_110 : _GEN_2798; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2800 = 7'h6f == out_payload_rob_idx[6:0] ? rob_flits_returned_111 : _GEN_2799; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2801 = 7'h70 == out_payload_rob_idx[6:0] ? rob_flits_returned_112 : _GEN_2800; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2802 = 7'h71 == out_payload_rob_idx[6:0] ? rob_flits_returned_113 : _GEN_2801; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2803 = 7'h72 == out_payload_rob_idx[6:0] ? rob_flits_returned_114 : _GEN_2802; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2804 = 7'h73 == out_payload_rob_idx[6:0] ? rob_flits_returned_115 : _GEN_2803; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2805 = 7'h74 == out_payload_rob_idx[6:0] ? rob_flits_returned_116 : _GEN_2804; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2806 = 7'h75 == out_payload_rob_idx[6:0] ? rob_flits_returned_117 : _GEN_2805; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2807 = 7'h76 == out_payload_rob_idx[6:0] ? rob_flits_returned_118 : _GEN_2806; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2808 = 7'h77 == out_payload_rob_idx[6:0] ? rob_flits_returned_119 : _GEN_2807; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2809 = 7'h78 == out_payload_rob_idx[6:0] ? rob_flits_returned_120 : _GEN_2808; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2810 = 7'h79 == out_payload_rob_idx[6:0] ? rob_flits_returned_121 : _GEN_2809; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2811 = 7'h7a == out_payload_rob_idx[6:0] ? rob_flits_returned_122 : _GEN_2810; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2812 = 7'h7b == out_payload_rob_idx[6:0] ? rob_flits_returned_123 : _GEN_2811; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2813 = 7'h7c == out_payload_rob_idx[6:0] ? rob_flits_returned_124 : _GEN_2812; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2814 = 7'h7d == out_payload_rob_idx[6:0] ? rob_flits_returned_125 : _GEN_2813; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2815 = 7'h7e == out_payload_rob_idx[6:0] ? rob_flits_returned_126 : _GEN_2814; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2816 = 7'h7f == out_payload_rob_idx[6:0] ? rob_flits_returned_127 : _GEN_2815; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2818 = 7'h1 == out_payload_rob_idx[6:0] ? rob_n_flits_1 : rob_n_flits_0; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2819 = 7'h2 == out_payload_rob_idx[6:0] ? rob_n_flits_2 : _GEN_2818; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2820 = 7'h3 == out_payload_rob_idx[6:0] ? rob_n_flits_3 : _GEN_2819; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2821 = 7'h4 == out_payload_rob_idx[6:0] ? rob_n_flits_4 : _GEN_2820; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2822 = 7'h5 == out_payload_rob_idx[6:0] ? rob_n_flits_5 : _GEN_2821; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2823 = 7'h6 == out_payload_rob_idx[6:0] ? rob_n_flits_6 : _GEN_2822; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2824 = 7'h7 == out_payload_rob_idx[6:0] ? rob_n_flits_7 : _GEN_2823; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2825 = 7'h8 == out_payload_rob_idx[6:0] ? rob_n_flits_8 : _GEN_2824; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2826 = 7'h9 == out_payload_rob_idx[6:0] ? rob_n_flits_9 : _GEN_2825; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2827 = 7'ha == out_payload_rob_idx[6:0] ? rob_n_flits_10 : _GEN_2826; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2828 = 7'hb == out_payload_rob_idx[6:0] ? rob_n_flits_11 : _GEN_2827; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2829 = 7'hc == out_payload_rob_idx[6:0] ? rob_n_flits_12 : _GEN_2828; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2830 = 7'hd == out_payload_rob_idx[6:0] ? rob_n_flits_13 : _GEN_2829; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2831 = 7'he == out_payload_rob_idx[6:0] ? rob_n_flits_14 : _GEN_2830; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2832 = 7'hf == out_payload_rob_idx[6:0] ? rob_n_flits_15 : _GEN_2831; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2833 = 7'h10 == out_payload_rob_idx[6:0] ? rob_n_flits_16 : _GEN_2832; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2834 = 7'h11 == out_payload_rob_idx[6:0] ? rob_n_flits_17 : _GEN_2833; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2835 = 7'h12 == out_payload_rob_idx[6:0] ? rob_n_flits_18 : _GEN_2834; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2836 = 7'h13 == out_payload_rob_idx[6:0] ? rob_n_flits_19 : _GEN_2835; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2837 = 7'h14 == out_payload_rob_idx[6:0] ? rob_n_flits_20 : _GEN_2836; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2838 = 7'h15 == out_payload_rob_idx[6:0] ? rob_n_flits_21 : _GEN_2837; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2839 = 7'h16 == out_payload_rob_idx[6:0] ? rob_n_flits_22 : _GEN_2838; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2840 = 7'h17 == out_payload_rob_idx[6:0] ? rob_n_flits_23 : _GEN_2839; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2841 = 7'h18 == out_payload_rob_idx[6:0] ? rob_n_flits_24 : _GEN_2840; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2842 = 7'h19 == out_payload_rob_idx[6:0] ? rob_n_flits_25 : _GEN_2841; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2843 = 7'h1a == out_payload_rob_idx[6:0] ? rob_n_flits_26 : _GEN_2842; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2844 = 7'h1b == out_payload_rob_idx[6:0] ? rob_n_flits_27 : _GEN_2843; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2845 = 7'h1c == out_payload_rob_idx[6:0] ? rob_n_flits_28 : _GEN_2844; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2846 = 7'h1d == out_payload_rob_idx[6:0] ? rob_n_flits_29 : _GEN_2845; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2847 = 7'h1e == out_payload_rob_idx[6:0] ? rob_n_flits_30 : _GEN_2846; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2848 = 7'h1f == out_payload_rob_idx[6:0] ? rob_n_flits_31 : _GEN_2847; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2849 = 7'h20 == out_payload_rob_idx[6:0] ? rob_n_flits_32 : _GEN_2848; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2850 = 7'h21 == out_payload_rob_idx[6:0] ? rob_n_flits_33 : _GEN_2849; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2851 = 7'h22 == out_payload_rob_idx[6:0] ? rob_n_flits_34 : _GEN_2850; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2852 = 7'h23 == out_payload_rob_idx[6:0] ? rob_n_flits_35 : _GEN_2851; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2853 = 7'h24 == out_payload_rob_idx[6:0] ? rob_n_flits_36 : _GEN_2852; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2854 = 7'h25 == out_payload_rob_idx[6:0] ? rob_n_flits_37 : _GEN_2853; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2855 = 7'h26 == out_payload_rob_idx[6:0] ? rob_n_flits_38 : _GEN_2854; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2856 = 7'h27 == out_payload_rob_idx[6:0] ? rob_n_flits_39 : _GEN_2855; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2857 = 7'h28 == out_payload_rob_idx[6:0] ? rob_n_flits_40 : _GEN_2856; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2858 = 7'h29 == out_payload_rob_idx[6:0] ? rob_n_flits_41 : _GEN_2857; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2859 = 7'h2a == out_payload_rob_idx[6:0] ? rob_n_flits_42 : _GEN_2858; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2860 = 7'h2b == out_payload_rob_idx[6:0] ? rob_n_flits_43 : _GEN_2859; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2861 = 7'h2c == out_payload_rob_idx[6:0] ? rob_n_flits_44 : _GEN_2860; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2862 = 7'h2d == out_payload_rob_idx[6:0] ? rob_n_flits_45 : _GEN_2861; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2863 = 7'h2e == out_payload_rob_idx[6:0] ? rob_n_flits_46 : _GEN_2862; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2864 = 7'h2f == out_payload_rob_idx[6:0] ? rob_n_flits_47 : _GEN_2863; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2865 = 7'h30 == out_payload_rob_idx[6:0] ? rob_n_flits_48 : _GEN_2864; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2866 = 7'h31 == out_payload_rob_idx[6:0] ? rob_n_flits_49 : _GEN_2865; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2867 = 7'h32 == out_payload_rob_idx[6:0] ? rob_n_flits_50 : _GEN_2866; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2868 = 7'h33 == out_payload_rob_idx[6:0] ? rob_n_flits_51 : _GEN_2867; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2869 = 7'h34 == out_payload_rob_idx[6:0] ? rob_n_flits_52 : _GEN_2868; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2870 = 7'h35 == out_payload_rob_idx[6:0] ? rob_n_flits_53 : _GEN_2869; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2871 = 7'h36 == out_payload_rob_idx[6:0] ? rob_n_flits_54 : _GEN_2870; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2872 = 7'h37 == out_payload_rob_idx[6:0] ? rob_n_flits_55 : _GEN_2871; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2873 = 7'h38 == out_payload_rob_idx[6:0] ? rob_n_flits_56 : _GEN_2872; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2874 = 7'h39 == out_payload_rob_idx[6:0] ? rob_n_flits_57 : _GEN_2873; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2875 = 7'h3a == out_payload_rob_idx[6:0] ? rob_n_flits_58 : _GEN_2874; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2876 = 7'h3b == out_payload_rob_idx[6:0] ? rob_n_flits_59 : _GEN_2875; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2877 = 7'h3c == out_payload_rob_idx[6:0] ? rob_n_flits_60 : _GEN_2876; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2878 = 7'h3d == out_payload_rob_idx[6:0] ? rob_n_flits_61 : _GEN_2877; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2879 = 7'h3e == out_payload_rob_idx[6:0] ? rob_n_flits_62 : _GEN_2878; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2880 = 7'h3f == out_payload_rob_idx[6:0] ? rob_n_flits_63 : _GEN_2879; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2881 = 7'h40 == out_payload_rob_idx[6:0] ? rob_n_flits_64 : _GEN_2880; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2882 = 7'h41 == out_payload_rob_idx[6:0] ? rob_n_flits_65 : _GEN_2881; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2883 = 7'h42 == out_payload_rob_idx[6:0] ? rob_n_flits_66 : _GEN_2882; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2884 = 7'h43 == out_payload_rob_idx[6:0] ? rob_n_flits_67 : _GEN_2883; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2885 = 7'h44 == out_payload_rob_idx[6:0] ? rob_n_flits_68 : _GEN_2884; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2886 = 7'h45 == out_payload_rob_idx[6:0] ? rob_n_flits_69 : _GEN_2885; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2887 = 7'h46 == out_payload_rob_idx[6:0] ? rob_n_flits_70 : _GEN_2886; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2888 = 7'h47 == out_payload_rob_idx[6:0] ? rob_n_flits_71 : _GEN_2887; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2889 = 7'h48 == out_payload_rob_idx[6:0] ? rob_n_flits_72 : _GEN_2888; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2890 = 7'h49 == out_payload_rob_idx[6:0] ? rob_n_flits_73 : _GEN_2889; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2891 = 7'h4a == out_payload_rob_idx[6:0] ? rob_n_flits_74 : _GEN_2890; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2892 = 7'h4b == out_payload_rob_idx[6:0] ? rob_n_flits_75 : _GEN_2891; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2893 = 7'h4c == out_payload_rob_idx[6:0] ? rob_n_flits_76 : _GEN_2892; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2894 = 7'h4d == out_payload_rob_idx[6:0] ? rob_n_flits_77 : _GEN_2893; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2895 = 7'h4e == out_payload_rob_idx[6:0] ? rob_n_flits_78 : _GEN_2894; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2896 = 7'h4f == out_payload_rob_idx[6:0] ? rob_n_flits_79 : _GEN_2895; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2897 = 7'h50 == out_payload_rob_idx[6:0] ? rob_n_flits_80 : _GEN_2896; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2898 = 7'h51 == out_payload_rob_idx[6:0] ? rob_n_flits_81 : _GEN_2897; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2899 = 7'h52 == out_payload_rob_idx[6:0] ? rob_n_flits_82 : _GEN_2898; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2900 = 7'h53 == out_payload_rob_idx[6:0] ? rob_n_flits_83 : _GEN_2899; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2901 = 7'h54 == out_payload_rob_idx[6:0] ? rob_n_flits_84 : _GEN_2900; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2902 = 7'h55 == out_payload_rob_idx[6:0] ? rob_n_flits_85 : _GEN_2901; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2903 = 7'h56 == out_payload_rob_idx[6:0] ? rob_n_flits_86 : _GEN_2902; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2904 = 7'h57 == out_payload_rob_idx[6:0] ? rob_n_flits_87 : _GEN_2903; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2905 = 7'h58 == out_payload_rob_idx[6:0] ? rob_n_flits_88 : _GEN_2904; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2906 = 7'h59 == out_payload_rob_idx[6:0] ? rob_n_flits_89 : _GEN_2905; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2907 = 7'h5a == out_payload_rob_idx[6:0] ? rob_n_flits_90 : _GEN_2906; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2908 = 7'h5b == out_payload_rob_idx[6:0] ? rob_n_flits_91 : _GEN_2907; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2909 = 7'h5c == out_payload_rob_idx[6:0] ? rob_n_flits_92 : _GEN_2908; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2910 = 7'h5d == out_payload_rob_idx[6:0] ? rob_n_flits_93 : _GEN_2909; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2911 = 7'h5e == out_payload_rob_idx[6:0] ? rob_n_flits_94 : _GEN_2910; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2912 = 7'h5f == out_payload_rob_idx[6:0] ? rob_n_flits_95 : _GEN_2911; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2913 = 7'h60 == out_payload_rob_idx[6:0] ? rob_n_flits_96 : _GEN_2912; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2914 = 7'h61 == out_payload_rob_idx[6:0] ? rob_n_flits_97 : _GEN_2913; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2915 = 7'h62 == out_payload_rob_idx[6:0] ? rob_n_flits_98 : _GEN_2914; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2916 = 7'h63 == out_payload_rob_idx[6:0] ? rob_n_flits_99 : _GEN_2915; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2917 = 7'h64 == out_payload_rob_idx[6:0] ? rob_n_flits_100 : _GEN_2916; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2918 = 7'h65 == out_payload_rob_idx[6:0] ? rob_n_flits_101 : _GEN_2917; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2919 = 7'h66 == out_payload_rob_idx[6:0] ? rob_n_flits_102 : _GEN_2918; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2920 = 7'h67 == out_payload_rob_idx[6:0] ? rob_n_flits_103 : _GEN_2919; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2921 = 7'h68 == out_payload_rob_idx[6:0] ? rob_n_flits_104 : _GEN_2920; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2922 = 7'h69 == out_payload_rob_idx[6:0] ? rob_n_flits_105 : _GEN_2921; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2923 = 7'h6a == out_payload_rob_idx[6:0] ? rob_n_flits_106 : _GEN_2922; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2924 = 7'h6b == out_payload_rob_idx[6:0] ? rob_n_flits_107 : _GEN_2923; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2925 = 7'h6c == out_payload_rob_idx[6:0] ? rob_n_flits_108 : _GEN_2924; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2926 = 7'h6d == out_payload_rob_idx[6:0] ? rob_n_flits_109 : _GEN_2925; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2927 = 7'h6e == out_payload_rob_idx[6:0] ? rob_n_flits_110 : _GEN_2926; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2928 = 7'h6f == out_payload_rob_idx[6:0] ? rob_n_flits_111 : _GEN_2927; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2929 = 7'h70 == out_payload_rob_idx[6:0] ? rob_n_flits_112 : _GEN_2928; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2930 = 7'h71 == out_payload_rob_idx[6:0] ? rob_n_flits_113 : _GEN_2929; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2931 = 7'h72 == out_payload_rob_idx[6:0] ? rob_n_flits_114 : _GEN_2930; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2932 = 7'h73 == out_payload_rob_idx[6:0] ? rob_n_flits_115 : _GEN_2931; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2933 = 7'h74 == out_payload_rob_idx[6:0] ? rob_n_flits_116 : _GEN_2932; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2934 = 7'h75 == out_payload_rob_idx[6:0] ? rob_n_flits_117 : _GEN_2933; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2935 = 7'h76 == out_payload_rob_idx[6:0] ? rob_n_flits_118 : _GEN_2934; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2936 = 7'h77 == out_payload_rob_idx[6:0] ? rob_n_flits_119 : _GEN_2935; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2937 = 7'h78 == out_payload_rob_idx[6:0] ? rob_n_flits_120 : _GEN_2936; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2938 = 7'h79 == out_payload_rob_idx[6:0] ? rob_n_flits_121 : _GEN_2937; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2939 = 7'h7a == out_payload_rob_idx[6:0] ? rob_n_flits_122 : _GEN_2938; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2940 = 7'h7b == out_payload_rob_idx[6:0] ? rob_n_flits_123 : _GEN_2939; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2941 = 7'h7c == out_payload_rob_idx[6:0] ? rob_n_flits_124 : _GEN_2940; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2942 = 7'h7d == out_payload_rob_idx[6:0] ? rob_n_flits_125 : _GEN_2941; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2943 = 7'h7e == out_payload_rob_idx[6:0] ? rob_n_flits_126 : _GEN_2942; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_2944 = 7'h7f == out_payload_rob_idx[6:0] ? rob_n_flits_127 : _GEN_2943; // @[TestHarness.scala 205:{42,42}]
  wire [15:0] _GEN_385 = {{9'd0}, packet_rob_idx}; // @[TestHarness.scala 206:61]
  wire  _T_59 = io_from_noc_0_flit_bits_head & enable_print_latency; // @[TestHarness.scala 208:30]
  wire [3:0] _rob_flits_returned_T_2 = _GEN_2816 + 4'h1; // @[TestHarness.scala 213:66]
  wire [15:0] _rob_payload_flits_fired_T_2 = _GEN_2432 + 16'h1; // @[TestHarness.scala 214:76]
  wire  _GEN_3585 = io_from_noc_0_flit_bits_head | packet_valid; // @[TestHarness.scala 196:31 215:{31,46}]
  wire [15:0] _GEN_3586 = io_from_noc_0_flit_bits_head ? out_payload_rob_idx : {{9'd0}, packet_rob_idx}; // @[TestHarness.scala 197:29 215:{31,72}]
  wire [15:0] _GEN_3845 = _T_67 ? _GEN_3586 : {{9'd0}, packet_rob_idx}; // @[TestHarness.scala 199:26 197:29]
  wire [127:0] _rob_valids_T = rob_valids | rob_allocs; // @[TestHarness.scala 222:29]
  wire [65535:0] _rob_valids_T_1 = ~rob_frees; // @[TestHarness.scala 222:45]
  wire [65535:0] _GEN_386 = {{65408'd0}, _rob_valids_T}; // @[TestHarness.scala 222:43]
  wire [65535:0] _rob_valids_T_2 = _GEN_386 & _rob_valids_T_1; // @[TestHarness.scala 222:43]
  wire [31:0] _GEN_387 = {{31'd0}, _T_67}; // @[TestHarness.scala 224:18]
  wire [31:0] _flits_T_2 = flits + _GEN_387; // @[TestHarness.scala 224:18]
  wire  tx_fire_0 = igen_io_fire; // @[TestHarness.scala 169:21 186:18]
  wire [31:0] _GEN_388 = {{31'd0}, tx_fire_0}; // @[TestHarness.scala 225:14]
  wire [31:0] _txs_T_1 = txs + _GEN_388; // @[TestHarness.scala 225:14]
  wire [63:0] _T_72 = _rob_tscs_T_22 - rob_tscs_0; // @[TestHarness.scala 229:18]
  wire [63:0] _T_79 = _rob_tscs_T_22 - rob_tscs_1; // @[TestHarness.scala 229:18]
  wire [63:0] _T_86 = _rob_tscs_T_22 - rob_tscs_2; // @[TestHarness.scala 229:18]
  wire [63:0] _T_93 = _rob_tscs_T_22 - rob_tscs_3; // @[TestHarness.scala 229:18]
  wire [63:0] _T_100 = _rob_tscs_T_22 - rob_tscs_4; // @[TestHarness.scala 229:18]
  wire [63:0] _T_107 = _rob_tscs_T_22 - rob_tscs_5; // @[TestHarness.scala 229:18]
  wire [63:0] _T_114 = _rob_tscs_T_22 - rob_tscs_6; // @[TestHarness.scala 229:18]
  wire [63:0] _T_121 = _rob_tscs_T_22 - rob_tscs_7; // @[TestHarness.scala 229:18]
  wire [63:0] _T_128 = _rob_tscs_T_22 - rob_tscs_8; // @[TestHarness.scala 229:18]
  wire [63:0] _T_135 = _rob_tscs_T_22 - rob_tscs_9; // @[TestHarness.scala 229:18]
  wire [63:0] _T_142 = _rob_tscs_T_22 - rob_tscs_10; // @[TestHarness.scala 229:18]
  wire [63:0] _T_149 = _rob_tscs_T_22 - rob_tscs_11; // @[TestHarness.scala 229:18]
  wire [63:0] _T_156 = _rob_tscs_T_22 - rob_tscs_12; // @[TestHarness.scala 229:18]
  wire [63:0] _T_163 = _rob_tscs_T_22 - rob_tscs_13; // @[TestHarness.scala 229:18]
  wire [63:0] _T_170 = _rob_tscs_T_22 - rob_tscs_14; // @[TestHarness.scala 229:18]
  wire [63:0] _T_177 = _rob_tscs_T_22 - rob_tscs_15; // @[TestHarness.scala 229:18]
  wire [63:0] _T_184 = _rob_tscs_T_22 - rob_tscs_16; // @[TestHarness.scala 229:18]
  wire [63:0] _T_191 = _rob_tscs_T_22 - rob_tscs_17; // @[TestHarness.scala 229:18]
  wire [63:0] _T_198 = _rob_tscs_T_22 - rob_tscs_18; // @[TestHarness.scala 229:18]
  wire [63:0] _T_205 = _rob_tscs_T_22 - rob_tscs_19; // @[TestHarness.scala 229:18]
  wire [63:0] _T_212 = _rob_tscs_T_22 - rob_tscs_20; // @[TestHarness.scala 229:18]
  wire [63:0] _T_219 = _rob_tscs_T_22 - rob_tscs_21; // @[TestHarness.scala 229:18]
  wire [63:0] _T_226 = _rob_tscs_T_22 - rob_tscs_22; // @[TestHarness.scala 229:18]
  wire [63:0] _T_233 = _rob_tscs_T_22 - rob_tscs_23; // @[TestHarness.scala 229:18]
  wire [63:0] _T_240 = _rob_tscs_T_22 - rob_tscs_24; // @[TestHarness.scala 229:18]
  wire [63:0] _T_247 = _rob_tscs_T_22 - rob_tscs_25; // @[TestHarness.scala 229:18]
  wire [63:0] _T_254 = _rob_tscs_T_22 - rob_tscs_26; // @[TestHarness.scala 229:18]
  wire [63:0] _T_261 = _rob_tscs_T_22 - rob_tscs_27; // @[TestHarness.scala 229:18]
  wire [63:0] _T_268 = _rob_tscs_T_22 - rob_tscs_28; // @[TestHarness.scala 229:18]
  wire [63:0] _T_275 = _rob_tscs_T_22 - rob_tscs_29; // @[TestHarness.scala 229:18]
  wire [63:0] _T_282 = _rob_tscs_T_22 - rob_tscs_30; // @[TestHarness.scala 229:18]
  wire [63:0] _T_289 = _rob_tscs_T_22 - rob_tscs_31; // @[TestHarness.scala 229:18]
  wire [63:0] _T_296 = _rob_tscs_T_22 - rob_tscs_32; // @[TestHarness.scala 229:18]
  wire [63:0] _T_303 = _rob_tscs_T_22 - rob_tscs_33; // @[TestHarness.scala 229:18]
  wire [63:0] _T_310 = _rob_tscs_T_22 - rob_tscs_34; // @[TestHarness.scala 229:18]
  wire [63:0] _T_317 = _rob_tscs_T_22 - rob_tscs_35; // @[TestHarness.scala 229:18]
  wire [63:0] _T_324 = _rob_tscs_T_22 - rob_tscs_36; // @[TestHarness.scala 229:18]
  wire [63:0] _T_331 = _rob_tscs_T_22 - rob_tscs_37; // @[TestHarness.scala 229:18]
  wire [63:0] _T_338 = _rob_tscs_T_22 - rob_tscs_38; // @[TestHarness.scala 229:18]
  wire [63:0] _T_345 = _rob_tscs_T_22 - rob_tscs_39; // @[TestHarness.scala 229:18]
  wire [63:0] _T_352 = _rob_tscs_T_22 - rob_tscs_40; // @[TestHarness.scala 229:18]
  wire [63:0] _T_359 = _rob_tscs_T_22 - rob_tscs_41; // @[TestHarness.scala 229:18]
  wire [63:0] _T_366 = _rob_tscs_T_22 - rob_tscs_42; // @[TestHarness.scala 229:18]
  wire [63:0] _T_373 = _rob_tscs_T_22 - rob_tscs_43; // @[TestHarness.scala 229:18]
  wire [63:0] _T_380 = _rob_tscs_T_22 - rob_tscs_44; // @[TestHarness.scala 229:18]
  wire [63:0] _T_387 = _rob_tscs_T_22 - rob_tscs_45; // @[TestHarness.scala 229:18]
  wire [63:0] _T_394 = _rob_tscs_T_22 - rob_tscs_46; // @[TestHarness.scala 229:18]
  wire [63:0] _T_401 = _rob_tscs_T_22 - rob_tscs_47; // @[TestHarness.scala 229:18]
  wire [63:0] _T_408 = _rob_tscs_T_22 - rob_tscs_48; // @[TestHarness.scala 229:18]
  wire [63:0] _T_415 = _rob_tscs_T_22 - rob_tscs_49; // @[TestHarness.scala 229:18]
  wire [63:0] _T_422 = _rob_tscs_T_22 - rob_tscs_50; // @[TestHarness.scala 229:18]
  wire [63:0] _T_429 = _rob_tscs_T_22 - rob_tscs_51; // @[TestHarness.scala 229:18]
  wire [63:0] _T_436 = _rob_tscs_T_22 - rob_tscs_52; // @[TestHarness.scala 229:18]
  wire [63:0] _T_443 = _rob_tscs_T_22 - rob_tscs_53; // @[TestHarness.scala 229:18]
  wire [63:0] _T_450 = _rob_tscs_T_22 - rob_tscs_54; // @[TestHarness.scala 229:18]
  wire [63:0] _T_457 = _rob_tscs_T_22 - rob_tscs_55; // @[TestHarness.scala 229:18]
  wire [63:0] _T_464 = _rob_tscs_T_22 - rob_tscs_56; // @[TestHarness.scala 229:18]
  wire [63:0] _T_471 = _rob_tscs_T_22 - rob_tscs_57; // @[TestHarness.scala 229:18]
  wire [63:0] _T_478 = _rob_tscs_T_22 - rob_tscs_58; // @[TestHarness.scala 229:18]
  wire [63:0] _T_485 = _rob_tscs_T_22 - rob_tscs_59; // @[TestHarness.scala 229:18]
  wire [63:0] _T_492 = _rob_tscs_T_22 - rob_tscs_60; // @[TestHarness.scala 229:18]
  wire [63:0] _T_499 = _rob_tscs_T_22 - rob_tscs_61; // @[TestHarness.scala 229:18]
  wire [63:0] _T_506 = _rob_tscs_T_22 - rob_tscs_62; // @[TestHarness.scala 229:18]
  wire [63:0] _T_513 = _rob_tscs_T_22 - rob_tscs_63; // @[TestHarness.scala 229:18]
  wire [63:0] _T_520 = _rob_tscs_T_22 - rob_tscs_64; // @[TestHarness.scala 229:18]
  wire [63:0] _T_527 = _rob_tscs_T_22 - rob_tscs_65; // @[TestHarness.scala 229:18]
  wire [63:0] _T_534 = _rob_tscs_T_22 - rob_tscs_66; // @[TestHarness.scala 229:18]
  wire [63:0] _T_541 = _rob_tscs_T_22 - rob_tscs_67; // @[TestHarness.scala 229:18]
  wire [63:0] _T_548 = _rob_tscs_T_22 - rob_tscs_68; // @[TestHarness.scala 229:18]
  wire [63:0] _T_555 = _rob_tscs_T_22 - rob_tscs_69; // @[TestHarness.scala 229:18]
  wire [63:0] _T_562 = _rob_tscs_T_22 - rob_tscs_70; // @[TestHarness.scala 229:18]
  wire [63:0] _T_569 = _rob_tscs_T_22 - rob_tscs_71; // @[TestHarness.scala 229:18]
  wire [63:0] _T_576 = _rob_tscs_T_22 - rob_tscs_72; // @[TestHarness.scala 229:18]
  wire [63:0] _T_583 = _rob_tscs_T_22 - rob_tscs_73; // @[TestHarness.scala 229:18]
  wire [63:0] _T_590 = _rob_tscs_T_22 - rob_tscs_74; // @[TestHarness.scala 229:18]
  wire [63:0] _T_597 = _rob_tscs_T_22 - rob_tscs_75; // @[TestHarness.scala 229:18]
  wire [63:0] _T_604 = _rob_tscs_T_22 - rob_tscs_76; // @[TestHarness.scala 229:18]
  wire [63:0] _T_611 = _rob_tscs_T_22 - rob_tscs_77; // @[TestHarness.scala 229:18]
  wire [63:0] _T_618 = _rob_tscs_T_22 - rob_tscs_78; // @[TestHarness.scala 229:18]
  wire [63:0] _T_625 = _rob_tscs_T_22 - rob_tscs_79; // @[TestHarness.scala 229:18]
  wire [63:0] _T_632 = _rob_tscs_T_22 - rob_tscs_80; // @[TestHarness.scala 229:18]
  wire [63:0] _T_639 = _rob_tscs_T_22 - rob_tscs_81; // @[TestHarness.scala 229:18]
  wire [63:0] _T_646 = _rob_tscs_T_22 - rob_tscs_82; // @[TestHarness.scala 229:18]
  wire [63:0] _T_653 = _rob_tscs_T_22 - rob_tscs_83; // @[TestHarness.scala 229:18]
  wire [63:0] _T_660 = _rob_tscs_T_22 - rob_tscs_84; // @[TestHarness.scala 229:18]
  wire [63:0] _T_667 = _rob_tscs_T_22 - rob_tscs_85; // @[TestHarness.scala 229:18]
  wire [63:0] _T_674 = _rob_tscs_T_22 - rob_tscs_86; // @[TestHarness.scala 229:18]
  wire [63:0] _T_681 = _rob_tscs_T_22 - rob_tscs_87; // @[TestHarness.scala 229:18]
  wire [63:0] _T_688 = _rob_tscs_T_22 - rob_tscs_88; // @[TestHarness.scala 229:18]
  wire [63:0] _T_695 = _rob_tscs_T_22 - rob_tscs_89; // @[TestHarness.scala 229:18]
  wire [63:0] _T_702 = _rob_tscs_T_22 - rob_tscs_90; // @[TestHarness.scala 229:18]
  wire [63:0] _T_709 = _rob_tscs_T_22 - rob_tscs_91; // @[TestHarness.scala 229:18]
  wire [63:0] _T_716 = _rob_tscs_T_22 - rob_tscs_92; // @[TestHarness.scala 229:18]
  wire [63:0] _T_723 = _rob_tscs_T_22 - rob_tscs_93; // @[TestHarness.scala 229:18]
  wire [63:0] _T_730 = _rob_tscs_T_22 - rob_tscs_94; // @[TestHarness.scala 229:18]
  wire [63:0] _T_737 = _rob_tscs_T_22 - rob_tscs_95; // @[TestHarness.scala 229:18]
  wire [63:0] _T_744 = _rob_tscs_T_22 - rob_tscs_96; // @[TestHarness.scala 229:18]
  wire [63:0] _T_751 = _rob_tscs_T_22 - rob_tscs_97; // @[TestHarness.scala 229:18]
  wire [63:0] _T_758 = _rob_tscs_T_22 - rob_tscs_98; // @[TestHarness.scala 229:18]
  wire [63:0] _T_765 = _rob_tscs_T_22 - rob_tscs_99; // @[TestHarness.scala 229:18]
  wire [63:0] _T_772 = _rob_tscs_T_22 - rob_tscs_100; // @[TestHarness.scala 229:18]
  wire [63:0] _T_779 = _rob_tscs_T_22 - rob_tscs_101; // @[TestHarness.scala 229:18]
  wire [63:0] _T_786 = _rob_tscs_T_22 - rob_tscs_102; // @[TestHarness.scala 229:18]
  wire [63:0] _T_793 = _rob_tscs_T_22 - rob_tscs_103; // @[TestHarness.scala 229:18]
  wire [63:0] _T_800 = _rob_tscs_T_22 - rob_tscs_104; // @[TestHarness.scala 229:18]
  wire [63:0] _T_807 = _rob_tscs_T_22 - rob_tscs_105; // @[TestHarness.scala 229:18]
  wire [63:0] _T_814 = _rob_tscs_T_22 - rob_tscs_106; // @[TestHarness.scala 229:18]
  wire [63:0] _T_821 = _rob_tscs_T_22 - rob_tscs_107; // @[TestHarness.scala 229:18]
  wire [63:0] _T_828 = _rob_tscs_T_22 - rob_tscs_108; // @[TestHarness.scala 229:18]
  wire [63:0] _T_835 = _rob_tscs_T_22 - rob_tscs_109; // @[TestHarness.scala 229:18]
  wire [63:0] _T_842 = _rob_tscs_T_22 - rob_tscs_110; // @[TestHarness.scala 229:18]
  wire [63:0] _T_849 = _rob_tscs_T_22 - rob_tscs_111; // @[TestHarness.scala 229:18]
  wire [63:0] _T_856 = _rob_tscs_T_22 - rob_tscs_112; // @[TestHarness.scala 229:18]
  wire [63:0] _T_863 = _rob_tscs_T_22 - rob_tscs_113; // @[TestHarness.scala 229:18]
  wire [63:0] _T_870 = _rob_tscs_T_22 - rob_tscs_114; // @[TestHarness.scala 229:18]
  wire [63:0] _T_877 = _rob_tscs_T_22 - rob_tscs_115; // @[TestHarness.scala 229:18]
  wire [63:0] _T_884 = _rob_tscs_T_22 - rob_tscs_116; // @[TestHarness.scala 229:18]
  wire [63:0] _T_891 = _rob_tscs_T_22 - rob_tscs_117; // @[TestHarness.scala 229:18]
  wire [63:0] _T_898 = _rob_tscs_T_22 - rob_tscs_118; // @[TestHarness.scala 229:18]
  wire [63:0] _T_905 = _rob_tscs_T_22 - rob_tscs_119; // @[TestHarness.scala 229:18]
  wire [63:0] _T_912 = _rob_tscs_T_22 - rob_tscs_120; // @[TestHarness.scala 229:18]
  wire [63:0] _T_919 = _rob_tscs_T_22 - rob_tscs_121; // @[TestHarness.scala 229:18]
  wire [63:0] _T_926 = _rob_tscs_T_22 - rob_tscs_122; // @[TestHarness.scala 229:18]
  wire [63:0] _T_933 = _rob_tscs_T_22 - rob_tscs_123; // @[TestHarness.scala 229:18]
  wire [63:0] _T_940 = _rob_tscs_T_22 - rob_tscs_124; // @[TestHarness.scala 229:18]
  wire [63:0] _T_947 = _rob_tscs_T_22 - rob_tscs_125; // @[TestHarness.scala 229:18]
  wire [63:0] _T_954 = _rob_tscs_T_22 - rob_tscs_126; // @[TestHarness.scala 229:18]
  wire [63:0] _T_961 = _rob_tscs_T_22 - rob_tscs_127; // @[TestHarness.scala 229:18]
  wire [65535:0] _GEN_517 = reset ? 65536'h0 : _rob_valids_T_2; // @[TestHarness.scala 156:{27,27} 222:14]
  wire  _GEN_518 = _T_67 & _T_3; // @[TestHarness.scala 201:13]
  InputGen igen ( // @[TestHarness.scala 171:22]
    .clock(igen_clock),
    .reset(igen_reset),
    .io_out_ready(igen_io_out_ready),
    .io_out_valid(igen_io_out_valid),
    .io_out_bits_head(igen_io_out_bits_head),
    .io_out_bits_tail(igen_io_out_bits_tail),
    .io_out_bits_payload(igen_io_out_bits_payload),
    .io_rob_ready(igen_io_rob_ready),
    .io_rob_idx(igen_io_rob_idx),
    .io_tsc(igen_io_tsc),
    .io_fire(igen_io_fire),
    .io_n_flits(igen_io_n_flits)
  );
  Queue_8 io_to_noc_0_flit_q ( // @[Decoupled.scala 375:21]
    .clock(io_to_noc_0_flit_q_clock),
    .reset(io_to_noc_0_flit_q_reset),
    .io_enq_ready(io_to_noc_0_flit_q_io_enq_ready),
    .io_enq_valid(io_to_noc_0_flit_q_io_enq_valid),
    .io_enq_bits_head(io_to_noc_0_flit_q_io_enq_bits_head),
    .io_enq_bits_tail(io_to_noc_0_flit_q_io_enq_bits_tail),
    .io_enq_bits_payload(io_to_noc_0_flit_q_io_enq_bits_payload),
    .io_deq_ready(io_to_noc_0_flit_q_io_deq_ready),
    .io_deq_valid(io_to_noc_0_flit_q_io_deq_valid),
    .io_deq_bits_head(io_to_noc_0_flit_q_io_deq_bits_head),
    .io_deq_bits_tail(io_to_noc_0_flit_q_io_deq_bits_tail),
    .io_deq_bits_payload(io_to_noc_0_flit_q_io_deq_bits_payload),
    .io_deq_bits_egress_id(io_to_noc_0_flit_q_io_deq_bits_egress_id)
  );
  plusarg_reader #(.FORMAT("noctest_enable_print=%d"), .DEFAULT(0), .WIDTH(1)) plusarg_reader ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_out)
  );
  MaxPeriodFibonacciLFSR io_from_noc_0_flit_ready_prng ( // @[PRNG.scala 91:22]
    .clock(io_from_noc_0_flit_ready_prng_clock),
    .reset(io_from_noc_0_flit_ready_prng_reset),
    .io_out_0(io_from_noc_0_flit_ready_prng_io_out_0),
    .io_out_1(io_from_noc_0_flit_ready_prng_io_out_1),
    .io_out_2(io_from_noc_0_flit_ready_prng_io_out_2),
    .io_out_3(io_from_noc_0_flit_ready_prng_io_out_3),
    .io_out_4(io_from_noc_0_flit_ready_prng_io_out_4),
    .io_out_5(io_from_noc_0_flit_ready_prng_io_out_5),
    .io_out_6(io_from_noc_0_flit_ready_prng_io_out_6),
    .io_out_7(io_from_noc_0_flit_ready_prng_io_out_7),
    .io_out_8(io_from_noc_0_flit_ready_prng_io_out_8),
    .io_out_9(io_from_noc_0_flit_ready_prng_io_out_9),
    .io_out_10(io_from_noc_0_flit_ready_prng_io_out_10),
    .io_out_11(io_from_noc_0_flit_ready_prng_io_out_11),
    .io_out_12(io_from_noc_0_flit_ready_prng_io_out_12),
    .io_out_13(io_from_noc_0_flit_ready_prng_io_out_13),
    .io_out_14(io_from_noc_0_flit_ready_prng_io_out_14),
    .io_out_15(io_from_noc_0_flit_ready_prng_io_out_15),
    .io_out_16(io_from_noc_0_flit_ready_prng_io_out_16),
    .io_out_17(io_from_noc_0_flit_ready_prng_io_out_17),
    .io_out_18(io_from_noc_0_flit_ready_prng_io_out_18),
    .io_out_19(io_from_noc_0_flit_ready_prng_io_out_19)
  );
  assign io_to_noc_0_flit_valid = io_to_noc_0_flit_q_io_deq_valid; // @[TestHarness.scala 177:12]
  assign io_to_noc_0_flit_bits_head = io_to_noc_0_flit_q_io_deq_bits_head; // @[TestHarness.scala 177:12]
  assign io_to_noc_0_flit_bits_tail = io_to_noc_0_flit_q_io_deq_bits_tail; // @[TestHarness.scala 177:12]
  assign io_to_noc_0_flit_bits_payload = io_to_noc_0_flit_q_io_deq_bits_payload; // @[TestHarness.scala 177:12]
  assign io_to_noc_0_flit_bits_egress_id = io_to_noc_0_flit_q_io_deq_bits_egress_id; // @[TestHarness.scala 177:12]
  assign io_from_noc_0_flit_ready = 1'h1; // @[TestHarness.scala 193:30]
  assign io_success = io_success_REG; // @[TestHarness.scala 164:14]
  assign igen_clock = clock;
  assign igen_reset = reset;
  assign igen_io_out_ready = io_to_noc_0_flit_q_io_enq_ready; // @[Decoupled.scala 379:17]
  assign igen_io_rob_ready = _igen_io_rob_ready_T_2 & txs < 32'hc350; // @[TestHarness.scala 175:19]
  assign igen_io_rob_idx = _T_5[0] ? 7'h0 : _sels_0_T_253; // @[Mux.scala 47:70]
  assign igen_io_tsc = tsc; // @[TestHarness.scala 176:17]
  assign io_to_noc_0_flit_q_clock = clock;
  assign io_to_noc_0_flit_q_reset = reset;
  assign io_to_noc_0_flit_q_io_enq_valid = igen_io_out_valid; // @[Decoupled.scala 377:22]
  assign io_to_noc_0_flit_q_io_enq_bits_head = igen_io_out_bits_head; // @[Decoupled.scala 378:21]
  assign io_to_noc_0_flit_q_io_enq_bits_tail = igen_io_out_bits_tail; // @[Decoupled.scala 378:21]
  assign io_to_noc_0_flit_q_io_enq_bits_payload = igen_io_out_bits_payload; // @[Decoupled.scala 378:21]
  assign io_to_noc_0_flit_q_io_deq_ready = io_to_noc_0_flit_ready; // @[TestHarness.scala 177:12]
  assign io_from_noc_0_flit_ready_prng_clock = clock;
  assign io_from_noc_0_flit_ready_prng_reset = reset;
  always @(posedge clock) begin
    if (reset) begin // @[TestHarness.scala 136:20]
      txs <= 32'h0; // @[TestHarness.scala 136:20]
    end else begin
      txs <= _txs_T_1; // @[TestHarness.scala 225:7]
    end
    if (reset) begin // @[TestHarness.scala 137:22]
      flits <= 32'h0; // @[TestHarness.scala 137:22]
    end else begin
      flits <= _flits_T_2; // @[TestHarness.scala 224:9]
    end
    if (reset) begin // @[TestHarness.scala 141:20]
      tsc <= 32'h0; // @[TestHarness.scala 141:20]
    end else begin
      tsc <= _tsc_T_1; // @[TestHarness.scala 142:7]
    end
    if (reset) begin // @[TestHarness.scala 144:29]
      idle_counter <= 11'h0; // @[TestHarness.scala 144:29]
    end else if (idle) begin // @[TestHarness.scala 146:15]
      idle_counter <= _idle_counter_T_1; // @[TestHarness.scala 146:30]
    end else begin
      idle_counter <= 11'h0; // @[TestHarness.scala 147:31]
    end
    rob_valids <= _GEN_517[127:0]; // @[TestHarness.scala 156:{27,27} 222:14]
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h0 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_0_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h0 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_0_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h0 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_0_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_0_flits_fired <= _GEN_1281;
      end
    end else begin
      rob_payload_0_flits_fired <= _GEN_1281;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_1_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_1_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h1 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_1_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_1_flits_fired <= _GEN_1282;
      end
    end else begin
      rob_payload_1_flits_fired <= _GEN_1282;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_2_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_2_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h2 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_2_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_2_flits_fired <= _GEN_1283;
      end
    end else begin
      rob_payload_2_flits_fired <= _GEN_1283;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_3_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_3_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h3 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_3_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_3_flits_fired <= _GEN_1284;
      end
    end else begin
      rob_payload_3_flits_fired <= _GEN_1284;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_4_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_4_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h4 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_4_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_4_flits_fired <= _GEN_1285;
      end
    end else begin
      rob_payload_4_flits_fired <= _GEN_1285;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_5_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_5_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h5 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_5_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_5_flits_fired <= _GEN_1286;
      end
    end else begin
      rob_payload_5_flits_fired <= _GEN_1286;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_6_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_6_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h6 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_6_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_6_flits_fired <= _GEN_1287;
      end
    end else begin
      rob_payload_6_flits_fired <= _GEN_1287;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_7_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_7_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h7 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_7_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_7_flits_fired <= _GEN_1288;
      end
    end else begin
      rob_payload_7_flits_fired <= _GEN_1288;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h8 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_8_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h8 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_8_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h8 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_8_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_8_flits_fired <= _GEN_1289;
      end
    end else begin
      rob_payload_8_flits_fired <= _GEN_1289;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h9 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_9_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h9 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_9_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h9 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_9_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_9_flits_fired <= _GEN_1290;
      end
    end else begin
      rob_payload_9_flits_fired <= _GEN_1290;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'ha == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_10_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'ha == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_10_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'ha == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_10_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_10_flits_fired <= _GEN_1291;
      end
    end else begin
      rob_payload_10_flits_fired <= _GEN_1291;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hb == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_11_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hb == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_11_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'hb == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_11_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_11_flits_fired <= _GEN_1292;
      end
    end else begin
      rob_payload_11_flits_fired <= _GEN_1292;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hc == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_12_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hc == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_12_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'hc == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_12_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_12_flits_fired <= _GEN_1293;
      end
    end else begin
      rob_payload_12_flits_fired <= _GEN_1293;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hd == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_13_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hd == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_13_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'hd == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_13_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_13_flits_fired <= _GEN_1294;
      end
    end else begin
      rob_payload_13_flits_fired <= _GEN_1294;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'he == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_14_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'he == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_14_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'he == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_14_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_14_flits_fired <= _GEN_1295;
      end
    end else begin
      rob_payload_14_flits_fired <= _GEN_1295;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hf == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_15_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hf == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_15_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'hf == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_15_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_15_flits_fired <= _GEN_1296;
      end
    end else begin
      rob_payload_15_flits_fired <= _GEN_1296;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h10 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_16_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h10 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_16_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h10 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_16_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_16_flits_fired <= _GEN_1297;
      end
    end else begin
      rob_payload_16_flits_fired <= _GEN_1297;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h11 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_17_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h11 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_17_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h11 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_17_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_17_flits_fired <= _GEN_1298;
      end
    end else begin
      rob_payload_17_flits_fired <= _GEN_1298;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h12 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_18_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h12 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_18_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h12 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_18_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_18_flits_fired <= _GEN_1299;
      end
    end else begin
      rob_payload_18_flits_fired <= _GEN_1299;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h13 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_19_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h13 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_19_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h13 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_19_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_19_flits_fired <= _GEN_1300;
      end
    end else begin
      rob_payload_19_flits_fired <= _GEN_1300;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h14 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_20_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h14 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_20_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h14 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_20_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_20_flits_fired <= _GEN_1301;
      end
    end else begin
      rob_payload_20_flits_fired <= _GEN_1301;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h15 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_21_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h15 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_21_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h15 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_21_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_21_flits_fired <= _GEN_1302;
      end
    end else begin
      rob_payload_21_flits_fired <= _GEN_1302;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h16 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_22_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h16 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_22_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h16 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_22_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_22_flits_fired <= _GEN_1303;
      end
    end else begin
      rob_payload_22_flits_fired <= _GEN_1303;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h17 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_23_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h17 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_23_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h17 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_23_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_23_flits_fired <= _GEN_1304;
      end
    end else begin
      rob_payload_23_flits_fired <= _GEN_1304;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h18 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_24_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h18 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_24_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h18 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_24_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_24_flits_fired <= _GEN_1305;
      end
    end else begin
      rob_payload_24_flits_fired <= _GEN_1305;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h19 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_25_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h19 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_25_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h19 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_25_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_25_flits_fired <= _GEN_1306;
      end
    end else begin
      rob_payload_25_flits_fired <= _GEN_1306;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1a == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_26_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1a == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_26_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h1a == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_26_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_26_flits_fired <= _GEN_1307;
      end
    end else begin
      rob_payload_26_flits_fired <= _GEN_1307;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1b == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_27_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1b == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_27_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h1b == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_27_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_27_flits_fired <= _GEN_1308;
      end
    end else begin
      rob_payload_27_flits_fired <= _GEN_1308;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1c == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_28_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1c == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_28_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h1c == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_28_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_28_flits_fired <= _GEN_1309;
      end
    end else begin
      rob_payload_28_flits_fired <= _GEN_1309;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1d == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_29_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1d == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_29_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h1d == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_29_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_29_flits_fired <= _GEN_1310;
      end
    end else begin
      rob_payload_29_flits_fired <= _GEN_1310;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1e == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_30_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1e == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_30_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h1e == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_30_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_30_flits_fired <= _GEN_1311;
      end
    end else begin
      rob_payload_30_flits_fired <= _GEN_1311;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1f == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_31_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1f == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_31_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h1f == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_31_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_31_flits_fired <= _GEN_1312;
      end
    end else begin
      rob_payload_31_flits_fired <= _GEN_1312;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h20 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_32_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h20 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_32_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h20 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_32_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_32_flits_fired <= _GEN_1313;
      end
    end else begin
      rob_payload_32_flits_fired <= _GEN_1313;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h21 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_33_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h21 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_33_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h21 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_33_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_33_flits_fired <= _GEN_1314;
      end
    end else begin
      rob_payload_33_flits_fired <= _GEN_1314;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h22 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_34_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h22 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_34_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h22 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_34_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_34_flits_fired <= _GEN_1315;
      end
    end else begin
      rob_payload_34_flits_fired <= _GEN_1315;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h23 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_35_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h23 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_35_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h23 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_35_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_35_flits_fired <= _GEN_1316;
      end
    end else begin
      rob_payload_35_flits_fired <= _GEN_1316;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h24 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_36_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h24 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_36_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h24 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_36_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_36_flits_fired <= _GEN_1317;
      end
    end else begin
      rob_payload_36_flits_fired <= _GEN_1317;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h25 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_37_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h25 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_37_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h25 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_37_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_37_flits_fired <= _GEN_1318;
      end
    end else begin
      rob_payload_37_flits_fired <= _GEN_1318;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h26 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_38_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h26 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_38_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h26 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_38_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_38_flits_fired <= _GEN_1319;
      end
    end else begin
      rob_payload_38_flits_fired <= _GEN_1319;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h27 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_39_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h27 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_39_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h27 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_39_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_39_flits_fired <= _GEN_1320;
      end
    end else begin
      rob_payload_39_flits_fired <= _GEN_1320;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h28 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_40_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h28 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_40_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h28 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_40_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_40_flits_fired <= _GEN_1321;
      end
    end else begin
      rob_payload_40_flits_fired <= _GEN_1321;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h29 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_41_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h29 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_41_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h29 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_41_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_41_flits_fired <= _GEN_1322;
      end
    end else begin
      rob_payload_41_flits_fired <= _GEN_1322;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2a == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_42_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2a == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_42_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h2a == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_42_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_42_flits_fired <= _GEN_1323;
      end
    end else begin
      rob_payload_42_flits_fired <= _GEN_1323;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2b == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_43_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2b == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_43_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h2b == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_43_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_43_flits_fired <= _GEN_1324;
      end
    end else begin
      rob_payload_43_flits_fired <= _GEN_1324;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2c == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_44_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2c == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_44_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h2c == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_44_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_44_flits_fired <= _GEN_1325;
      end
    end else begin
      rob_payload_44_flits_fired <= _GEN_1325;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2d == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_45_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2d == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_45_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h2d == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_45_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_45_flits_fired <= _GEN_1326;
      end
    end else begin
      rob_payload_45_flits_fired <= _GEN_1326;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2e == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_46_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2e == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_46_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h2e == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_46_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_46_flits_fired <= _GEN_1327;
      end
    end else begin
      rob_payload_46_flits_fired <= _GEN_1327;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2f == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_47_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2f == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_47_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h2f == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_47_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_47_flits_fired <= _GEN_1328;
      end
    end else begin
      rob_payload_47_flits_fired <= _GEN_1328;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h30 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_48_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h30 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_48_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h30 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_48_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_48_flits_fired <= _GEN_1329;
      end
    end else begin
      rob_payload_48_flits_fired <= _GEN_1329;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h31 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_49_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h31 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_49_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h31 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_49_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_49_flits_fired <= _GEN_1330;
      end
    end else begin
      rob_payload_49_flits_fired <= _GEN_1330;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h32 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_50_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h32 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_50_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h32 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_50_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_50_flits_fired <= _GEN_1331;
      end
    end else begin
      rob_payload_50_flits_fired <= _GEN_1331;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h33 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_51_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h33 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_51_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h33 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_51_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_51_flits_fired <= _GEN_1332;
      end
    end else begin
      rob_payload_51_flits_fired <= _GEN_1332;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h34 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_52_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h34 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_52_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h34 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_52_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_52_flits_fired <= _GEN_1333;
      end
    end else begin
      rob_payload_52_flits_fired <= _GEN_1333;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h35 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_53_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h35 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_53_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h35 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_53_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_53_flits_fired <= _GEN_1334;
      end
    end else begin
      rob_payload_53_flits_fired <= _GEN_1334;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h36 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_54_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h36 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_54_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h36 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_54_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_54_flits_fired <= _GEN_1335;
      end
    end else begin
      rob_payload_54_flits_fired <= _GEN_1335;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h37 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_55_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h37 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_55_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h37 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_55_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_55_flits_fired <= _GEN_1336;
      end
    end else begin
      rob_payload_55_flits_fired <= _GEN_1336;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h38 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_56_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h38 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_56_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h38 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_56_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_56_flits_fired <= _GEN_1337;
      end
    end else begin
      rob_payload_56_flits_fired <= _GEN_1337;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h39 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_57_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h39 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_57_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h39 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_57_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_57_flits_fired <= _GEN_1338;
      end
    end else begin
      rob_payload_57_flits_fired <= _GEN_1338;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3a == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_58_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3a == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_58_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h3a == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_58_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_58_flits_fired <= _GEN_1339;
      end
    end else begin
      rob_payload_58_flits_fired <= _GEN_1339;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3b == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_59_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3b == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_59_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h3b == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_59_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_59_flits_fired <= _GEN_1340;
      end
    end else begin
      rob_payload_59_flits_fired <= _GEN_1340;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3c == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_60_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3c == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_60_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h3c == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_60_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_60_flits_fired <= _GEN_1341;
      end
    end else begin
      rob_payload_60_flits_fired <= _GEN_1341;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3d == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_61_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3d == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_61_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h3d == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_61_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_61_flits_fired <= _GEN_1342;
      end
    end else begin
      rob_payload_61_flits_fired <= _GEN_1342;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3e == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_62_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3e == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_62_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h3e == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_62_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_62_flits_fired <= _GEN_1343;
      end
    end else begin
      rob_payload_62_flits_fired <= _GEN_1343;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3f == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_63_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3f == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_63_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h3f == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_63_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_63_flits_fired <= _GEN_1344;
      end
    end else begin
      rob_payload_63_flits_fired <= _GEN_1344;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h40 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_64_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h40 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_64_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h40 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_64_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_64_flits_fired <= _GEN_1345;
      end
    end else begin
      rob_payload_64_flits_fired <= _GEN_1345;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h41 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_65_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h41 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_65_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h41 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_65_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_65_flits_fired <= _GEN_1346;
      end
    end else begin
      rob_payload_65_flits_fired <= _GEN_1346;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h42 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_66_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h42 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_66_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h42 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_66_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_66_flits_fired <= _GEN_1347;
      end
    end else begin
      rob_payload_66_flits_fired <= _GEN_1347;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h43 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_67_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h43 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_67_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h43 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_67_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_67_flits_fired <= _GEN_1348;
      end
    end else begin
      rob_payload_67_flits_fired <= _GEN_1348;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h44 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_68_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h44 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_68_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h44 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_68_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_68_flits_fired <= _GEN_1349;
      end
    end else begin
      rob_payload_68_flits_fired <= _GEN_1349;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h45 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_69_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h45 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_69_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h45 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_69_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_69_flits_fired <= _GEN_1350;
      end
    end else begin
      rob_payload_69_flits_fired <= _GEN_1350;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h46 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_70_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h46 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_70_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h46 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_70_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_70_flits_fired <= _GEN_1351;
      end
    end else begin
      rob_payload_70_flits_fired <= _GEN_1351;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h47 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_71_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h47 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_71_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h47 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_71_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_71_flits_fired <= _GEN_1352;
      end
    end else begin
      rob_payload_71_flits_fired <= _GEN_1352;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h48 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_72_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h48 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_72_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h48 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_72_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_72_flits_fired <= _GEN_1353;
      end
    end else begin
      rob_payload_72_flits_fired <= _GEN_1353;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h49 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_73_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h49 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_73_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h49 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_73_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_73_flits_fired <= _GEN_1354;
      end
    end else begin
      rob_payload_73_flits_fired <= _GEN_1354;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4a == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_74_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4a == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_74_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h4a == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_74_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_74_flits_fired <= _GEN_1355;
      end
    end else begin
      rob_payload_74_flits_fired <= _GEN_1355;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4b == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_75_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4b == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_75_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h4b == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_75_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_75_flits_fired <= _GEN_1356;
      end
    end else begin
      rob_payload_75_flits_fired <= _GEN_1356;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4c == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_76_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4c == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_76_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h4c == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_76_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_76_flits_fired <= _GEN_1357;
      end
    end else begin
      rob_payload_76_flits_fired <= _GEN_1357;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4d == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_77_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4d == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_77_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h4d == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_77_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_77_flits_fired <= _GEN_1358;
      end
    end else begin
      rob_payload_77_flits_fired <= _GEN_1358;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4e == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_78_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4e == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_78_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h4e == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_78_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_78_flits_fired <= _GEN_1359;
      end
    end else begin
      rob_payload_78_flits_fired <= _GEN_1359;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4f == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_79_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4f == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_79_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h4f == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_79_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_79_flits_fired <= _GEN_1360;
      end
    end else begin
      rob_payload_79_flits_fired <= _GEN_1360;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h50 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_80_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h50 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_80_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h50 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_80_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_80_flits_fired <= _GEN_1361;
      end
    end else begin
      rob_payload_80_flits_fired <= _GEN_1361;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h51 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_81_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h51 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_81_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h51 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_81_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_81_flits_fired <= _GEN_1362;
      end
    end else begin
      rob_payload_81_flits_fired <= _GEN_1362;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h52 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_82_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h52 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_82_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h52 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_82_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_82_flits_fired <= _GEN_1363;
      end
    end else begin
      rob_payload_82_flits_fired <= _GEN_1363;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h53 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_83_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h53 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_83_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h53 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_83_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_83_flits_fired <= _GEN_1364;
      end
    end else begin
      rob_payload_83_flits_fired <= _GEN_1364;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h54 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_84_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h54 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_84_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h54 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_84_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_84_flits_fired <= _GEN_1365;
      end
    end else begin
      rob_payload_84_flits_fired <= _GEN_1365;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h55 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_85_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h55 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_85_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h55 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_85_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_85_flits_fired <= _GEN_1366;
      end
    end else begin
      rob_payload_85_flits_fired <= _GEN_1366;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h56 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_86_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h56 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_86_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h56 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_86_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_86_flits_fired <= _GEN_1367;
      end
    end else begin
      rob_payload_86_flits_fired <= _GEN_1367;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h57 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_87_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h57 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_87_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h57 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_87_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_87_flits_fired <= _GEN_1368;
      end
    end else begin
      rob_payload_87_flits_fired <= _GEN_1368;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h58 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_88_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h58 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_88_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h58 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_88_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_88_flits_fired <= _GEN_1369;
      end
    end else begin
      rob_payload_88_flits_fired <= _GEN_1369;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h59 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_89_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h59 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_89_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h59 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_89_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_89_flits_fired <= _GEN_1370;
      end
    end else begin
      rob_payload_89_flits_fired <= _GEN_1370;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5a == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_90_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5a == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_90_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h5a == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_90_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_90_flits_fired <= _GEN_1371;
      end
    end else begin
      rob_payload_90_flits_fired <= _GEN_1371;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5b == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_91_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5b == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_91_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h5b == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_91_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_91_flits_fired <= _GEN_1372;
      end
    end else begin
      rob_payload_91_flits_fired <= _GEN_1372;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5c == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_92_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5c == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_92_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h5c == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_92_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_92_flits_fired <= _GEN_1373;
      end
    end else begin
      rob_payload_92_flits_fired <= _GEN_1373;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5d == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_93_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5d == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_93_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h5d == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_93_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_93_flits_fired <= _GEN_1374;
      end
    end else begin
      rob_payload_93_flits_fired <= _GEN_1374;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5e == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_94_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5e == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_94_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h5e == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_94_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_94_flits_fired <= _GEN_1375;
      end
    end else begin
      rob_payload_94_flits_fired <= _GEN_1375;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5f == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_95_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5f == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_95_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h5f == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_95_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_95_flits_fired <= _GEN_1376;
      end
    end else begin
      rob_payload_95_flits_fired <= _GEN_1376;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h60 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_96_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h60 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_96_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h60 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_96_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_96_flits_fired <= _GEN_1377;
      end
    end else begin
      rob_payload_96_flits_fired <= _GEN_1377;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h61 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_97_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h61 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_97_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h61 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_97_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_97_flits_fired <= _GEN_1378;
      end
    end else begin
      rob_payload_97_flits_fired <= _GEN_1378;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h62 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_98_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h62 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_98_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h62 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_98_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_98_flits_fired <= _GEN_1379;
      end
    end else begin
      rob_payload_98_flits_fired <= _GEN_1379;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h63 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_99_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h63 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_99_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h63 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_99_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_99_flits_fired <= _GEN_1380;
      end
    end else begin
      rob_payload_99_flits_fired <= _GEN_1380;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h64 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_100_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h64 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_100_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h64 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_100_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_100_flits_fired <= _GEN_1381;
      end
    end else begin
      rob_payload_100_flits_fired <= _GEN_1381;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h65 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_101_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h65 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_101_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h65 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_101_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_101_flits_fired <= _GEN_1382;
      end
    end else begin
      rob_payload_101_flits_fired <= _GEN_1382;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h66 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_102_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h66 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_102_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h66 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_102_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_102_flits_fired <= _GEN_1383;
      end
    end else begin
      rob_payload_102_flits_fired <= _GEN_1383;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h67 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_103_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h67 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_103_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h67 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_103_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_103_flits_fired <= _GEN_1384;
      end
    end else begin
      rob_payload_103_flits_fired <= _GEN_1384;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h68 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_104_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h68 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_104_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h68 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_104_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_104_flits_fired <= _GEN_1385;
      end
    end else begin
      rob_payload_104_flits_fired <= _GEN_1385;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h69 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_105_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h69 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_105_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h69 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_105_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_105_flits_fired <= _GEN_1386;
      end
    end else begin
      rob_payload_105_flits_fired <= _GEN_1386;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6a == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_106_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6a == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_106_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h6a == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_106_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_106_flits_fired <= _GEN_1387;
      end
    end else begin
      rob_payload_106_flits_fired <= _GEN_1387;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6b == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_107_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6b == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_107_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h6b == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_107_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_107_flits_fired <= _GEN_1388;
      end
    end else begin
      rob_payload_107_flits_fired <= _GEN_1388;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6c == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_108_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6c == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_108_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h6c == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_108_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_108_flits_fired <= _GEN_1389;
      end
    end else begin
      rob_payload_108_flits_fired <= _GEN_1389;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6d == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_109_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6d == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_109_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h6d == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_109_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_109_flits_fired <= _GEN_1390;
      end
    end else begin
      rob_payload_109_flits_fired <= _GEN_1390;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6e == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_110_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6e == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_110_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h6e == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_110_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_110_flits_fired <= _GEN_1391;
      end
    end else begin
      rob_payload_110_flits_fired <= _GEN_1391;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6f == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_111_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6f == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_111_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h6f == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_111_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_111_flits_fired <= _GEN_1392;
      end
    end else begin
      rob_payload_111_flits_fired <= _GEN_1392;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h70 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_112_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h70 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_112_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h70 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_112_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_112_flits_fired <= _GEN_1393;
      end
    end else begin
      rob_payload_112_flits_fired <= _GEN_1393;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h71 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_113_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h71 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_113_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h71 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_113_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_113_flits_fired <= _GEN_1394;
      end
    end else begin
      rob_payload_113_flits_fired <= _GEN_1394;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h72 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_114_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h72 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_114_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h72 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_114_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_114_flits_fired <= _GEN_1395;
      end
    end else begin
      rob_payload_114_flits_fired <= _GEN_1395;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h73 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_115_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h73 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_115_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h73 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_115_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_115_flits_fired <= _GEN_1396;
      end
    end else begin
      rob_payload_115_flits_fired <= _GEN_1396;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h74 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_116_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h74 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_116_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h74 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_116_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_116_flits_fired <= _GEN_1397;
      end
    end else begin
      rob_payload_116_flits_fired <= _GEN_1397;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h75 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_117_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h75 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_117_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h75 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_117_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_117_flits_fired <= _GEN_1398;
      end
    end else begin
      rob_payload_117_flits_fired <= _GEN_1398;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h76 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_118_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h76 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_118_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h76 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_118_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_118_flits_fired <= _GEN_1399;
      end
    end else begin
      rob_payload_118_flits_fired <= _GEN_1399;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h77 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_119_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h77 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_119_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h77 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_119_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_119_flits_fired <= _GEN_1400;
      end
    end else begin
      rob_payload_119_flits_fired <= _GEN_1400;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h78 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_120_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h78 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_120_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h78 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_120_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_120_flits_fired <= _GEN_1401;
      end
    end else begin
      rob_payload_120_flits_fired <= _GEN_1401;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h79 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_121_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h79 == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_121_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h79 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_121_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_121_flits_fired <= _GEN_1402;
      end
    end else begin
      rob_payload_121_flits_fired <= _GEN_1402;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7a == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_122_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7a == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_122_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h7a == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_122_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_122_flits_fired <= _GEN_1403;
      end
    end else begin
      rob_payload_122_flits_fired <= _GEN_1403;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7b == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_123_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7b == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_123_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h7b == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_123_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_123_flits_fired <= _GEN_1404;
      end
    end else begin
      rob_payload_123_flits_fired <= _GEN_1404;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7c == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_124_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7c == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_124_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h7c == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_124_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_124_flits_fired <= _GEN_1405;
      end
    end else begin
      rob_payload_124_flits_fired <= _GEN_1405;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7d == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_125_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7d == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_125_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h7d == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_125_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_125_flits_fired <= _GEN_1406;
      end
    end else begin
      rob_payload_125_flits_fired <= _GEN_1406;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7e == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_126_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7e == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_126_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h7e == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_126_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_126_flits_fired <= _GEN_1407;
      end
    end else begin
      rob_payload_126_flits_fired <= _GEN_1407;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7f == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_127_tsc <= _rob_payload_WIRE_1[63:32]; // @[TestHarness.scala 179:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7f == rob_alloc_ids_0) begin // @[TestHarness.scala 179:36]
        rob_payload_127_rob_idx <= _rob_payload_WIRE_1[31:16]; // @[TestHarness.scala 179:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h7f == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_127_flits_fired <= _rob_payload_flits_fired_T_2; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_127_flits_fired <= _GEN_1408;
      end
    end else begin
      rob_payload_127_flits_fired <= _GEN_1408;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h0 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_0 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_1 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_2 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_3 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_4 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_5 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_6 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_7 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h8 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_8 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h9 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_9 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'ha == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_10 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hb == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_11 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hc == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_12 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hd == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_13 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'he == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_14 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hf == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_15 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h10 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_16 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h11 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_17 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h12 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_18 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h13 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_19 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h14 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_20 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h15 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_21 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h16 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_22 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h17 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_23 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h18 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_24 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h19 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_25 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1a == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_26 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1b == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_27 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1c == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_28 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1d == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_29 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1e == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_30 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1f == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_31 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h20 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_32 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h21 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_33 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h22 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_34 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h23 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_35 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h24 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_36 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h25 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_37 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h26 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_38 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h27 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_39 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h28 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_40 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h29 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_41 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2a == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_42 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2b == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_43 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2c == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_44 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2d == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_45 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2e == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_46 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2f == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_47 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h30 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_48 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h31 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_49 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h32 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_50 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h33 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_51 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h34 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_52 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h35 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_53 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h36 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_54 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h37 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_55 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h38 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_56 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h39 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_57 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3a == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_58 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3b == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_59 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3c == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_60 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3d == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_61 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3e == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_62 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3f == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_63 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h40 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_64 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h41 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_65 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h42 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_66 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h43 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_67 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h44 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_68 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h45 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_69 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h46 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_70 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h47 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_71 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h48 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_72 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h49 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_73 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4a == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_74 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4b == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_75 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4c == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_76 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4d == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_77 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4e == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_78 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4f == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_79 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h50 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_80 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h51 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_81 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h52 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_82 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h53 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_83 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h54 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_84 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h55 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_85 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h56 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_86 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h57 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_87 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h58 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_88 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h59 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_89 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5a == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_90 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5b == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_91 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5c == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_92 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5d == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_93 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5e == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_94 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5f == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_95 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h60 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_96 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h61 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_97 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h62 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_98 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h63 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_99 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h64 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_100 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h65 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_101 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h66 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_102 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h67 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_103 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h68 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_104 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h69 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_105 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6a == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_106 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6b == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_107 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6c == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_108 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6d == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_109 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6e == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_110 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6f == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_111 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h70 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_112 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h71 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_113 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h72 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_114 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h73 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_115 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h74 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_116 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h75 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_117 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h76 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_118 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h77 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_119 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h78 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_120 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h79 == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_121 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7a == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_122 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7b == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_123 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7c == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_124 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7d == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_125 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7e == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_126 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7f == rob_alloc_ids_0) begin // @[TestHarness.scala 182:36]
        rob_n_flits_127 <= _rob_n_flits_T_18; // @[TestHarness.scala 182:36]
      end
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h0 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_0 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_0 <= _GEN_1793;
      end
    end else begin
      rob_flits_returned_0 <= _GEN_1793;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h1 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_1 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_1 <= _GEN_1794;
      end
    end else begin
      rob_flits_returned_1 <= _GEN_1794;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h2 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_2 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_2 <= _GEN_1795;
      end
    end else begin
      rob_flits_returned_2 <= _GEN_1795;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h3 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_3 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_3 <= _GEN_1796;
      end
    end else begin
      rob_flits_returned_3 <= _GEN_1796;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h4 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_4 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_4 <= _GEN_1797;
      end
    end else begin
      rob_flits_returned_4 <= _GEN_1797;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h5 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_5 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_5 <= _GEN_1798;
      end
    end else begin
      rob_flits_returned_5 <= _GEN_1798;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h6 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_6 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_6 <= _GEN_1799;
      end
    end else begin
      rob_flits_returned_6 <= _GEN_1799;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h7 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_7 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_7 <= _GEN_1800;
      end
    end else begin
      rob_flits_returned_7 <= _GEN_1800;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h8 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_8 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_8 <= _GEN_1801;
      end
    end else begin
      rob_flits_returned_8 <= _GEN_1801;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h9 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_9 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_9 <= _GEN_1802;
      end
    end else begin
      rob_flits_returned_9 <= _GEN_1802;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'ha == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_10 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_10 <= _GEN_1803;
      end
    end else begin
      rob_flits_returned_10 <= _GEN_1803;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'hb == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_11 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_11 <= _GEN_1804;
      end
    end else begin
      rob_flits_returned_11 <= _GEN_1804;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'hc == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_12 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_12 <= _GEN_1805;
      end
    end else begin
      rob_flits_returned_12 <= _GEN_1805;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'hd == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_13 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_13 <= _GEN_1806;
      end
    end else begin
      rob_flits_returned_13 <= _GEN_1806;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'he == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_14 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_14 <= _GEN_1807;
      end
    end else begin
      rob_flits_returned_14 <= _GEN_1807;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'hf == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_15 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_15 <= _GEN_1808;
      end
    end else begin
      rob_flits_returned_15 <= _GEN_1808;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h10 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_16 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_16 <= _GEN_1809;
      end
    end else begin
      rob_flits_returned_16 <= _GEN_1809;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h11 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_17 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_17 <= _GEN_1810;
      end
    end else begin
      rob_flits_returned_17 <= _GEN_1810;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h12 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_18 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_18 <= _GEN_1811;
      end
    end else begin
      rob_flits_returned_18 <= _GEN_1811;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h13 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_19 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_19 <= _GEN_1812;
      end
    end else begin
      rob_flits_returned_19 <= _GEN_1812;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h14 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_20 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_20 <= _GEN_1813;
      end
    end else begin
      rob_flits_returned_20 <= _GEN_1813;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h15 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_21 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_21 <= _GEN_1814;
      end
    end else begin
      rob_flits_returned_21 <= _GEN_1814;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h16 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_22 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_22 <= _GEN_1815;
      end
    end else begin
      rob_flits_returned_22 <= _GEN_1815;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h17 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_23 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_23 <= _GEN_1816;
      end
    end else begin
      rob_flits_returned_23 <= _GEN_1816;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h18 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_24 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_24 <= _GEN_1817;
      end
    end else begin
      rob_flits_returned_24 <= _GEN_1817;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h19 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_25 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_25 <= _GEN_1818;
      end
    end else begin
      rob_flits_returned_25 <= _GEN_1818;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h1a == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_26 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_26 <= _GEN_1819;
      end
    end else begin
      rob_flits_returned_26 <= _GEN_1819;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h1b == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_27 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_27 <= _GEN_1820;
      end
    end else begin
      rob_flits_returned_27 <= _GEN_1820;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h1c == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_28 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_28 <= _GEN_1821;
      end
    end else begin
      rob_flits_returned_28 <= _GEN_1821;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h1d == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_29 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_29 <= _GEN_1822;
      end
    end else begin
      rob_flits_returned_29 <= _GEN_1822;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h1e == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_30 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_30 <= _GEN_1823;
      end
    end else begin
      rob_flits_returned_30 <= _GEN_1823;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h1f == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_31 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_31 <= _GEN_1824;
      end
    end else begin
      rob_flits_returned_31 <= _GEN_1824;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h20 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_32 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_32 <= _GEN_1825;
      end
    end else begin
      rob_flits_returned_32 <= _GEN_1825;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h21 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_33 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_33 <= _GEN_1826;
      end
    end else begin
      rob_flits_returned_33 <= _GEN_1826;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h22 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_34 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_34 <= _GEN_1827;
      end
    end else begin
      rob_flits_returned_34 <= _GEN_1827;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h23 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_35 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_35 <= _GEN_1828;
      end
    end else begin
      rob_flits_returned_35 <= _GEN_1828;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h24 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_36 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_36 <= _GEN_1829;
      end
    end else begin
      rob_flits_returned_36 <= _GEN_1829;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h25 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_37 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_37 <= _GEN_1830;
      end
    end else begin
      rob_flits_returned_37 <= _GEN_1830;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h26 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_38 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_38 <= _GEN_1831;
      end
    end else begin
      rob_flits_returned_38 <= _GEN_1831;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h27 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_39 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_39 <= _GEN_1832;
      end
    end else begin
      rob_flits_returned_39 <= _GEN_1832;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h28 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_40 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_40 <= _GEN_1833;
      end
    end else begin
      rob_flits_returned_40 <= _GEN_1833;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h29 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_41 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_41 <= _GEN_1834;
      end
    end else begin
      rob_flits_returned_41 <= _GEN_1834;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h2a == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_42 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_42 <= _GEN_1835;
      end
    end else begin
      rob_flits_returned_42 <= _GEN_1835;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h2b == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_43 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_43 <= _GEN_1836;
      end
    end else begin
      rob_flits_returned_43 <= _GEN_1836;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h2c == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_44 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_44 <= _GEN_1837;
      end
    end else begin
      rob_flits_returned_44 <= _GEN_1837;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h2d == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_45 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_45 <= _GEN_1838;
      end
    end else begin
      rob_flits_returned_45 <= _GEN_1838;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h2e == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_46 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_46 <= _GEN_1839;
      end
    end else begin
      rob_flits_returned_46 <= _GEN_1839;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h2f == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_47 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_47 <= _GEN_1840;
      end
    end else begin
      rob_flits_returned_47 <= _GEN_1840;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h30 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_48 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_48 <= _GEN_1841;
      end
    end else begin
      rob_flits_returned_48 <= _GEN_1841;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h31 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_49 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_49 <= _GEN_1842;
      end
    end else begin
      rob_flits_returned_49 <= _GEN_1842;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h32 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_50 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_50 <= _GEN_1843;
      end
    end else begin
      rob_flits_returned_50 <= _GEN_1843;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h33 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_51 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_51 <= _GEN_1844;
      end
    end else begin
      rob_flits_returned_51 <= _GEN_1844;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h34 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_52 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_52 <= _GEN_1845;
      end
    end else begin
      rob_flits_returned_52 <= _GEN_1845;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h35 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_53 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_53 <= _GEN_1846;
      end
    end else begin
      rob_flits_returned_53 <= _GEN_1846;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h36 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_54 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_54 <= _GEN_1847;
      end
    end else begin
      rob_flits_returned_54 <= _GEN_1847;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h37 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_55 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_55 <= _GEN_1848;
      end
    end else begin
      rob_flits_returned_55 <= _GEN_1848;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h38 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_56 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_56 <= _GEN_1849;
      end
    end else begin
      rob_flits_returned_56 <= _GEN_1849;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h39 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_57 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_57 <= _GEN_1850;
      end
    end else begin
      rob_flits_returned_57 <= _GEN_1850;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h3a == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_58 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_58 <= _GEN_1851;
      end
    end else begin
      rob_flits_returned_58 <= _GEN_1851;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h3b == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_59 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_59 <= _GEN_1852;
      end
    end else begin
      rob_flits_returned_59 <= _GEN_1852;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h3c == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_60 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_60 <= _GEN_1853;
      end
    end else begin
      rob_flits_returned_60 <= _GEN_1853;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h3d == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_61 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_61 <= _GEN_1854;
      end
    end else begin
      rob_flits_returned_61 <= _GEN_1854;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h3e == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_62 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_62 <= _GEN_1855;
      end
    end else begin
      rob_flits_returned_62 <= _GEN_1855;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h3f == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_63 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_63 <= _GEN_1856;
      end
    end else begin
      rob_flits_returned_63 <= _GEN_1856;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h40 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_64 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_64 <= _GEN_1857;
      end
    end else begin
      rob_flits_returned_64 <= _GEN_1857;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h41 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_65 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_65 <= _GEN_1858;
      end
    end else begin
      rob_flits_returned_65 <= _GEN_1858;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h42 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_66 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_66 <= _GEN_1859;
      end
    end else begin
      rob_flits_returned_66 <= _GEN_1859;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h43 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_67 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_67 <= _GEN_1860;
      end
    end else begin
      rob_flits_returned_67 <= _GEN_1860;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h44 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_68 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_68 <= _GEN_1861;
      end
    end else begin
      rob_flits_returned_68 <= _GEN_1861;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h45 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_69 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_69 <= _GEN_1862;
      end
    end else begin
      rob_flits_returned_69 <= _GEN_1862;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h46 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_70 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_70 <= _GEN_1863;
      end
    end else begin
      rob_flits_returned_70 <= _GEN_1863;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h47 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_71 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_71 <= _GEN_1864;
      end
    end else begin
      rob_flits_returned_71 <= _GEN_1864;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h48 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_72 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_72 <= _GEN_1865;
      end
    end else begin
      rob_flits_returned_72 <= _GEN_1865;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h49 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_73 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_73 <= _GEN_1866;
      end
    end else begin
      rob_flits_returned_73 <= _GEN_1866;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h4a == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_74 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_74 <= _GEN_1867;
      end
    end else begin
      rob_flits_returned_74 <= _GEN_1867;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h4b == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_75 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_75 <= _GEN_1868;
      end
    end else begin
      rob_flits_returned_75 <= _GEN_1868;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h4c == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_76 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_76 <= _GEN_1869;
      end
    end else begin
      rob_flits_returned_76 <= _GEN_1869;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h4d == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_77 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_77 <= _GEN_1870;
      end
    end else begin
      rob_flits_returned_77 <= _GEN_1870;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h4e == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_78 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_78 <= _GEN_1871;
      end
    end else begin
      rob_flits_returned_78 <= _GEN_1871;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h4f == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_79 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_79 <= _GEN_1872;
      end
    end else begin
      rob_flits_returned_79 <= _GEN_1872;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h50 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_80 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_80 <= _GEN_1873;
      end
    end else begin
      rob_flits_returned_80 <= _GEN_1873;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h51 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_81 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_81 <= _GEN_1874;
      end
    end else begin
      rob_flits_returned_81 <= _GEN_1874;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h52 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_82 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_82 <= _GEN_1875;
      end
    end else begin
      rob_flits_returned_82 <= _GEN_1875;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h53 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_83 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_83 <= _GEN_1876;
      end
    end else begin
      rob_flits_returned_83 <= _GEN_1876;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h54 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_84 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_84 <= _GEN_1877;
      end
    end else begin
      rob_flits_returned_84 <= _GEN_1877;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h55 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_85 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_85 <= _GEN_1878;
      end
    end else begin
      rob_flits_returned_85 <= _GEN_1878;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h56 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_86 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_86 <= _GEN_1879;
      end
    end else begin
      rob_flits_returned_86 <= _GEN_1879;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h57 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_87 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_87 <= _GEN_1880;
      end
    end else begin
      rob_flits_returned_87 <= _GEN_1880;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h58 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_88 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_88 <= _GEN_1881;
      end
    end else begin
      rob_flits_returned_88 <= _GEN_1881;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h59 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_89 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_89 <= _GEN_1882;
      end
    end else begin
      rob_flits_returned_89 <= _GEN_1882;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h5a == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_90 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_90 <= _GEN_1883;
      end
    end else begin
      rob_flits_returned_90 <= _GEN_1883;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h5b == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_91 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_91 <= _GEN_1884;
      end
    end else begin
      rob_flits_returned_91 <= _GEN_1884;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h5c == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_92 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_92 <= _GEN_1885;
      end
    end else begin
      rob_flits_returned_92 <= _GEN_1885;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h5d == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_93 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_93 <= _GEN_1886;
      end
    end else begin
      rob_flits_returned_93 <= _GEN_1886;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h5e == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_94 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_94 <= _GEN_1887;
      end
    end else begin
      rob_flits_returned_94 <= _GEN_1887;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h5f == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_95 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_95 <= _GEN_1888;
      end
    end else begin
      rob_flits_returned_95 <= _GEN_1888;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h60 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_96 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_96 <= _GEN_1889;
      end
    end else begin
      rob_flits_returned_96 <= _GEN_1889;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h61 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_97 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_97 <= _GEN_1890;
      end
    end else begin
      rob_flits_returned_97 <= _GEN_1890;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h62 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_98 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_98 <= _GEN_1891;
      end
    end else begin
      rob_flits_returned_98 <= _GEN_1891;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h63 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_99 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_99 <= _GEN_1892;
      end
    end else begin
      rob_flits_returned_99 <= _GEN_1892;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h64 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_100 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_100 <= _GEN_1893;
      end
    end else begin
      rob_flits_returned_100 <= _GEN_1893;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h65 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_101 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_101 <= _GEN_1894;
      end
    end else begin
      rob_flits_returned_101 <= _GEN_1894;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h66 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_102 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_102 <= _GEN_1895;
      end
    end else begin
      rob_flits_returned_102 <= _GEN_1895;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h67 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_103 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_103 <= _GEN_1896;
      end
    end else begin
      rob_flits_returned_103 <= _GEN_1896;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h68 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_104 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_104 <= _GEN_1897;
      end
    end else begin
      rob_flits_returned_104 <= _GEN_1897;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h69 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_105 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_105 <= _GEN_1898;
      end
    end else begin
      rob_flits_returned_105 <= _GEN_1898;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h6a == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_106 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_106 <= _GEN_1899;
      end
    end else begin
      rob_flits_returned_106 <= _GEN_1899;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h6b == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_107 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_107 <= _GEN_1900;
      end
    end else begin
      rob_flits_returned_107 <= _GEN_1900;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h6c == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_108 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_108 <= _GEN_1901;
      end
    end else begin
      rob_flits_returned_108 <= _GEN_1901;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h6d == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_109 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_109 <= _GEN_1902;
      end
    end else begin
      rob_flits_returned_109 <= _GEN_1902;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h6e == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_110 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_110 <= _GEN_1903;
      end
    end else begin
      rob_flits_returned_110 <= _GEN_1903;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h6f == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_111 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_111 <= _GEN_1904;
      end
    end else begin
      rob_flits_returned_111 <= _GEN_1904;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h70 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_112 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_112 <= _GEN_1905;
      end
    end else begin
      rob_flits_returned_112 <= _GEN_1905;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h71 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_113 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_113 <= _GEN_1906;
      end
    end else begin
      rob_flits_returned_113 <= _GEN_1906;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h72 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_114 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_114 <= _GEN_1907;
      end
    end else begin
      rob_flits_returned_114 <= _GEN_1907;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h73 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_115 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_115 <= _GEN_1908;
      end
    end else begin
      rob_flits_returned_115 <= _GEN_1908;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h74 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_116 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_116 <= _GEN_1909;
      end
    end else begin
      rob_flits_returned_116 <= _GEN_1909;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h75 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_117 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_117 <= _GEN_1910;
      end
    end else begin
      rob_flits_returned_117 <= _GEN_1910;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h76 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_118 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_118 <= _GEN_1911;
      end
    end else begin
      rob_flits_returned_118 <= _GEN_1911;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h77 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_119 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_119 <= _GEN_1912;
      end
    end else begin
      rob_flits_returned_119 <= _GEN_1912;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h78 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_120 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_120 <= _GEN_1913;
      end
    end else begin
      rob_flits_returned_120 <= _GEN_1913;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h79 == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_121 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_121 <= _GEN_1914;
      end
    end else begin
      rob_flits_returned_121 <= _GEN_1914;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h7a == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_122 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_122 <= _GEN_1915;
      end
    end else begin
      rob_flits_returned_122 <= _GEN_1915;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h7b == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_123 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_123 <= _GEN_1916;
      end
    end else begin
      rob_flits_returned_123 <= _GEN_1916;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h7c == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_124 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_124 <= _GEN_1917;
      end
    end else begin
      rob_flits_returned_124 <= _GEN_1917;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h7d == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_125 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_125 <= _GEN_1918;
      end
    end else begin
      rob_flits_returned_125 <= _GEN_1918;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h7e == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_126 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_126 <= _GEN_1919;
      end
    end else begin
      rob_flits_returned_126 <= _GEN_1919;
    end
    if (_T_67) begin // @[TestHarness.scala 199:26]
      if (7'h7f == out_payload_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_127 <= _rob_flits_returned_T_2; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_127 <= _GEN_1920;
      end
    end else begin
      rob_flits_returned_127 <= _GEN_1920;
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h0 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_0 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_1 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_2 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_3 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_4 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_5 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_6 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_7 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h8 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_8 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h9 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_9 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'ha == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_10 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hb == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_11 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hc == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_12 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hd == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_13 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'he == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_14 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hf == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_15 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h10 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_16 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h11 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_17 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h12 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_18 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h13 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_19 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h14 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_20 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h15 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_21 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h16 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_22 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h17 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_23 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h18 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_24 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h19 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_25 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1a == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_26 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1b == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_27 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1c == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_28 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1d == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_29 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1e == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_30 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1f == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_31 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h20 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_32 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h21 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_33 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h22 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_34 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h23 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_35 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h24 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_36 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h25 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_37 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h26 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_38 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h27 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_39 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h28 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_40 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h29 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_41 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2a == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_42 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2b == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_43 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2c == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_44 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2d == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_45 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2e == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_46 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2f == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_47 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h30 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_48 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h31 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_49 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h32 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_50 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h33 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_51 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h34 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_52 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h35 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_53 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h36 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_54 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h37 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_55 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h38 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_56 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h39 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_57 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3a == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_58 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3b == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_59 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3c == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_60 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3d == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_61 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3e == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_62 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3f == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_63 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h40 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_64 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h41 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_65 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h42 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_66 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h43 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_67 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h44 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_68 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h45 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_69 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h46 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_70 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h47 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_71 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h48 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_72 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h49 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_73 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4a == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_74 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4b == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_75 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4c == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_76 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4d == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_77 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4e == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_78 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4f == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_79 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h50 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_80 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h51 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_81 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h52 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_82 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h53 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_83 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h54 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_84 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h55 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_85 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h56 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_86 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h57 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_87 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h58 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_88 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h59 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_89 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5a == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_90 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5b == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_91 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5c == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_92 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5d == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_93 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5e == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_94 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5f == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_95 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h60 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_96 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h61 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_97 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h62 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_98 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h63 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_99 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h64 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_100 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h65 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_101 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h66 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_102 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h67 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_103 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h68 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_104 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h69 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_105 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6a == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_106 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6b == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_107 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6c == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_108 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6d == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_109 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6e == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_110 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6f == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_111 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h70 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_112 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h71 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_113 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h72 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_114 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h73 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_115 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h74 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_116 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h75 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_117 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h76 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_118 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h77 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_119 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h78 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_120 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h79 == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_121 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7a == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_122 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7b == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_123 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7c == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_124 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7d == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_125 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7e == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_126 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7f == rob_alloc_ids_0) begin // @[TestHarness.scala 184:36]
        rob_tscs_127 <= _rob_tscs_T_22; // @[TestHarness.scala 184:36]
      end
    end
    if (reset) begin // @[TestHarness.scala 164:24]
      io_success_REG <= 1'h0; // @[TestHarness.scala 164:24]
    end else begin
      io_success_REG <= success; // @[TestHarness.scala 164:24]
    end
    if (reset) begin // @[TestHarness.scala 196:31]
      packet_valid <= 1'h0; // @[TestHarness.scala 196:31]
    end else if (_T_67) begin // @[TestHarness.scala 199:26]
      if (io_from_noc_0_flit_bits_tail) begin // @[TestHarness.scala 216:31]
        packet_valid <= 1'h0; // @[TestHarness.scala 216:46]
      end else begin
        packet_valid <= _GEN_3585;
      end
    end
    packet_rob_idx <= _GEN_3845[6:0];
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~idle_counter[10])) begin
          $fwrite(32'h80000002,"Assertion failed\n    at TestHarness.scala:148 assert(!idle_counter(10))\n"); // @[TestHarness.scala 148:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (success & _T_3) begin
          $fwrite(32'h80000002,"%d flits, %d cycles\n",flits,tsc); // @[TestHarness.scala 166:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_67 & _T_3 & ~_T_25[0]) begin
          $fwrite(32'h80000002,
            "Assertion failed: out[0] unexpected response\n    at TestHarness.scala:201 assert(rob_valids(rob_idx), cf\"out[${i.toString}] unexpected response\")\n"
            ); // @[TestHarness.scala 201:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_518 & ~(_T_31 == io_from_noc_0_flit_bits_payload)) begin
          $fwrite(32'h80000002,
            "Assertion failed: out[0] incorrect payload\n    at TestHarness.scala:202 assert(rob_payload(rob_idx).asUInt === o.flit.bits.payload.asUInt, cf\"out[${i.toString}] incorrect payload\");\n"
            ); // @[TestHarness.scala 202:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_518 & ~(~io_from_noc_0_flit_bits_ingress_id)) begin
          $fwrite(32'h80000002,
            "Assertion failed: out[0] incorrect source\n    at TestHarness.scala:203 assert(o.flit.bits.ingress_id === rob_ingress_id(rob_idx), cf\"out[${i.toString}] incorrect source\")\n"
            ); // @[TestHarness.scala 203:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_518 & ~(_GEN_2816 < _GEN_2944)) begin
          $fwrite(32'h80000002,
            "Assertion failed: out[0] too many flits returned\n    at TestHarness.scala:205 assert(rob_flits_returned(rob_idx) < rob_n_flits(rob_idx), cf\"out[${i.toString}] too many flits returned\")\n"
            ); // @[TestHarness.scala 205:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_518 & ~(~packet_valid & io_from_noc_0_flit_bits_head | out_payload_rob_idx == _GEN_385)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at TestHarness.scala:206 assert((!packet_valid && o.flit.bits.head) || rob_idx === packet_rob_idx)\n"
            ); // @[TestHarness.scala 206:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_67 & _T_59 & _T_3) begin
          $fwrite(32'h80000002,"%d, 0, %d\n",1'h0,tsc - out_payload_tsc); // @[TestHarness.scala 210:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[0] & _T_3 & ~(_T_72 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 0 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[1] & _T_3 & ~(_T_79 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 1 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[2] & _T_3 & ~(_T_86 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 2 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[3] & _T_3 & ~(_T_93 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 3 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[4] & _T_3 & ~(_T_100 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 4 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[5] & _T_3 & ~(_T_107 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 5 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[6] & _T_3 & ~(_T_114 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 6 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[7] & _T_3 & ~(_T_121 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 7 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[8] & _T_3 & ~(_T_128 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 8 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[9] & _T_3 & ~(_T_135 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 9 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[10] & _T_3 & ~(_T_142 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 10 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[11] & _T_3 & ~(_T_149 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 11 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[12] & _T_3 & ~(_T_156 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 12 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[13] & _T_3 & ~(_T_163 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 13 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[14] & _T_3 & ~(_T_170 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 14 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[15] & _T_3 & ~(_T_177 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 15 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[16] & _T_3 & ~(_T_184 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 16 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[17] & _T_3 & ~(_T_191 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 17 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[18] & _T_3 & ~(_T_198 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 18 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[19] & _T_3 & ~(_T_205 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 19 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[20] & _T_3 & ~(_T_212 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 20 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[21] & _T_3 & ~(_T_219 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 21 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[22] & _T_3 & ~(_T_226 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 22 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[23] & _T_3 & ~(_T_233 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 23 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[24] & _T_3 & ~(_T_240 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 24 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[25] & _T_3 & ~(_T_247 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 25 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[26] & _T_3 & ~(_T_254 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 26 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[27] & _T_3 & ~(_T_261 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 27 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[28] & _T_3 & ~(_T_268 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 28 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[29] & _T_3 & ~(_T_275 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 29 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[30] & _T_3 & ~(_T_282 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 30 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[31] & _T_3 & ~(_T_289 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 31 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[32] & _T_3 & ~(_T_296 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 32 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[33] & _T_3 & ~(_T_303 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 33 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[34] & _T_3 & ~(_T_310 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 34 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[35] & _T_3 & ~(_T_317 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 35 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[36] & _T_3 & ~(_T_324 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 36 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[37] & _T_3 & ~(_T_331 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 37 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[38] & _T_3 & ~(_T_338 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 38 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[39] & _T_3 & ~(_T_345 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 39 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[40] & _T_3 & ~(_T_352 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 40 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[41] & _T_3 & ~(_T_359 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 41 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[42] & _T_3 & ~(_T_366 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 42 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[43] & _T_3 & ~(_T_373 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 43 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[44] & _T_3 & ~(_T_380 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 44 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[45] & _T_3 & ~(_T_387 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 45 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[46] & _T_3 & ~(_T_394 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 46 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[47] & _T_3 & ~(_T_401 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 47 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[48] & _T_3 & ~(_T_408 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 48 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[49] & _T_3 & ~(_T_415 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 49 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[50] & _T_3 & ~(_T_422 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 50 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[51] & _T_3 & ~(_T_429 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 51 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[52] & _T_3 & ~(_T_436 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 52 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[53] & _T_3 & ~(_T_443 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 53 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[54] & _T_3 & ~(_T_450 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 54 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[55] & _T_3 & ~(_T_457 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 55 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[56] & _T_3 & ~(_T_464 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 56 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[57] & _T_3 & ~(_T_471 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 57 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[58] & _T_3 & ~(_T_478 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 58 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[59] & _T_3 & ~(_T_485 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 59 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[60] & _T_3 & ~(_T_492 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 60 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[61] & _T_3 & ~(_T_499 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 61 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[62] & _T_3 & ~(_T_506 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 62 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[63] & _T_3 & ~(_T_513 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 63 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[64] & _T_3 & ~(_T_520 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 64 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[65] & _T_3 & ~(_T_527 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 65 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[66] & _T_3 & ~(_T_534 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 66 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[67] & _T_3 & ~(_T_541 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 67 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[68] & _T_3 & ~(_T_548 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 68 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[69] & _T_3 & ~(_T_555 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 69 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[70] & _T_3 & ~(_T_562 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 70 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[71] & _T_3 & ~(_T_569 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 71 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[72] & _T_3 & ~(_T_576 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 72 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[73] & _T_3 & ~(_T_583 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 73 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[74] & _T_3 & ~(_T_590 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 74 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[75] & _T_3 & ~(_T_597 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 75 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[76] & _T_3 & ~(_T_604 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 76 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[77] & _T_3 & ~(_T_611 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 77 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[78] & _T_3 & ~(_T_618 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 78 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[79] & _T_3 & ~(_T_625 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 79 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[80] & _T_3 & ~(_T_632 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 80 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[81] & _T_3 & ~(_T_639 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 81 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[82] & _T_3 & ~(_T_646 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 82 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[83] & _T_3 & ~(_T_653 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 83 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[84] & _T_3 & ~(_T_660 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 84 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[85] & _T_3 & ~(_T_667 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 85 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[86] & _T_3 & ~(_T_674 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 86 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[87] & _T_3 & ~(_T_681 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 87 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[88] & _T_3 & ~(_T_688 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 88 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[89] & _T_3 & ~(_T_695 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 89 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[90] & _T_3 & ~(_T_702 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 90 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[91] & _T_3 & ~(_T_709 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 91 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[92] & _T_3 & ~(_T_716 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 92 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[93] & _T_3 & ~(_T_723 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 93 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[94] & _T_3 & ~(_T_730 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 94 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[95] & _T_3 & ~(_T_737 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 95 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[96] & _T_3 & ~(_T_744 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 96 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[97] & _T_3 & ~(_T_751 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 97 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[98] & _T_3 & ~(_T_758 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 98 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[99] & _T_3 & ~(_T_765 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 99 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[100] & _T_3 & ~(_T_772 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 100 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[101] & _T_3 & ~(_T_779 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 101 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[102] & _T_3 & ~(_T_786 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 102 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[103] & _T_3 & ~(_T_793 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 103 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[104] & _T_3 & ~(_T_800 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 104 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[105] & _T_3 & ~(_T_807 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 105 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[106] & _T_3 & ~(_T_814 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 106 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[107] & _T_3 & ~(_T_821 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 107 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[108] & _T_3 & ~(_T_828 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 108 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[109] & _T_3 & ~(_T_835 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 109 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[110] & _T_3 & ~(_T_842 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 110 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[111] & _T_3 & ~(_T_849 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 111 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[112] & _T_3 & ~(_T_856 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 112 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[113] & _T_3 & ~(_T_863 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 113 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[114] & _T_3 & ~(_T_870 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 114 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[115] & _T_3 & ~(_T_877 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 115 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[116] & _T_3 & ~(_T_884 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 116 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[117] & _T_3 & ~(_T_891 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 117 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[118] & _T_3 & ~(_T_898 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 118 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[119] & _T_3 & ~(_T_905 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 119 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[120] & _T_3 & ~(_T_912 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 120 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[121] & _T_3 & ~(_T_919 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 121 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[122] & _T_3 & ~(_T_926 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 122 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[123] & _T_3 & ~(_T_933 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 123 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[124] & _T_3 & ~(_T_940 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 124 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[125] & _T_3 & ~(_T_947 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 125 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[126] & _T_3 & ~(_T_954 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 126 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[127] & _T_3 & ~(_T_961 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 127 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  txs = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  flits = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  tsc = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  idle_counter = _RAND_3[10:0];
  _RAND_4 = {4{`RANDOM}};
  rob_valids = _RAND_4[127:0];
  _RAND_5 = {1{`RANDOM}};
  rob_payload_0_tsc = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  rob_payload_0_rob_idx = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  rob_payload_0_flits_fired = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  rob_payload_1_tsc = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  rob_payload_1_rob_idx = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  rob_payload_1_flits_fired = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  rob_payload_2_tsc = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  rob_payload_2_rob_idx = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  rob_payload_2_flits_fired = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  rob_payload_3_tsc = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  rob_payload_3_rob_idx = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  rob_payload_3_flits_fired = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  rob_payload_4_tsc = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  rob_payload_4_rob_idx = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  rob_payload_4_flits_fired = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  rob_payload_5_tsc = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  rob_payload_5_rob_idx = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  rob_payload_5_flits_fired = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  rob_payload_6_tsc = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  rob_payload_6_rob_idx = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  rob_payload_6_flits_fired = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  rob_payload_7_tsc = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  rob_payload_7_rob_idx = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  rob_payload_7_flits_fired = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  rob_payload_8_tsc = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  rob_payload_8_rob_idx = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  rob_payload_8_flits_fired = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  rob_payload_9_tsc = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  rob_payload_9_rob_idx = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  rob_payload_9_flits_fired = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  rob_payload_10_tsc = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  rob_payload_10_rob_idx = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  rob_payload_10_flits_fired = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  rob_payload_11_tsc = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  rob_payload_11_rob_idx = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  rob_payload_11_flits_fired = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  rob_payload_12_tsc = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  rob_payload_12_rob_idx = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  rob_payload_12_flits_fired = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  rob_payload_13_tsc = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  rob_payload_13_rob_idx = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  rob_payload_13_flits_fired = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  rob_payload_14_tsc = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  rob_payload_14_rob_idx = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  rob_payload_14_flits_fired = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  rob_payload_15_tsc = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  rob_payload_15_rob_idx = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  rob_payload_15_flits_fired = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  rob_payload_16_tsc = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  rob_payload_16_rob_idx = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  rob_payload_16_flits_fired = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  rob_payload_17_tsc = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  rob_payload_17_rob_idx = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  rob_payload_17_flits_fired = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  rob_payload_18_tsc = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  rob_payload_18_rob_idx = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  rob_payload_18_flits_fired = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  rob_payload_19_tsc = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  rob_payload_19_rob_idx = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  rob_payload_19_flits_fired = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  rob_payload_20_tsc = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  rob_payload_20_rob_idx = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  rob_payload_20_flits_fired = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  rob_payload_21_tsc = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  rob_payload_21_rob_idx = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  rob_payload_21_flits_fired = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  rob_payload_22_tsc = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  rob_payload_22_rob_idx = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  rob_payload_22_flits_fired = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  rob_payload_23_tsc = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  rob_payload_23_rob_idx = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  rob_payload_23_flits_fired = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  rob_payload_24_tsc = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  rob_payload_24_rob_idx = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  rob_payload_24_flits_fired = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  rob_payload_25_tsc = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  rob_payload_25_rob_idx = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  rob_payload_25_flits_fired = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  rob_payload_26_tsc = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  rob_payload_26_rob_idx = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  rob_payload_26_flits_fired = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  rob_payload_27_tsc = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  rob_payload_27_rob_idx = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  rob_payload_27_flits_fired = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  rob_payload_28_tsc = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  rob_payload_28_rob_idx = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  rob_payload_28_flits_fired = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  rob_payload_29_tsc = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  rob_payload_29_rob_idx = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  rob_payload_29_flits_fired = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  rob_payload_30_tsc = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  rob_payload_30_rob_idx = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  rob_payload_30_flits_fired = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  rob_payload_31_tsc = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  rob_payload_31_rob_idx = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  rob_payload_31_flits_fired = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  rob_payload_32_tsc = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  rob_payload_32_rob_idx = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  rob_payload_32_flits_fired = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  rob_payload_33_tsc = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  rob_payload_33_rob_idx = _RAND_105[15:0];
  _RAND_106 = {1{`RANDOM}};
  rob_payload_33_flits_fired = _RAND_106[15:0];
  _RAND_107 = {1{`RANDOM}};
  rob_payload_34_tsc = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  rob_payload_34_rob_idx = _RAND_108[15:0];
  _RAND_109 = {1{`RANDOM}};
  rob_payload_34_flits_fired = _RAND_109[15:0];
  _RAND_110 = {1{`RANDOM}};
  rob_payload_35_tsc = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  rob_payload_35_rob_idx = _RAND_111[15:0];
  _RAND_112 = {1{`RANDOM}};
  rob_payload_35_flits_fired = _RAND_112[15:0];
  _RAND_113 = {1{`RANDOM}};
  rob_payload_36_tsc = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  rob_payload_36_rob_idx = _RAND_114[15:0];
  _RAND_115 = {1{`RANDOM}};
  rob_payload_36_flits_fired = _RAND_115[15:0];
  _RAND_116 = {1{`RANDOM}};
  rob_payload_37_tsc = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  rob_payload_37_rob_idx = _RAND_117[15:0];
  _RAND_118 = {1{`RANDOM}};
  rob_payload_37_flits_fired = _RAND_118[15:0];
  _RAND_119 = {1{`RANDOM}};
  rob_payload_38_tsc = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  rob_payload_38_rob_idx = _RAND_120[15:0];
  _RAND_121 = {1{`RANDOM}};
  rob_payload_38_flits_fired = _RAND_121[15:0];
  _RAND_122 = {1{`RANDOM}};
  rob_payload_39_tsc = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  rob_payload_39_rob_idx = _RAND_123[15:0];
  _RAND_124 = {1{`RANDOM}};
  rob_payload_39_flits_fired = _RAND_124[15:0];
  _RAND_125 = {1{`RANDOM}};
  rob_payload_40_tsc = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  rob_payload_40_rob_idx = _RAND_126[15:0];
  _RAND_127 = {1{`RANDOM}};
  rob_payload_40_flits_fired = _RAND_127[15:0];
  _RAND_128 = {1{`RANDOM}};
  rob_payload_41_tsc = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  rob_payload_41_rob_idx = _RAND_129[15:0];
  _RAND_130 = {1{`RANDOM}};
  rob_payload_41_flits_fired = _RAND_130[15:0];
  _RAND_131 = {1{`RANDOM}};
  rob_payload_42_tsc = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  rob_payload_42_rob_idx = _RAND_132[15:0];
  _RAND_133 = {1{`RANDOM}};
  rob_payload_42_flits_fired = _RAND_133[15:0];
  _RAND_134 = {1{`RANDOM}};
  rob_payload_43_tsc = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  rob_payload_43_rob_idx = _RAND_135[15:0];
  _RAND_136 = {1{`RANDOM}};
  rob_payload_43_flits_fired = _RAND_136[15:0];
  _RAND_137 = {1{`RANDOM}};
  rob_payload_44_tsc = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  rob_payload_44_rob_idx = _RAND_138[15:0];
  _RAND_139 = {1{`RANDOM}};
  rob_payload_44_flits_fired = _RAND_139[15:0];
  _RAND_140 = {1{`RANDOM}};
  rob_payload_45_tsc = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  rob_payload_45_rob_idx = _RAND_141[15:0];
  _RAND_142 = {1{`RANDOM}};
  rob_payload_45_flits_fired = _RAND_142[15:0];
  _RAND_143 = {1{`RANDOM}};
  rob_payload_46_tsc = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  rob_payload_46_rob_idx = _RAND_144[15:0];
  _RAND_145 = {1{`RANDOM}};
  rob_payload_46_flits_fired = _RAND_145[15:0];
  _RAND_146 = {1{`RANDOM}};
  rob_payload_47_tsc = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  rob_payload_47_rob_idx = _RAND_147[15:0];
  _RAND_148 = {1{`RANDOM}};
  rob_payload_47_flits_fired = _RAND_148[15:0];
  _RAND_149 = {1{`RANDOM}};
  rob_payload_48_tsc = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  rob_payload_48_rob_idx = _RAND_150[15:0];
  _RAND_151 = {1{`RANDOM}};
  rob_payload_48_flits_fired = _RAND_151[15:0];
  _RAND_152 = {1{`RANDOM}};
  rob_payload_49_tsc = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  rob_payload_49_rob_idx = _RAND_153[15:0];
  _RAND_154 = {1{`RANDOM}};
  rob_payload_49_flits_fired = _RAND_154[15:0];
  _RAND_155 = {1{`RANDOM}};
  rob_payload_50_tsc = _RAND_155[31:0];
  _RAND_156 = {1{`RANDOM}};
  rob_payload_50_rob_idx = _RAND_156[15:0];
  _RAND_157 = {1{`RANDOM}};
  rob_payload_50_flits_fired = _RAND_157[15:0];
  _RAND_158 = {1{`RANDOM}};
  rob_payload_51_tsc = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  rob_payload_51_rob_idx = _RAND_159[15:0];
  _RAND_160 = {1{`RANDOM}};
  rob_payload_51_flits_fired = _RAND_160[15:0];
  _RAND_161 = {1{`RANDOM}};
  rob_payload_52_tsc = _RAND_161[31:0];
  _RAND_162 = {1{`RANDOM}};
  rob_payload_52_rob_idx = _RAND_162[15:0];
  _RAND_163 = {1{`RANDOM}};
  rob_payload_52_flits_fired = _RAND_163[15:0];
  _RAND_164 = {1{`RANDOM}};
  rob_payload_53_tsc = _RAND_164[31:0];
  _RAND_165 = {1{`RANDOM}};
  rob_payload_53_rob_idx = _RAND_165[15:0];
  _RAND_166 = {1{`RANDOM}};
  rob_payload_53_flits_fired = _RAND_166[15:0];
  _RAND_167 = {1{`RANDOM}};
  rob_payload_54_tsc = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  rob_payload_54_rob_idx = _RAND_168[15:0];
  _RAND_169 = {1{`RANDOM}};
  rob_payload_54_flits_fired = _RAND_169[15:0];
  _RAND_170 = {1{`RANDOM}};
  rob_payload_55_tsc = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  rob_payload_55_rob_idx = _RAND_171[15:0];
  _RAND_172 = {1{`RANDOM}};
  rob_payload_55_flits_fired = _RAND_172[15:0];
  _RAND_173 = {1{`RANDOM}};
  rob_payload_56_tsc = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  rob_payload_56_rob_idx = _RAND_174[15:0];
  _RAND_175 = {1{`RANDOM}};
  rob_payload_56_flits_fired = _RAND_175[15:0];
  _RAND_176 = {1{`RANDOM}};
  rob_payload_57_tsc = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  rob_payload_57_rob_idx = _RAND_177[15:0];
  _RAND_178 = {1{`RANDOM}};
  rob_payload_57_flits_fired = _RAND_178[15:0];
  _RAND_179 = {1{`RANDOM}};
  rob_payload_58_tsc = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  rob_payload_58_rob_idx = _RAND_180[15:0];
  _RAND_181 = {1{`RANDOM}};
  rob_payload_58_flits_fired = _RAND_181[15:0];
  _RAND_182 = {1{`RANDOM}};
  rob_payload_59_tsc = _RAND_182[31:0];
  _RAND_183 = {1{`RANDOM}};
  rob_payload_59_rob_idx = _RAND_183[15:0];
  _RAND_184 = {1{`RANDOM}};
  rob_payload_59_flits_fired = _RAND_184[15:0];
  _RAND_185 = {1{`RANDOM}};
  rob_payload_60_tsc = _RAND_185[31:0];
  _RAND_186 = {1{`RANDOM}};
  rob_payload_60_rob_idx = _RAND_186[15:0];
  _RAND_187 = {1{`RANDOM}};
  rob_payload_60_flits_fired = _RAND_187[15:0];
  _RAND_188 = {1{`RANDOM}};
  rob_payload_61_tsc = _RAND_188[31:0];
  _RAND_189 = {1{`RANDOM}};
  rob_payload_61_rob_idx = _RAND_189[15:0];
  _RAND_190 = {1{`RANDOM}};
  rob_payload_61_flits_fired = _RAND_190[15:0];
  _RAND_191 = {1{`RANDOM}};
  rob_payload_62_tsc = _RAND_191[31:0];
  _RAND_192 = {1{`RANDOM}};
  rob_payload_62_rob_idx = _RAND_192[15:0];
  _RAND_193 = {1{`RANDOM}};
  rob_payload_62_flits_fired = _RAND_193[15:0];
  _RAND_194 = {1{`RANDOM}};
  rob_payload_63_tsc = _RAND_194[31:0];
  _RAND_195 = {1{`RANDOM}};
  rob_payload_63_rob_idx = _RAND_195[15:0];
  _RAND_196 = {1{`RANDOM}};
  rob_payload_63_flits_fired = _RAND_196[15:0];
  _RAND_197 = {1{`RANDOM}};
  rob_payload_64_tsc = _RAND_197[31:0];
  _RAND_198 = {1{`RANDOM}};
  rob_payload_64_rob_idx = _RAND_198[15:0];
  _RAND_199 = {1{`RANDOM}};
  rob_payload_64_flits_fired = _RAND_199[15:0];
  _RAND_200 = {1{`RANDOM}};
  rob_payload_65_tsc = _RAND_200[31:0];
  _RAND_201 = {1{`RANDOM}};
  rob_payload_65_rob_idx = _RAND_201[15:0];
  _RAND_202 = {1{`RANDOM}};
  rob_payload_65_flits_fired = _RAND_202[15:0];
  _RAND_203 = {1{`RANDOM}};
  rob_payload_66_tsc = _RAND_203[31:0];
  _RAND_204 = {1{`RANDOM}};
  rob_payload_66_rob_idx = _RAND_204[15:0];
  _RAND_205 = {1{`RANDOM}};
  rob_payload_66_flits_fired = _RAND_205[15:0];
  _RAND_206 = {1{`RANDOM}};
  rob_payload_67_tsc = _RAND_206[31:0];
  _RAND_207 = {1{`RANDOM}};
  rob_payload_67_rob_idx = _RAND_207[15:0];
  _RAND_208 = {1{`RANDOM}};
  rob_payload_67_flits_fired = _RAND_208[15:0];
  _RAND_209 = {1{`RANDOM}};
  rob_payload_68_tsc = _RAND_209[31:0];
  _RAND_210 = {1{`RANDOM}};
  rob_payload_68_rob_idx = _RAND_210[15:0];
  _RAND_211 = {1{`RANDOM}};
  rob_payload_68_flits_fired = _RAND_211[15:0];
  _RAND_212 = {1{`RANDOM}};
  rob_payload_69_tsc = _RAND_212[31:0];
  _RAND_213 = {1{`RANDOM}};
  rob_payload_69_rob_idx = _RAND_213[15:0];
  _RAND_214 = {1{`RANDOM}};
  rob_payload_69_flits_fired = _RAND_214[15:0];
  _RAND_215 = {1{`RANDOM}};
  rob_payload_70_tsc = _RAND_215[31:0];
  _RAND_216 = {1{`RANDOM}};
  rob_payload_70_rob_idx = _RAND_216[15:0];
  _RAND_217 = {1{`RANDOM}};
  rob_payload_70_flits_fired = _RAND_217[15:0];
  _RAND_218 = {1{`RANDOM}};
  rob_payload_71_tsc = _RAND_218[31:0];
  _RAND_219 = {1{`RANDOM}};
  rob_payload_71_rob_idx = _RAND_219[15:0];
  _RAND_220 = {1{`RANDOM}};
  rob_payload_71_flits_fired = _RAND_220[15:0];
  _RAND_221 = {1{`RANDOM}};
  rob_payload_72_tsc = _RAND_221[31:0];
  _RAND_222 = {1{`RANDOM}};
  rob_payload_72_rob_idx = _RAND_222[15:0];
  _RAND_223 = {1{`RANDOM}};
  rob_payload_72_flits_fired = _RAND_223[15:0];
  _RAND_224 = {1{`RANDOM}};
  rob_payload_73_tsc = _RAND_224[31:0];
  _RAND_225 = {1{`RANDOM}};
  rob_payload_73_rob_idx = _RAND_225[15:0];
  _RAND_226 = {1{`RANDOM}};
  rob_payload_73_flits_fired = _RAND_226[15:0];
  _RAND_227 = {1{`RANDOM}};
  rob_payload_74_tsc = _RAND_227[31:0];
  _RAND_228 = {1{`RANDOM}};
  rob_payload_74_rob_idx = _RAND_228[15:0];
  _RAND_229 = {1{`RANDOM}};
  rob_payload_74_flits_fired = _RAND_229[15:0];
  _RAND_230 = {1{`RANDOM}};
  rob_payload_75_tsc = _RAND_230[31:0];
  _RAND_231 = {1{`RANDOM}};
  rob_payload_75_rob_idx = _RAND_231[15:0];
  _RAND_232 = {1{`RANDOM}};
  rob_payload_75_flits_fired = _RAND_232[15:0];
  _RAND_233 = {1{`RANDOM}};
  rob_payload_76_tsc = _RAND_233[31:0];
  _RAND_234 = {1{`RANDOM}};
  rob_payload_76_rob_idx = _RAND_234[15:0];
  _RAND_235 = {1{`RANDOM}};
  rob_payload_76_flits_fired = _RAND_235[15:0];
  _RAND_236 = {1{`RANDOM}};
  rob_payload_77_tsc = _RAND_236[31:0];
  _RAND_237 = {1{`RANDOM}};
  rob_payload_77_rob_idx = _RAND_237[15:0];
  _RAND_238 = {1{`RANDOM}};
  rob_payload_77_flits_fired = _RAND_238[15:0];
  _RAND_239 = {1{`RANDOM}};
  rob_payload_78_tsc = _RAND_239[31:0];
  _RAND_240 = {1{`RANDOM}};
  rob_payload_78_rob_idx = _RAND_240[15:0];
  _RAND_241 = {1{`RANDOM}};
  rob_payload_78_flits_fired = _RAND_241[15:0];
  _RAND_242 = {1{`RANDOM}};
  rob_payload_79_tsc = _RAND_242[31:0];
  _RAND_243 = {1{`RANDOM}};
  rob_payload_79_rob_idx = _RAND_243[15:0];
  _RAND_244 = {1{`RANDOM}};
  rob_payload_79_flits_fired = _RAND_244[15:0];
  _RAND_245 = {1{`RANDOM}};
  rob_payload_80_tsc = _RAND_245[31:0];
  _RAND_246 = {1{`RANDOM}};
  rob_payload_80_rob_idx = _RAND_246[15:0];
  _RAND_247 = {1{`RANDOM}};
  rob_payload_80_flits_fired = _RAND_247[15:0];
  _RAND_248 = {1{`RANDOM}};
  rob_payload_81_tsc = _RAND_248[31:0];
  _RAND_249 = {1{`RANDOM}};
  rob_payload_81_rob_idx = _RAND_249[15:0];
  _RAND_250 = {1{`RANDOM}};
  rob_payload_81_flits_fired = _RAND_250[15:0];
  _RAND_251 = {1{`RANDOM}};
  rob_payload_82_tsc = _RAND_251[31:0];
  _RAND_252 = {1{`RANDOM}};
  rob_payload_82_rob_idx = _RAND_252[15:0];
  _RAND_253 = {1{`RANDOM}};
  rob_payload_82_flits_fired = _RAND_253[15:0];
  _RAND_254 = {1{`RANDOM}};
  rob_payload_83_tsc = _RAND_254[31:0];
  _RAND_255 = {1{`RANDOM}};
  rob_payload_83_rob_idx = _RAND_255[15:0];
  _RAND_256 = {1{`RANDOM}};
  rob_payload_83_flits_fired = _RAND_256[15:0];
  _RAND_257 = {1{`RANDOM}};
  rob_payload_84_tsc = _RAND_257[31:0];
  _RAND_258 = {1{`RANDOM}};
  rob_payload_84_rob_idx = _RAND_258[15:0];
  _RAND_259 = {1{`RANDOM}};
  rob_payload_84_flits_fired = _RAND_259[15:0];
  _RAND_260 = {1{`RANDOM}};
  rob_payload_85_tsc = _RAND_260[31:0];
  _RAND_261 = {1{`RANDOM}};
  rob_payload_85_rob_idx = _RAND_261[15:0];
  _RAND_262 = {1{`RANDOM}};
  rob_payload_85_flits_fired = _RAND_262[15:0];
  _RAND_263 = {1{`RANDOM}};
  rob_payload_86_tsc = _RAND_263[31:0];
  _RAND_264 = {1{`RANDOM}};
  rob_payload_86_rob_idx = _RAND_264[15:0];
  _RAND_265 = {1{`RANDOM}};
  rob_payload_86_flits_fired = _RAND_265[15:0];
  _RAND_266 = {1{`RANDOM}};
  rob_payload_87_tsc = _RAND_266[31:0];
  _RAND_267 = {1{`RANDOM}};
  rob_payload_87_rob_idx = _RAND_267[15:0];
  _RAND_268 = {1{`RANDOM}};
  rob_payload_87_flits_fired = _RAND_268[15:0];
  _RAND_269 = {1{`RANDOM}};
  rob_payload_88_tsc = _RAND_269[31:0];
  _RAND_270 = {1{`RANDOM}};
  rob_payload_88_rob_idx = _RAND_270[15:0];
  _RAND_271 = {1{`RANDOM}};
  rob_payload_88_flits_fired = _RAND_271[15:0];
  _RAND_272 = {1{`RANDOM}};
  rob_payload_89_tsc = _RAND_272[31:0];
  _RAND_273 = {1{`RANDOM}};
  rob_payload_89_rob_idx = _RAND_273[15:0];
  _RAND_274 = {1{`RANDOM}};
  rob_payload_89_flits_fired = _RAND_274[15:0];
  _RAND_275 = {1{`RANDOM}};
  rob_payload_90_tsc = _RAND_275[31:0];
  _RAND_276 = {1{`RANDOM}};
  rob_payload_90_rob_idx = _RAND_276[15:0];
  _RAND_277 = {1{`RANDOM}};
  rob_payload_90_flits_fired = _RAND_277[15:0];
  _RAND_278 = {1{`RANDOM}};
  rob_payload_91_tsc = _RAND_278[31:0];
  _RAND_279 = {1{`RANDOM}};
  rob_payload_91_rob_idx = _RAND_279[15:0];
  _RAND_280 = {1{`RANDOM}};
  rob_payload_91_flits_fired = _RAND_280[15:0];
  _RAND_281 = {1{`RANDOM}};
  rob_payload_92_tsc = _RAND_281[31:0];
  _RAND_282 = {1{`RANDOM}};
  rob_payload_92_rob_idx = _RAND_282[15:0];
  _RAND_283 = {1{`RANDOM}};
  rob_payload_92_flits_fired = _RAND_283[15:0];
  _RAND_284 = {1{`RANDOM}};
  rob_payload_93_tsc = _RAND_284[31:0];
  _RAND_285 = {1{`RANDOM}};
  rob_payload_93_rob_idx = _RAND_285[15:0];
  _RAND_286 = {1{`RANDOM}};
  rob_payload_93_flits_fired = _RAND_286[15:0];
  _RAND_287 = {1{`RANDOM}};
  rob_payload_94_tsc = _RAND_287[31:0];
  _RAND_288 = {1{`RANDOM}};
  rob_payload_94_rob_idx = _RAND_288[15:0];
  _RAND_289 = {1{`RANDOM}};
  rob_payload_94_flits_fired = _RAND_289[15:0];
  _RAND_290 = {1{`RANDOM}};
  rob_payload_95_tsc = _RAND_290[31:0];
  _RAND_291 = {1{`RANDOM}};
  rob_payload_95_rob_idx = _RAND_291[15:0];
  _RAND_292 = {1{`RANDOM}};
  rob_payload_95_flits_fired = _RAND_292[15:0];
  _RAND_293 = {1{`RANDOM}};
  rob_payload_96_tsc = _RAND_293[31:0];
  _RAND_294 = {1{`RANDOM}};
  rob_payload_96_rob_idx = _RAND_294[15:0];
  _RAND_295 = {1{`RANDOM}};
  rob_payload_96_flits_fired = _RAND_295[15:0];
  _RAND_296 = {1{`RANDOM}};
  rob_payload_97_tsc = _RAND_296[31:0];
  _RAND_297 = {1{`RANDOM}};
  rob_payload_97_rob_idx = _RAND_297[15:0];
  _RAND_298 = {1{`RANDOM}};
  rob_payload_97_flits_fired = _RAND_298[15:0];
  _RAND_299 = {1{`RANDOM}};
  rob_payload_98_tsc = _RAND_299[31:0];
  _RAND_300 = {1{`RANDOM}};
  rob_payload_98_rob_idx = _RAND_300[15:0];
  _RAND_301 = {1{`RANDOM}};
  rob_payload_98_flits_fired = _RAND_301[15:0];
  _RAND_302 = {1{`RANDOM}};
  rob_payload_99_tsc = _RAND_302[31:0];
  _RAND_303 = {1{`RANDOM}};
  rob_payload_99_rob_idx = _RAND_303[15:0];
  _RAND_304 = {1{`RANDOM}};
  rob_payload_99_flits_fired = _RAND_304[15:0];
  _RAND_305 = {1{`RANDOM}};
  rob_payload_100_tsc = _RAND_305[31:0];
  _RAND_306 = {1{`RANDOM}};
  rob_payload_100_rob_idx = _RAND_306[15:0];
  _RAND_307 = {1{`RANDOM}};
  rob_payload_100_flits_fired = _RAND_307[15:0];
  _RAND_308 = {1{`RANDOM}};
  rob_payload_101_tsc = _RAND_308[31:0];
  _RAND_309 = {1{`RANDOM}};
  rob_payload_101_rob_idx = _RAND_309[15:0];
  _RAND_310 = {1{`RANDOM}};
  rob_payload_101_flits_fired = _RAND_310[15:0];
  _RAND_311 = {1{`RANDOM}};
  rob_payload_102_tsc = _RAND_311[31:0];
  _RAND_312 = {1{`RANDOM}};
  rob_payload_102_rob_idx = _RAND_312[15:0];
  _RAND_313 = {1{`RANDOM}};
  rob_payload_102_flits_fired = _RAND_313[15:0];
  _RAND_314 = {1{`RANDOM}};
  rob_payload_103_tsc = _RAND_314[31:0];
  _RAND_315 = {1{`RANDOM}};
  rob_payload_103_rob_idx = _RAND_315[15:0];
  _RAND_316 = {1{`RANDOM}};
  rob_payload_103_flits_fired = _RAND_316[15:0];
  _RAND_317 = {1{`RANDOM}};
  rob_payload_104_tsc = _RAND_317[31:0];
  _RAND_318 = {1{`RANDOM}};
  rob_payload_104_rob_idx = _RAND_318[15:0];
  _RAND_319 = {1{`RANDOM}};
  rob_payload_104_flits_fired = _RAND_319[15:0];
  _RAND_320 = {1{`RANDOM}};
  rob_payload_105_tsc = _RAND_320[31:0];
  _RAND_321 = {1{`RANDOM}};
  rob_payload_105_rob_idx = _RAND_321[15:0];
  _RAND_322 = {1{`RANDOM}};
  rob_payload_105_flits_fired = _RAND_322[15:0];
  _RAND_323 = {1{`RANDOM}};
  rob_payload_106_tsc = _RAND_323[31:0];
  _RAND_324 = {1{`RANDOM}};
  rob_payload_106_rob_idx = _RAND_324[15:0];
  _RAND_325 = {1{`RANDOM}};
  rob_payload_106_flits_fired = _RAND_325[15:0];
  _RAND_326 = {1{`RANDOM}};
  rob_payload_107_tsc = _RAND_326[31:0];
  _RAND_327 = {1{`RANDOM}};
  rob_payload_107_rob_idx = _RAND_327[15:0];
  _RAND_328 = {1{`RANDOM}};
  rob_payload_107_flits_fired = _RAND_328[15:0];
  _RAND_329 = {1{`RANDOM}};
  rob_payload_108_tsc = _RAND_329[31:0];
  _RAND_330 = {1{`RANDOM}};
  rob_payload_108_rob_idx = _RAND_330[15:0];
  _RAND_331 = {1{`RANDOM}};
  rob_payload_108_flits_fired = _RAND_331[15:0];
  _RAND_332 = {1{`RANDOM}};
  rob_payload_109_tsc = _RAND_332[31:0];
  _RAND_333 = {1{`RANDOM}};
  rob_payload_109_rob_idx = _RAND_333[15:0];
  _RAND_334 = {1{`RANDOM}};
  rob_payload_109_flits_fired = _RAND_334[15:0];
  _RAND_335 = {1{`RANDOM}};
  rob_payload_110_tsc = _RAND_335[31:0];
  _RAND_336 = {1{`RANDOM}};
  rob_payload_110_rob_idx = _RAND_336[15:0];
  _RAND_337 = {1{`RANDOM}};
  rob_payload_110_flits_fired = _RAND_337[15:0];
  _RAND_338 = {1{`RANDOM}};
  rob_payload_111_tsc = _RAND_338[31:0];
  _RAND_339 = {1{`RANDOM}};
  rob_payload_111_rob_idx = _RAND_339[15:0];
  _RAND_340 = {1{`RANDOM}};
  rob_payload_111_flits_fired = _RAND_340[15:0];
  _RAND_341 = {1{`RANDOM}};
  rob_payload_112_tsc = _RAND_341[31:0];
  _RAND_342 = {1{`RANDOM}};
  rob_payload_112_rob_idx = _RAND_342[15:0];
  _RAND_343 = {1{`RANDOM}};
  rob_payload_112_flits_fired = _RAND_343[15:0];
  _RAND_344 = {1{`RANDOM}};
  rob_payload_113_tsc = _RAND_344[31:0];
  _RAND_345 = {1{`RANDOM}};
  rob_payload_113_rob_idx = _RAND_345[15:0];
  _RAND_346 = {1{`RANDOM}};
  rob_payload_113_flits_fired = _RAND_346[15:0];
  _RAND_347 = {1{`RANDOM}};
  rob_payload_114_tsc = _RAND_347[31:0];
  _RAND_348 = {1{`RANDOM}};
  rob_payload_114_rob_idx = _RAND_348[15:0];
  _RAND_349 = {1{`RANDOM}};
  rob_payload_114_flits_fired = _RAND_349[15:0];
  _RAND_350 = {1{`RANDOM}};
  rob_payload_115_tsc = _RAND_350[31:0];
  _RAND_351 = {1{`RANDOM}};
  rob_payload_115_rob_idx = _RAND_351[15:0];
  _RAND_352 = {1{`RANDOM}};
  rob_payload_115_flits_fired = _RAND_352[15:0];
  _RAND_353 = {1{`RANDOM}};
  rob_payload_116_tsc = _RAND_353[31:0];
  _RAND_354 = {1{`RANDOM}};
  rob_payload_116_rob_idx = _RAND_354[15:0];
  _RAND_355 = {1{`RANDOM}};
  rob_payload_116_flits_fired = _RAND_355[15:0];
  _RAND_356 = {1{`RANDOM}};
  rob_payload_117_tsc = _RAND_356[31:0];
  _RAND_357 = {1{`RANDOM}};
  rob_payload_117_rob_idx = _RAND_357[15:0];
  _RAND_358 = {1{`RANDOM}};
  rob_payload_117_flits_fired = _RAND_358[15:0];
  _RAND_359 = {1{`RANDOM}};
  rob_payload_118_tsc = _RAND_359[31:0];
  _RAND_360 = {1{`RANDOM}};
  rob_payload_118_rob_idx = _RAND_360[15:0];
  _RAND_361 = {1{`RANDOM}};
  rob_payload_118_flits_fired = _RAND_361[15:0];
  _RAND_362 = {1{`RANDOM}};
  rob_payload_119_tsc = _RAND_362[31:0];
  _RAND_363 = {1{`RANDOM}};
  rob_payload_119_rob_idx = _RAND_363[15:0];
  _RAND_364 = {1{`RANDOM}};
  rob_payload_119_flits_fired = _RAND_364[15:0];
  _RAND_365 = {1{`RANDOM}};
  rob_payload_120_tsc = _RAND_365[31:0];
  _RAND_366 = {1{`RANDOM}};
  rob_payload_120_rob_idx = _RAND_366[15:0];
  _RAND_367 = {1{`RANDOM}};
  rob_payload_120_flits_fired = _RAND_367[15:0];
  _RAND_368 = {1{`RANDOM}};
  rob_payload_121_tsc = _RAND_368[31:0];
  _RAND_369 = {1{`RANDOM}};
  rob_payload_121_rob_idx = _RAND_369[15:0];
  _RAND_370 = {1{`RANDOM}};
  rob_payload_121_flits_fired = _RAND_370[15:0];
  _RAND_371 = {1{`RANDOM}};
  rob_payload_122_tsc = _RAND_371[31:0];
  _RAND_372 = {1{`RANDOM}};
  rob_payload_122_rob_idx = _RAND_372[15:0];
  _RAND_373 = {1{`RANDOM}};
  rob_payload_122_flits_fired = _RAND_373[15:0];
  _RAND_374 = {1{`RANDOM}};
  rob_payload_123_tsc = _RAND_374[31:0];
  _RAND_375 = {1{`RANDOM}};
  rob_payload_123_rob_idx = _RAND_375[15:0];
  _RAND_376 = {1{`RANDOM}};
  rob_payload_123_flits_fired = _RAND_376[15:0];
  _RAND_377 = {1{`RANDOM}};
  rob_payload_124_tsc = _RAND_377[31:0];
  _RAND_378 = {1{`RANDOM}};
  rob_payload_124_rob_idx = _RAND_378[15:0];
  _RAND_379 = {1{`RANDOM}};
  rob_payload_124_flits_fired = _RAND_379[15:0];
  _RAND_380 = {1{`RANDOM}};
  rob_payload_125_tsc = _RAND_380[31:0];
  _RAND_381 = {1{`RANDOM}};
  rob_payload_125_rob_idx = _RAND_381[15:0];
  _RAND_382 = {1{`RANDOM}};
  rob_payload_125_flits_fired = _RAND_382[15:0];
  _RAND_383 = {1{`RANDOM}};
  rob_payload_126_tsc = _RAND_383[31:0];
  _RAND_384 = {1{`RANDOM}};
  rob_payload_126_rob_idx = _RAND_384[15:0];
  _RAND_385 = {1{`RANDOM}};
  rob_payload_126_flits_fired = _RAND_385[15:0];
  _RAND_386 = {1{`RANDOM}};
  rob_payload_127_tsc = _RAND_386[31:0];
  _RAND_387 = {1{`RANDOM}};
  rob_payload_127_rob_idx = _RAND_387[15:0];
  _RAND_388 = {1{`RANDOM}};
  rob_payload_127_flits_fired = _RAND_388[15:0];
  _RAND_389 = {1{`RANDOM}};
  rob_n_flits_0 = _RAND_389[3:0];
  _RAND_390 = {1{`RANDOM}};
  rob_n_flits_1 = _RAND_390[3:0];
  _RAND_391 = {1{`RANDOM}};
  rob_n_flits_2 = _RAND_391[3:0];
  _RAND_392 = {1{`RANDOM}};
  rob_n_flits_3 = _RAND_392[3:0];
  _RAND_393 = {1{`RANDOM}};
  rob_n_flits_4 = _RAND_393[3:0];
  _RAND_394 = {1{`RANDOM}};
  rob_n_flits_5 = _RAND_394[3:0];
  _RAND_395 = {1{`RANDOM}};
  rob_n_flits_6 = _RAND_395[3:0];
  _RAND_396 = {1{`RANDOM}};
  rob_n_flits_7 = _RAND_396[3:0];
  _RAND_397 = {1{`RANDOM}};
  rob_n_flits_8 = _RAND_397[3:0];
  _RAND_398 = {1{`RANDOM}};
  rob_n_flits_9 = _RAND_398[3:0];
  _RAND_399 = {1{`RANDOM}};
  rob_n_flits_10 = _RAND_399[3:0];
  _RAND_400 = {1{`RANDOM}};
  rob_n_flits_11 = _RAND_400[3:0];
  _RAND_401 = {1{`RANDOM}};
  rob_n_flits_12 = _RAND_401[3:0];
  _RAND_402 = {1{`RANDOM}};
  rob_n_flits_13 = _RAND_402[3:0];
  _RAND_403 = {1{`RANDOM}};
  rob_n_flits_14 = _RAND_403[3:0];
  _RAND_404 = {1{`RANDOM}};
  rob_n_flits_15 = _RAND_404[3:0];
  _RAND_405 = {1{`RANDOM}};
  rob_n_flits_16 = _RAND_405[3:0];
  _RAND_406 = {1{`RANDOM}};
  rob_n_flits_17 = _RAND_406[3:0];
  _RAND_407 = {1{`RANDOM}};
  rob_n_flits_18 = _RAND_407[3:0];
  _RAND_408 = {1{`RANDOM}};
  rob_n_flits_19 = _RAND_408[3:0];
  _RAND_409 = {1{`RANDOM}};
  rob_n_flits_20 = _RAND_409[3:0];
  _RAND_410 = {1{`RANDOM}};
  rob_n_flits_21 = _RAND_410[3:0];
  _RAND_411 = {1{`RANDOM}};
  rob_n_flits_22 = _RAND_411[3:0];
  _RAND_412 = {1{`RANDOM}};
  rob_n_flits_23 = _RAND_412[3:0];
  _RAND_413 = {1{`RANDOM}};
  rob_n_flits_24 = _RAND_413[3:0];
  _RAND_414 = {1{`RANDOM}};
  rob_n_flits_25 = _RAND_414[3:0];
  _RAND_415 = {1{`RANDOM}};
  rob_n_flits_26 = _RAND_415[3:0];
  _RAND_416 = {1{`RANDOM}};
  rob_n_flits_27 = _RAND_416[3:0];
  _RAND_417 = {1{`RANDOM}};
  rob_n_flits_28 = _RAND_417[3:0];
  _RAND_418 = {1{`RANDOM}};
  rob_n_flits_29 = _RAND_418[3:0];
  _RAND_419 = {1{`RANDOM}};
  rob_n_flits_30 = _RAND_419[3:0];
  _RAND_420 = {1{`RANDOM}};
  rob_n_flits_31 = _RAND_420[3:0];
  _RAND_421 = {1{`RANDOM}};
  rob_n_flits_32 = _RAND_421[3:0];
  _RAND_422 = {1{`RANDOM}};
  rob_n_flits_33 = _RAND_422[3:0];
  _RAND_423 = {1{`RANDOM}};
  rob_n_flits_34 = _RAND_423[3:0];
  _RAND_424 = {1{`RANDOM}};
  rob_n_flits_35 = _RAND_424[3:0];
  _RAND_425 = {1{`RANDOM}};
  rob_n_flits_36 = _RAND_425[3:0];
  _RAND_426 = {1{`RANDOM}};
  rob_n_flits_37 = _RAND_426[3:0];
  _RAND_427 = {1{`RANDOM}};
  rob_n_flits_38 = _RAND_427[3:0];
  _RAND_428 = {1{`RANDOM}};
  rob_n_flits_39 = _RAND_428[3:0];
  _RAND_429 = {1{`RANDOM}};
  rob_n_flits_40 = _RAND_429[3:0];
  _RAND_430 = {1{`RANDOM}};
  rob_n_flits_41 = _RAND_430[3:0];
  _RAND_431 = {1{`RANDOM}};
  rob_n_flits_42 = _RAND_431[3:0];
  _RAND_432 = {1{`RANDOM}};
  rob_n_flits_43 = _RAND_432[3:0];
  _RAND_433 = {1{`RANDOM}};
  rob_n_flits_44 = _RAND_433[3:0];
  _RAND_434 = {1{`RANDOM}};
  rob_n_flits_45 = _RAND_434[3:0];
  _RAND_435 = {1{`RANDOM}};
  rob_n_flits_46 = _RAND_435[3:0];
  _RAND_436 = {1{`RANDOM}};
  rob_n_flits_47 = _RAND_436[3:0];
  _RAND_437 = {1{`RANDOM}};
  rob_n_flits_48 = _RAND_437[3:0];
  _RAND_438 = {1{`RANDOM}};
  rob_n_flits_49 = _RAND_438[3:0];
  _RAND_439 = {1{`RANDOM}};
  rob_n_flits_50 = _RAND_439[3:0];
  _RAND_440 = {1{`RANDOM}};
  rob_n_flits_51 = _RAND_440[3:0];
  _RAND_441 = {1{`RANDOM}};
  rob_n_flits_52 = _RAND_441[3:0];
  _RAND_442 = {1{`RANDOM}};
  rob_n_flits_53 = _RAND_442[3:0];
  _RAND_443 = {1{`RANDOM}};
  rob_n_flits_54 = _RAND_443[3:0];
  _RAND_444 = {1{`RANDOM}};
  rob_n_flits_55 = _RAND_444[3:0];
  _RAND_445 = {1{`RANDOM}};
  rob_n_flits_56 = _RAND_445[3:0];
  _RAND_446 = {1{`RANDOM}};
  rob_n_flits_57 = _RAND_446[3:0];
  _RAND_447 = {1{`RANDOM}};
  rob_n_flits_58 = _RAND_447[3:0];
  _RAND_448 = {1{`RANDOM}};
  rob_n_flits_59 = _RAND_448[3:0];
  _RAND_449 = {1{`RANDOM}};
  rob_n_flits_60 = _RAND_449[3:0];
  _RAND_450 = {1{`RANDOM}};
  rob_n_flits_61 = _RAND_450[3:0];
  _RAND_451 = {1{`RANDOM}};
  rob_n_flits_62 = _RAND_451[3:0];
  _RAND_452 = {1{`RANDOM}};
  rob_n_flits_63 = _RAND_452[3:0];
  _RAND_453 = {1{`RANDOM}};
  rob_n_flits_64 = _RAND_453[3:0];
  _RAND_454 = {1{`RANDOM}};
  rob_n_flits_65 = _RAND_454[3:0];
  _RAND_455 = {1{`RANDOM}};
  rob_n_flits_66 = _RAND_455[3:0];
  _RAND_456 = {1{`RANDOM}};
  rob_n_flits_67 = _RAND_456[3:0];
  _RAND_457 = {1{`RANDOM}};
  rob_n_flits_68 = _RAND_457[3:0];
  _RAND_458 = {1{`RANDOM}};
  rob_n_flits_69 = _RAND_458[3:0];
  _RAND_459 = {1{`RANDOM}};
  rob_n_flits_70 = _RAND_459[3:0];
  _RAND_460 = {1{`RANDOM}};
  rob_n_flits_71 = _RAND_460[3:0];
  _RAND_461 = {1{`RANDOM}};
  rob_n_flits_72 = _RAND_461[3:0];
  _RAND_462 = {1{`RANDOM}};
  rob_n_flits_73 = _RAND_462[3:0];
  _RAND_463 = {1{`RANDOM}};
  rob_n_flits_74 = _RAND_463[3:0];
  _RAND_464 = {1{`RANDOM}};
  rob_n_flits_75 = _RAND_464[3:0];
  _RAND_465 = {1{`RANDOM}};
  rob_n_flits_76 = _RAND_465[3:0];
  _RAND_466 = {1{`RANDOM}};
  rob_n_flits_77 = _RAND_466[3:0];
  _RAND_467 = {1{`RANDOM}};
  rob_n_flits_78 = _RAND_467[3:0];
  _RAND_468 = {1{`RANDOM}};
  rob_n_flits_79 = _RAND_468[3:0];
  _RAND_469 = {1{`RANDOM}};
  rob_n_flits_80 = _RAND_469[3:0];
  _RAND_470 = {1{`RANDOM}};
  rob_n_flits_81 = _RAND_470[3:0];
  _RAND_471 = {1{`RANDOM}};
  rob_n_flits_82 = _RAND_471[3:0];
  _RAND_472 = {1{`RANDOM}};
  rob_n_flits_83 = _RAND_472[3:0];
  _RAND_473 = {1{`RANDOM}};
  rob_n_flits_84 = _RAND_473[3:0];
  _RAND_474 = {1{`RANDOM}};
  rob_n_flits_85 = _RAND_474[3:0];
  _RAND_475 = {1{`RANDOM}};
  rob_n_flits_86 = _RAND_475[3:0];
  _RAND_476 = {1{`RANDOM}};
  rob_n_flits_87 = _RAND_476[3:0];
  _RAND_477 = {1{`RANDOM}};
  rob_n_flits_88 = _RAND_477[3:0];
  _RAND_478 = {1{`RANDOM}};
  rob_n_flits_89 = _RAND_478[3:0];
  _RAND_479 = {1{`RANDOM}};
  rob_n_flits_90 = _RAND_479[3:0];
  _RAND_480 = {1{`RANDOM}};
  rob_n_flits_91 = _RAND_480[3:0];
  _RAND_481 = {1{`RANDOM}};
  rob_n_flits_92 = _RAND_481[3:0];
  _RAND_482 = {1{`RANDOM}};
  rob_n_flits_93 = _RAND_482[3:0];
  _RAND_483 = {1{`RANDOM}};
  rob_n_flits_94 = _RAND_483[3:0];
  _RAND_484 = {1{`RANDOM}};
  rob_n_flits_95 = _RAND_484[3:0];
  _RAND_485 = {1{`RANDOM}};
  rob_n_flits_96 = _RAND_485[3:0];
  _RAND_486 = {1{`RANDOM}};
  rob_n_flits_97 = _RAND_486[3:0];
  _RAND_487 = {1{`RANDOM}};
  rob_n_flits_98 = _RAND_487[3:0];
  _RAND_488 = {1{`RANDOM}};
  rob_n_flits_99 = _RAND_488[3:0];
  _RAND_489 = {1{`RANDOM}};
  rob_n_flits_100 = _RAND_489[3:0];
  _RAND_490 = {1{`RANDOM}};
  rob_n_flits_101 = _RAND_490[3:0];
  _RAND_491 = {1{`RANDOM}};
  rob_n_flits_102 = _RAND_491[3:0];
  _RAND_492 = {1{`RANDOM}};
  rob_n_flits_103 = _RAND_492[3:0];
  _RAND_493 = {1{`RANDOM}};
  rob_n_flits_104 = _RAND_493[3:0];
  _RAND_494 = {1{`RANDOM}};
  rob_n_flits_105 = _RAND_494[3:0];
  _RAND_495 = {1{`RANDOM}};
  rob_n_flits_106 = _RAND_495[3:0];
  _RAND_496 = {1{`RANDOM}};
  rob_n_flits_107 = _RAND_496[3:0];
  _RAND_497 = {1{`RANDOM}};
  rob_n_flits_108 = _RAND_497[3:0];
  _RAND_498 = {1{`RANDOM}};
  rob_n_flits_109 = _RAND_498[3:0];
  _RAND_499 = {1{`RANDOM}};
  rob_n_flits_110 = _RAND_499[3:0];
  _RAND_500 = {1{`RANDOM}};
  rob_n_flits_111 = _RAND_500[3:0];
  _RAND_501 = {1{`RANDOM}};
  rob_n_flits_112 = _RAND_501[3:0];
  _RAND_502 = {1{`RANDOM}};
  rob_n_flits_113 = _RAND_502[3:0];
  _RAND_503 = {1{`RANDOM}};
  rob_n_flits_114 = _RAND_503[3:0];
  _RAND_504 = {1{`RANDOM}};
  rob_n_flits_115 = _RAND_504[3:0];
  _RAND_505 = {1{`RANDOM}};
  rob_n_flits_116 = _RAND_505[3:0];
  _RAND_506 = {1{`RANDOM}};
  rob_n_flits_117 = _RAND_506[3:0];
  _RAND_507 = {1{`RANDOM}};
  rob_n_flits_118 = _RAND_507[3:0];
  _RAND_508 = {1{`RANDOM}};
  rob_n_flits_119 = _RAND_508[3:0];
  _RAND_509 = {1{`RANDOM}};
  rob_n_flits_120 = _RAND_509[3:0];
  _RAND_510 = {1{`RANDOM}};
  rob_n_flits_121 = _RAND_510[3:0];
  _RAND_511 = {1{`RANDOM}};
  rob_n_flits_122 = _RAND_511[3:0];
  _RAND_512 = {1{`RANDOM}};
  rob_n_flits_123 = _RAND_512[3:0];
  _RAND_513 = {1{`RANDOM}};
  rob_n_flits_124 = _RAND_513[3:0];
  _RAND_514 = {1{`RANDOM}};
  rob_n_flits_125 = _RAND_514[3:0];
  _RAND_515 = {1{`RANDOM}};
  rob_n_flits_126 = _RAND_515[3:0];
  _RAND_516 = {1{`RANDOM}};
  rob_n_flits_127 = _RAND_516[3:0];
  _RAND_517 = {1{`RANDOM}};
  rob_flits_returned_0 = _RAND_517[3:0];
  _RAND_518 = {1{`RANDOM}};
  rob_flits_returned_1 = _RAND_518[3:0];
  _RAND_519 = {1{`RANDOM}};
  rob_flits_returned_2 = _RAND_519[3:0];
  _RAND_520 = {1{`RANDOM}};
  rob_flits_returned_3 = _RAND_520[3:0];
  _RAND_521 = {1{`RANDOM}};
  rob_flits_returned_4 = _RAND_521[3:0];
  _RAND_522 = {1{`RANDOM}};
  rob_flits_returned_5 = _RAND_522[3:0];
  _RAND_523 = {1{`RANDOM}};
  rob_flits_returned_6 = _RAND_523[3:0];
  _RAND_524 = {1{`RANDOM}};
  rob_flits_returned_7 = _RAND_524[3:0];
  _RAND_525 = {1{`RANDOM}};
  rob_flits_returned_8 = _RAND_525[3:0];
  _RAND_526 = {1{`RANDOM}};
  rob_flits_returned_9 = _RAND_526[3:0];
  _RAND_527 = {1{`RANDOM}};
  rob_flits_returned_10 = _RAND_527[3:0];
  _RAND_528 = {1{`RANDOM}};
  rob_flits_returned_11 = _RAND_528[3:0];
  _RAND_529 = {1{`RANDOM}};
  rob_flits_returned_12 = _RAND_529[3:0];
  _RAND_530 = {1{`RANDOM}};
  rob_flits_returned_13 = _RAND_530[3:0];
  _RAND_531 = {1{`RANDOM}};
  rob_flits_returned_14 = _RAND_531[3:0];
  _RAND_532 = {1{`RANDOM}};
  rob_flits_returned_15 = _RAND_532[3:0];
  _RAND_533 = {1{`RANDOM}};
  rob_flits_returned_16 = _RAND_533[3:0];
  _RAND_534 = {1{`RANDOM}};
  rob_flits_returned_17 = _RAND_534[3:0];
  _RAND_535 = {1{`RANDOM}};
  rob_flits_returned_18 = _RAND_535[3:0];
  _RAND_536 = {1{`RANDOM}};
  rob_flits_returned_19 = _RAND_536[3:0];
  _RAND_537 = {1{`RANDOM}};
  rob_flits_returned_20 = _RAND_537[3:0];
  _RAND_538 = {1{`RANDOM}};
  rob_flits_returned_21 = _RAND_538[3:0];
  _RAND_539 = {1{`RANDOM}};
  rob_flits_returned_22 = _RAND_539[3:0];
  _RAND_540 = {1{`RANDOM}};
  rob_flits_returned_23 = _RAND_540[3:0];
  _RAND_541 = {1{`RANDOM}};
  rob_flits_returned_24 = _RAND_541[3:0];
  _RAND_542 = {1{`RANDOM}};
  rob_flits_returned_25 = _RAND_542[3:0];
  _RAND_543 = {1{`RANDOM}};
  rob_flits_returned_26 = _RAND_543[3:0];
  _RAND_544 = {1{`RANDOM}};
  rob_flits_returned_27 = _RAND_544[3:0];
  _RAND_545 = {1{`RANDOM}};
  rob_flits_returned_28 = _RAND_545[3:0];
  _RAND_546 = {1{`RANDOM}};
  rob_flits_returned_29 = _RAND_546[3:0];
  _RAND_547 = {1{`RANDOM}};
  rob_flits_returned_30 = _RAND_547[3:0];
  _RAND_548 = {1{`RANDOM}};
  rob_flits_returned_31 = _RAND_548[3:0];
  _RAND_549 = {1{`RANDOM}};
  rob_flits_returned_32 = _RAND_549[3:0];
  _RAND_550 = {1{`RANDOM}};
  rob_flits_returned_33 = _RAND_550[3:0];
  _RAND_551 = {1{`RANDOM}};
  rob_flits_returned_34 = _RAND_551[3:0];
  _RAND_552 = {1{`RANDOM}};
  rob_flits_returned_35 = _RAND_552[3:0];
  _RAND_553 = {1{`RANDOM}};
  rob_flits_returned_36 = _RAND_553[3:0];
  _RAND_554 = {1{`RANDOM}};
  rob_flits_returned_37 = _RAND_554[3:0];
  _RAND_555 = {1{`RANDOM}};
  rob_flits_returned_38 = _RAND_555[3:0];
  _RAND_556 = {1{`RANDOM}};
  rob_flits_returned_39 = _RAND_556[3:0];
  _RAND_557 = {1{`RANDOM}};
  rob_flits_returned_40 = _RAND_557[3:0];
  _RAND_558 = {1{`RANDOM}};
  rob_flits_returned_41 = _RAND_558[3:0];
  _RAND_559 = {1{`RANDOM}};
  rob_flits_returned_42 = _RAND_559[3:0];
  _RAND_560 = {1{`RANDOM}};
  rob_flits_returned_43 = _RAND_560[3:0];
  _RAND_561 = {1{`RANDOM}};
  rob_flits_returned_44 = _RAND_561[3:0];
  _RAND_562 = {1{`RANDOM}};
  rob_flits_returned_45 = _RAND_562[3:0];
  _RAND_563 = {1{`RANDOM}};
  rob_flits_returned_46 = _RAND_563[3:0];
  _RAND_564 = {1{`RANDOM}};
  rob_flits_returned_47 = _RAND_564[3:0];
  _RAND_565 = {1{`RANDOM}};
  rob_flits_returned_48 = _RAND_565[3:0];
  _RAND_566 = {1{`RANDOM}};
  rob_flits_returned_49 = _RAND_566[3:0];
  _RAND_567 = {1{`RANDOM}};
  rob_flits_returned_50 = _RAND_567[3:0];
  _RAND_568 = {1{`RANDOM}};
  rob_flits_returned_51 = _RAND_568[3:0];
  _RAND_569 = {1{`RANDOM}};
  rob_flits_returned_52 = _RAND_569[3:0];
  _RAND_570 = {1{`RANDOM}};
  rob_flits_returned_53 = _RAND_570[3:0];
  _RAND_571 = {1{`RANDOM}};
  rob_flits_returned_54 = _RAND_571[3:0];
  _RAND_572 = {1{`RANDOM}};
  rob_flits_returned_55 = _RAND_572[3:0];
  _RAND_573 = {1{`RANDOM}};
  rob_flits_returned_56 = _RAND_573[3:0];
  _RAND_574 = {1{`RANDOM}};
  rob_flits_returned_57 = _RAND_574[3:0];
  _RAND_575 = {1{`RANDOM}};
  rob_flits_returned_58 = _RAND_575[3:0];
  _RAND_576 = {1{`RANDOM}};
  rob_flits_returned_59 = _RAND_576[3:0];
  _RAND_577 = {1{`RANDOM}};
  rob_flits_returned_60 = _RAND_577[3:0];
  _RAND_578 = {1{`RANDOM}};
  rob_flits_returned_61 = _RAND_578[3:0];
  _RAND_579 = {1{`RANDOM}};
  rob_flits_returned_62 = _RAND_579[3:0];
  _RAND_580 = {1{`RANDOM}};
  rob_flits_returned_63 = _RAND_580[3:0];
  _RAND_581 = {1{`RANDOM}};
  rob_flits_returned_64 = _RAND_581[3:0];
  _RAND_582 = {1{`RANDOM}};
  rob_flits_returned_65 = _RAND_582[3:0];
  _RAND_583 = {1{`RANDOM}};
  rob_flits_returned_66 = _RAND_583[3:0];
  _RAND_584 = {1{`RANDOM}};
  rob_flits_returned_67 = _RAND_584[3:0];
  _RAND_585 = {1{`RANDOM}};
  rob_flits_returned_68 = _RAND_585[3:0];
  _RAND_586 = {1{`RANDOM}};
  rob_flits_returned_69 = _RAND_586[3:0];
  _RAND_587 = {1{`RANDOM}};
  rob_flits_returned_70 = _RAND_587[3:0];
  _RAND_588 = {1{`RANDOM}};
  rob_flits_returned_71 = _RAND_588[3:0];
  _RAND_589 = {1{`RANDOM}};
  rob_flits_returned_72 = _RAND_589[3:0];
  _RAND_590 = {1{`RANDOM}};
  rob_flits_returned_73 = _RAND_590[3:0];
  _RAND_591 = {1{`RANDOM}};
  rob_flits_returned_74 = _RAND_591[3:0];
  _RAND_592 = {1{`RANDOM}};
  rob_flits_returned_75 = _RAND_592[3:0];
  _RAND_593 = {1{`RANDOM}};
  rob_flits_returned_76 = _RAND_593[3:0];
  _RAND_594 = {1{`RANDOM}};
  rob_flits_returned_77 = _RAND_594[3:0];
  _RAND_595 = {1{`RANDOM}};
  rob_flits_returned_78 = _RAND_595[3:0];
  _RAND_596 = {1{`RANDOM}};
  rob_flits_returned_79 = _RAND_596[3:0];
  _RAND_597 = {1{`RANDOM}};
  rob_flits_returned_80 = _RAND_597[3:0];
  _RAND_598 = {1{`RANDOM}};
  rob_flits_returned_81 = _RAND_598[3:0];
  _RAND_599 = {1{`RANDOM}};
  rob_flits_returned_82 = _RAND_599[3:0];
  _RAND_600 = {1{`RANDOM}};
  rob_flits_returned_83 = _RAND_600[3:0];
  _RAND_601 = {1{`RANDOM}};
  rob_flits_returned_84 = _RAND_601[3:0];
  _RAND_602 = {1{`RANDOM}};
  rob_flits_returned_85 = _RAND_602[3:0];
  _RAND_603 = {1{`RANDOM}};
  rob_flits_returned_86 = _RAND_603[3:0];
  _RAND_604 = {1{`RANDOM}};
  rob_flits_returned_87 = _RAND_604[3:0];
  _RAND_605 = {1{`RANDOM}};
  rob_flits_returned_88 = _RAND_605[3:0];
  _RAND_606 = {1{`RANDOM}};
  rob_flits_returned_89 = _RAND_606[3:0];
  _RAND_607 = {1{`RANDOM}};
  rob_flits_returned_90 = _RAND_607[3:0];
  _RAND_608 = {1{`RANDOM}};
  rob_flits_returned_91 = _RAND_608[3:0];
  _RAND_609 = {1{`RANDOM}};
  rob_flits_returned_92 = _RAND_609[3:0];
  _RAND_610 = {1{`RANDOM}};
  rob_flits_returned_93 = _RAND_610[3:0];
  _RAND_611 = {1{`RANDOM}};
  rob_flits_returned_94 = _RAND_611[3:0];
  _RAND_612 = {1{`RANDOM}};
  rob_flits_returned_95 = _RAND_612[3:0];
  _RAND_613 = {1{`RANDOM}};
  rob_flits_returned_96 = _RAND_613[3:0];
  _RAND_614 = {1{`RANDOM}};
  rob_flits_returned_97 = _RAND_614[3:0];
  _RAND_615 = {1{`RANDOM}};
  rob_flits_returned_98 = _RAND_615[3:0];
  _RAND_616 = {1{`RANDOM}};
  rob_flits_returned_99 = _RAND_616[3:0];
  _RAND_617 = {1{`RANDOM}};
  rob_flits_returned_100 = _RAND_617[3:0];
  _RAND_618 = {1{`RANDOM}};
  rob_flits_returned_101 = _RAND_618[3:0];
  _RAND_619 = {1{`RANDOM}};
  rob_flits_returned_102 = _RAND_619[3:0];
  _RAND_620 = {1{`RANDOM}};
  rob_flits_returned_103 = _RAND_620[3:0];
  _RAND_621 = {1{`RANDOM}};
  rob_flits_returned_104 = _RAND_621[3:0];
  _RAND_622 = {1{`RANDOM}};
  rob_flits_returned_105 = _RAND_622[3:0];
  _RAND_623 = {1{`RANDOM}};
  rob_flits_returned_106 = _RAND_623[3:0];
  _RAND_624 = {1{`RANDOM}};
  rob_flits_returned_107 = _RAND_624[3:0];
  _RAND_625 = {1{`RANDOM}};
  rob_flits_returned_108 = _RAND_625[3:0];
  _RAND_626 = {1{`RANDOM}};
  rob_flits_returned_109 = _RAND_626[3:0];
  _RAND_627 = {1{`RANDOM}};
  rob_flits_returned_110 = _RAND_627[3:0];
  _RAND_628 = {1{`RANDOM}};
  rob_flits_returned_111 = _RAND_628[3:0];
  _RAND_629 = {1{`RANDOM}};
  rob_flits_returned_112 = _RAND_629[3:0];
  _RAND_630 = {1{`RANDOM}};
  rob_flits_returned_113 = _RAND_630[3:0];
  _RAND_631 = {1{`RANDOM}};
  rob_flits_returned_114 = _RAND_631[3:0];
  _RAND_632 = {1{`RANDOM}};
  rob_flits_returned_115 = _RAND_632[3:0];
  _RAND_633 = {1{`RANDOM}};
  rob_flits_returned_116 = _RAND_633[3:0];
  _RAND_634 = {1{`RANDOM}};
  rob_flits_returned_117 = _RAND_634[3:0];
  _RAND_635 = {1{`RANDOM}};
  rob_flits_returned_118 = _RAND_635[3:0];
  _RAND_636 = {1{`RANDOM}};
  rob_flits_returned_119 = _RAND_636[3:0];
  _RAND_637 = {1{`RANDOM}};
  rob_flits_returned_120 = _RAND_637[3:0];
  _RAND_638 = {1{`RANDOM}};
  rob_flits_returned_121 = _RAND_638[3:0];
  _RAND_639 = {1{`RANDOM}};
  rob_flits_returned_122 = _RAND_639[3:0];
  _RAND_640 = {1{`RANDOM}};
  rob_flits_returned_123 = _RAND_640[3:0];
  _RAND_641 = {1{`RANDOM}};
  rob_flits_returned_124 = _RAND_641[3:0];
  _RAND_642 = {1{`RANDOM}};
  rob_flits_returned_125 = _RAND_642[3:0];
  _RAND_643 = {1{`RANDOM}};
  rob_flits_returned_126 = _RAND_643[3:0];
  _RAND_644 = {1{`RANDOM}};
  rob_flits_returned_127 = _RAND_644[3:0];
  _RAND_645 = {2{`RANDOM}};
  rob_tscs_0 = _RAND_645[63:0];
  _RAND_646 = {2{`RANDOM}};
  rob_tscs_1 = _RAND_646[63:0];
  _RAND_647 = {2{`RANDOM}};
  rob_tscs_2 = _RAND_647[63:0];
  _RAND_648 = {2{`RANDOM}};
  rob_tscs_3 = _RAND_648[63:0];
  _RAND_649 = {2{`RANDOM}};
  rob_tscs_4 = _RAND_649[63:0];
  _RAND_650 = {2{`RANDOM}};
  rob_tscs_5 = _RAND_650[63:0];
  _RAND_651 = {2{`RANDOM}};
  rob_tscs_6 = _RAND_651[63:0];
  _RAND_652 = {2{`RANDOM}};
  rob_tscs_7 = _RAND_652[63:0];
  _RAND_653 = {2{`RANDOM}};
  rob_tscs_8 = _RAND_653[63:0];
  _RAND_654 = {2{`RANDOM}};
  rob_tscs_9 = _RAND_654[63:0];
  _RAND_655 = {2{`RANDOM}};
  rob_tscs_10 = _RAND_655[63:0];
  _RAND_656 = {2{`RANDOM}};
  rob_tscs_11 = _RAND_656[63:0];
  _RAND_657 = {2{`RANDOM}};
  rob_tscs_12 = _RAND_657[63:0];
  _RAND_658 = {2{`RANDOM}};
  rob_tscs_13 = _RAND_658[63:0];
  _RAND_659 = {2{`RANDOM}};
  rob_tscs_14 = _RAND_659[63:0];
  _RAND_660 = {2{`RANDOM}};
  rob_tscs_15 = _RAND_660[63:0];
  _RAND_661 = {2{`RANDOM}};
  rob_tscs_16 = _RAND_661[63:0];
  _RAND_662 = {2{`RANDOM}};
  rob_tscs_17 = _RAND_662[63:0];
  _RAND_663 = {2{`RANDOM}};
  rob_tscs_18 = _RAND_663[63:0];
  _RAND_664 = {2{`RANDOM}};
  rob_tscs_19 = _RAND_664[63:0];
  _RAND_665 = {2{`RANDOM}};
  rob_tscs_20 = _RAND_665[63:0];
  _RAND_666 = {2{`RANDOM}};
  rob_tscs_21 = _RAND_666[63:0];
  _RAND_667 = {2{`RANDOM}};
  rob_tscs_22 = _RAND_667[63:0];
  _RAND_668 = {2{`RANDOM}};
  rob_tscs_23 = _RAND_668[63:0];
  _RAND_669 = {2{`RANDOM}};
  rob_tscs_24 = _RAND_669[63:0];
  _RAND_670 = {2{`RANDOM}};
  rob_tscs_25 = _RAND_670[63:0];
  _RAND_671 = {2{`RANDOM}};
  rob_tscs_26 = _RAND_671[63:0];
  _RAND_672 = {2{`RANDOM}};
  rob_tscs_27 = _RAND_672[63:0];
  _RAND_673 = {2{`RANDOM}};
  rob_tscs_28 = _RAND_673[63:0];
  _RAND_674 = {2{`RANDOM}};
  rob_tscs_29 = _RAND_674[63:0];
  _RAND_675 = {2{`RANDOM}};
  rob_tscs_30 = _RAND_675[63:0];
  _RAND_676 = {2{`RANDOM}};
  rob_tscs_31 = _RAND_676[63:0];
  _RAND_677 = {2{`RANDOM}};
  rob_tscs_32 = _RAND_677[63:0];
  _RAND_678 = {2{`RANDOM}};
  rob_tscs_33 = _RAND_678[63:0];
  _RAND_679 = {2{`RANDOM}};
  rob_tscs_34 = _RAND_679[63:0];
  _RAND_680 = {2{`RANDOM}};
  rob_tscs_35 = _RAND_680[63:0];
  _RAND_681 = {2{`RANDOM}};
  rob_tscs_36 = _RAND_681[63:0];
  _RAND_682 = {2{`RANDOM}};
  rob_tscs_37 = _RAND_682[63:0];
  _RAND_683 = {2{`RANDOM}};
  rob_tscs_38 = _RAND_683[63:0];
  _RAND_684 = {2{`RANDOM}};
  rob_tscs_39 = _RAND_684[63:0];
  _RAND_685 = {2{`RANDOM}};
  rob_tscs_40 = _RAND_685[63:0];
  _RAND_686 = {2{`RANDOM}};
  rob_tscs_41 = _RAND_686[63:0];
  _RAND_687 = {2{`RANDOM}};
  rob_tscs_42 = _RAND_687[63:0];
  _RAND_688 = {2{`RANDOM}};
  rob_tscs_43 = _RAND_688[63:0];
  _RAND_689 = {2{`RANDOM}};
  rob_tscs_44 = _RAND_689[63:0];
  _RAND_690 = {2{`RANDOM}};
  rob_tscs_45 = _RAND_690[63:0];
  _RAND_691 = {2{`RANDOM}};
  rob_tscs_46 = _RAND_691[63:0];
  _RAND_692 = {2{`RANDOM}};
  rob_tscs_47 = _RAND_692[63:0];
  _RAND_693 = {2{`RANDOM}};
  rob_tscs_48 = _RAND_693[63:0];
  _RAND_694 = {2{`RANDOM}};
  rob_tscs_49 = _RAND_694[63:0];
  _RAND_695 = {2{`RANDOM}};
  rob_tscs_50 = _RAND_695[63:0];
  _RAND_696 = {2{`RANDOM}};
  rob_tscs_51 = _RAND_696[63:0];
  _RAND_697 = {2{`RANDOM}};
  rob_tscs_52 = _RAND_697[63:0];
  _RAND_698 = {2{`RANDOM}};
  rob_tscs_53 = _RAND_698[63:0];
  _RAND_699 = {2{`RANDOM}};
  rob_tscs_54 = _RAND_699[63:0];
  _RAND_700 = {2{`RANDOM}};
  rob_tscs_55 = _RAND_700[63:0];
  _RAND_701 = {2{`RANDOM}};
  rob_tscs_56 = _RAND_701[63:0];
  _RAND_702 = {2{`RANDOM}};
  rob_tscs_57 = _RAND_702[63:0];
  _RAND_703 = {2{`RANDOM}};
  rob_tscs_58 = _RAND_703[63:0];
  _RAND_704 = {2{`RANDOM}};
  rob_tscs_59 = _RAND_704[63:0];
  _RAND_705 = {2{`RANDOM}};
  rob_tscs_60 = _RAND_705[63:0];
  _RAND_706 = {2{`RANDOM}};
  rob_tscs_61 = _RAND_706[63:0];
  _RAND_707 = {2{`RANDOM}};
  rob_tscs_62 = _RAND_707[63:0];
  _RAND_708 = {2{`RANDOM}};
  rob_tscs_63 = _RAND_708[63:0];
  _RAND_709 = {2{`RANDOM}};
  rob_tscs_64 = _RAND_709[63:0];
  _RAND_710 = {2{`RANDOM}};
  rob_tscs_65 = _RAND_710[63:0];
  _RAND_711 = {2{`RANDOM}};
  rob_tscs_66 = _RAND_711[63:0];
  _RAND_712 = {2{`RANDOM}};
  rob_tscs_67 = _RAND_712[63:0];
  _RAND_713 = {2{`RANDOM}};
  rob_tscs_68 = _RAND_713[63:0];
  _RAND_714 = {2{`RANDOM}};
  rob_tscs_69 = _RAND_714[63:0];
  _RAND_715 = {2{`RANDOM}};
  rob_tscs_70 = _RAND_715[63:0];
  _RAND_716 = {2{`RANDOM}};
  rob_tscs_71 = _RAND_716[63:0];
  _RAND_717 = {2{`RANDOM}};
  rob_tscs_72 = _RAND_717[63:0];
  _RAND_718 = {2{`RANDOM}};
  rob_tscs_73 = _RAND_718[63:0];
  _RAND_719 = {2{`RANDOM}};
  rob_tscs_74 = _RAND_719[63:0];
  _RAND_720 = {2{`RANDOM}};
  rob_tscs_75 = _RAND_720[63:0];
  _RAND_721 = {2{`RANDOM}};
  rob_tscs_76 = _RAND_721[63:0];
  _RAND_722 = {2{`RANDOM}};
  rob_tscs_77 = _RAND_722[63:0];
  _RAND_723 = {2{`RANDOM}};
  rob_tscs_78 = _RAND_723[63:0];
  _RAND_724 = {2{`RANDOM}};
  rob_tscs_79 = _RAND_724[63:0];
  _RAND_725 = {2{`RANDOM}};
  rob_tscs_80 = _RAND_725[63:0];
  _RAND_726 = {2{`RANDOM}};
  rob_tscs_81 = _RAND_726[63:0];
  _RAND_727 = {2{`RANDOM}};
  rob_tscs_82 = _RAND_727[63:0];
  _RAND_728 = {2{`RANDOM}};
  rob_tscs_83 = _RAND_728[63:0];
  _RAND_729 = {2{`RANDOM}};
  rob_tscs_84 = _RAND_729[63:0];
  _RAND_730 = {2{`RANDOM}};
  rob_tscs_85 = _RAND_730[63:0];
  _RAND_731 = {2{`RANDOM}};
  rob_tscs_86 = _RAND_731[63:0];
  _RAND_732 = {2{`RANDOM}};
  rob_tscs_87 = _RAND_732[63:0];
  _RAND_733 = {2{`RANDOM}};
  rob_tscs_88 = _RAND_733[63:0];
  _RAND_734 = {2{`RANDOM}};
  rob_tscs_89 = _RAND_734[63:0];
  _RAND_735 = {2{`RANDOM}};
  rob_tscs_90 = _RAND_735[63:0];
  _RAND_736 = {2{`RANDOM}};
  rob_tscs_91 = _RAND_736[63:0];
  _RAND_737 = {2{`RANDOM}};
  rob_tscs_92 = _RAND_737[63:0];
  _RAND_738 = {2{`RANDOM}};
  rob_tscs_93 = _RAND_738[63:0];
  _RAND_739 = {2{`RANDOM}};
  rob_tscs_94 = _RAND_739[63:0];
  _RAND_740 = {2{`RANDOM}};
  rob_tscs_95 = _RAND_740[63:0];
  _RAND_741 = {2{`RANDOM}};
  rob_tscs_96 = _RAND_741[63:0];
  _RAND_742 = {2{`RANDOM}};
  rob_tscs_97 = _RAND_742[63:0];
  _RAND_743 = {2{`RANDOM}};
  rob_tscs_98 = _RAND_743[63:0];
  _RAND_744 = {2{`RANDOM}};
  rob_tscs_99 = _RAND_744[63:0];
  _RAND_745 = {2{`RANDOM}};
  rob_tscs_100 = _RAND_745[63:0];
  _RAND_746 = {2{`RANDOM}};
  rob_tscs_101 = _RAND_746[63:0];
  _RAND_747 = {2{`RANDOM}};
  rob_tscs_102 = _RAND_747[63:0];
  _RAND_748 = {2{`RANDOM}};
  rob_tscs_103 = _RAND_748[63:0];
  _RAND_749 = {2{`RANDOM}};
  rob_tscs_104 = _RAND_749[63:0];
  _RAND_750 = {2{`RANDOM}};
  rob_tscs_105 = _RAND_750[63:0];
  _RAND_751 = {2{`RANDOM}};
  rob_tscs_106 = _RAND_751[63:0];
  _RAND_752 = {2{`RANDOM}};
  rob_tscs_107 = _RAND_752[63:0];
  _RAND_753 = {2{`RANDOM}};
  rob_tscs_108 = _RAND_753[63:0];
  _RAND_754 = {2{`RANDOM}};
  rob_tscs_109 = _RAND_754[63:0];
  _RAND_755 = {2{`RANDOM}};
  rob_tscs_110 = _RAND_755[63:0];
  _RAND_756 = {2{`RANDOM}};
  rob_tscs_111 = _RAND_756[63:0];
  _RAND_757 = {2{`RANDOM}};
  rob_tscs_112 = _RAND_757[63:0];
  _RAND_758 = {2{`RANDOM}};
  rob_tscs_113 = _RAND_758[63:0];
  _RAND_759 = {2{`RANDOM}};
  rob_tscs_114 = _RAND_759[63:0];
  _RAND_760 = {2{`RANDOM}};
  rob_tscs_115 = _RAND_760[63:0];
  _RAND_761 = {2{`RANDOM}};
  rob_tscs_116 = _RAND_761[63:0];
  _RAND_762 = {2{`RANDOM}};
  rob_tscs_117 = _RAND_762[63:0];
  _RAND_763 = {2{`RANDOM}};
  rob_tscs_118 = _RAND_763[63:0];
  _RAND_764 = {2{`RANDOM}};
  rob_tscs_119 = _RAND_764[63:0];
  _RAND_765 = {2{`RANDOM}};
  rob_tscs_120 = _RAND_765[63:0];
  _RAND_766 = {2{`RANDOM}};
  rob_tscs_121 = _RAND_766[63:0];
  _RAND_767 = {2{`RANDOM}};
  rob_tscs_122 = _RAND_767[63:0];
  _RAND_768 = {2{`RANDOM}};
  rob_tscs_123 = _RAND_768[63:0];
  _RAND_769 = {2{`RANDOM}};
  rob_tscs_124 = _RAND_769[63:0];
  _RAND_770 = {2{`RANDOM}};
  rob_tscs_125 = _RAND_770[63:0];
  _RAND_771 = {2{`RANDOM}};
  rob_tscs_126 = _RAND_771[63:0];
  _RAND_772 = {2{`RANDOM}};
  rob_tscs_127 = _RAND_772[63:0];
  _RAND_773 = {1{`RANDOM}};
  io_success_REG = _RAND_773[0:0];
  _RAND_774 = {1{`RANDOM}};
  packet_valid = _RAND_774[0:0];
  _RAND_775 = {1{`RANDOM}};
  packet_rob_idx = _RAND_775[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(~idle_counter[10]); // @[TestHarness.scala 148:9]
    end
    //
    if (_T_67 & _T_3) begin
      assert(_T_25[0]); // @[TestHarness.scala 201:13]
    end
    //
    if (_T_67 & _T_3) begin
      assert(_T_31 == io_from_noc_0_flit_bits_payload); // @[TestHarness.scala 202:13]
    end
    //
    if (_T_67 & _T_3) begin
      assert(~io_from_noc_0_flit_bits_ingress_id); // @[TestHarness.scala 203:13]
    end
    //
    if (_T_67 & _T_3) begin
      assert(1'h1); // @[TestHarness.scala 204:13]
    end
    //
    if (_T_67 & _T_3) begin
      assert(_GEN_2816 < _GEN_2944); // @[TestHarness.scala 205:13]
    end
    //
    if (_T_67 & _T_3) begin
      assert(~packet_valid & io_from_noc_0_flit_bits_head | out_payload_rob_idx == _GEN_385); // @[TestHarness.scala 206:13]
    end
    //
    if (rob_valids[0] & _T_3) begin
      assert(_T_72 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[1] & _T_3) begin
      assert(_T_79 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[2] & _T_3) begin
      assert(_T_86 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[3] & _T_3) begin
      assert(_T_93 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[4] & _T_3) begin
      assert(_T_100 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[5] & _T_3) begin
      assert(_T_107 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[6] & _T_3) begin
      assert(_T_114 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[7] & _T_3) begin
      assert(_T_121 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[8] & _T_3) begin
      assert(_T_128 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[9] & _T_3) begin
      assert(_T_135 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[10] & _T_3) begin
      assert(_T_142 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[11] & _T_3) begin
      assert(_T_149 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[12] & _T_3) begin
      assert(_T_156 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[13] & _T_3) begin
      assert(_T_163 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[14] & _T_3) begin
      assert(_T_170 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[15] & _T_3) begin
      assert(_T_177 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[16] & _T_3) begin
      assert(_T_184 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[17] & _T_3) begin
      assert(_T_191 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[18] & _T_3) begin
      assert(_T_198 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[19] & _T_3) begin
      assert(_T_205 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[20] & _T_3) begin
      assert(_T_212 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[21] & _T_3) begin
      assert(_T_219 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[22] & _T_3) begin
      assert(_T_226 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[23] & _T_3) begin
      assert(_T_233 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[24] & _T_3) begin
      assert(_T_240 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[25] & _T_3) begin
      assert(_T_247 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[26] & _T_3) begin
      assert(_T_254 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[27] & _T_3) begin
      assert(_T_261 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[28] & _T_3) begin
      assert(_T_268 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[29] & _T_3) begin
      assert(_T_275 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[30] & _T_3) begin
      assert(_T_282 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[31] & _T_3) begin
      assert(_T_289 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[32] & _T_3) begin
      assert(_T_296 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[33] & _T_3) begin
      assert(_T_303 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[34] & _T_3) begin
      assert(_T_310 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[35] & _T_3) begin
      assert(_T_317 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[36] & _T_3) begin
      assert(_T_324 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[37] & _T_3) begin
      assert(_T_331 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[38] & _T_3) begin
      assert(_T_338 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[39] & _T_3) begin
      assert(_T_345 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[40] & _T_3) begin
      assert(_T_352 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[41] & _T_3) begin
      assert(_T_359 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[42] & _T_3) begin
      assert(_T_366 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[43] & _T_3) begin
      assert(_T_373 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[44] & _T_3) begin
      assert(_T_380 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[45] & _T_3) begin
      assert(_T_387 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[46] & _T_3) begin
      assert(_T_394 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[47] & _T_3) begin
      assert(_T_401 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[48] & _T_3) begin
      assert(_T_408 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[49] & _T_3) begin
      assert(_T_415 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[50] & _T_3) begin
      assert(_T_422 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[51] & _T_3) begin
      assert(_T_429 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[52] & _T_3) begin
      assert(_T_436 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[53] & _T_3) begin
      assert(_T_443 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[54] & _T_3) begin
      assert(_T_450 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[55] & _T_3) begin
      assert(_T_457 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[56] & _T_3) begin
      assert(_T_464 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[57] & _T_3) begin
      assert(_T_471 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[58] & _T_3) begin
      assert(_T_478 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[59] & _T_3) begin
      assert(_T_485 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[60] & _T_3) begin
      assert(_T_492 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[61] & _T_3) begin
      assert(_T_499 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[62] & _T_3) begin
      assert(_T_506 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[63] & _T_3) begin
      assert(_T_513 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[64] & _T_3) begin
      assert(_T_520 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[65] & _T_3) begin
      assert(_T_527 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[66] & _T_3) begin
      assert(_T_534 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[67] & _T_3) begin
      assert(_T_541 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[68] & _T_3) begin
      assert(_T_548 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[69] & _T_3) begin
      assert(_T_555 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[70] & _T_3) begin
      assert(_T_562 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[71] & _T_3) begin
      assert(_T_569 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[72] & _T_3) begin
      assert(_T_576 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[73] & _T_3) begin
      assert(_T_583 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[74] & _T_3) begin
      assert(_T_590 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[75] & _T_3) begin
      assert(_T_597 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[76] & _T_3) begin
      assert(_T_604 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[77] & _T_3) begin
      assert(_T_611 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[78] & _T_3) begin
      assert(_T_618 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[79] & _T_3) begin
      assert(_T_625 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[80] & _T_3) begin
      assert(_T_632 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[81] & _T_3) begin
      assert(_T_639 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[82] & _T_3) begin
      assert(_T_646 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[83] & _T_3) begin
      assert(_T_653 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[84] & _T_3) begin
      assert(_T_660 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[85] & _T_3) begin
      assert(_T_667 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[86] & _T_3) begin
      assert(_T_674 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[87] & _T_3) begin
      assert(_T_681 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[88] & _T_3) begin
      assert(_T_688 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[89] & _T_3) begin
      assert(_T_695 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[90] & _T_3) begin
      assert(_T_702 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[91] & _T_3) begin
      assert(_T_709 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[92] & _T_3) begin
      assert(_T_716 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[93] & _T_3) begin
      assert(_T_723 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[94] & _T_3) begin
      assert(_T_730 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[95] & _T_3) begin
      assert(_T_737 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[96] & _T_3) begin
      assert(_T_744 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[97] & _T_3) begin
      assert(_T_751 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[98] & _T_3) begin
      assert(_T_758 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[99] & _T_3) begin
      assert(_T_765 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[100] & _T_3) begin
      assert(_T_772 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[101] & _T_3) begin
      assert(_T_779 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[102] & _T_3) begin
      assert(_T_786 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[103] & _T_3) begin
      assert(_T_793 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[104] & _T_3) begin
      assert(_T_800 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[105] & _T_3) begin
      assert(_T_807 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[106] & _T_3) begin
      assert(_T_814 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[107] & _T_3) begin
      assert(_T_821 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[108] & _T_3) begin
      assert(_T_828 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[109] & _T_3) begin
      assert(_T_835 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[110] & _T_3) begin
      assert(_T_842 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[111] & _T_3) begin
      assert(_T_849 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[112] & _T_3) begin
      assert(_T_856 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[113] & _T_3) begin
      assert(_T_863 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[114] & _T_3) begin
      assert(_T_870 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[115] & _T_3) begin
      assert(_T_877 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[116] & _T_3) begin
      assert(_T_884 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[117] & _T_3) begin
      assert(_T_891 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[118] & _T_3) begin
      assert(_T_898 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[119] & _T_3) begin
      assert(_T_905 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[120] & _T_3) begin
      assert(_T_912 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[121] & _T_3) begin
      assert(_T_919 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[122] & _T_3) begin
      assert(_T_926 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[123] & _T_3) begin
      assert(_T_933 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[124] & _T_3) begin
      assert(_T_940 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[125] & _T_3) begin
      assert(_T_947 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[126] & _T_3) begin
      assert(_T_954 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[127] & _T_3) begin
      assert(_T_961 < 64'h4000); // @[TestHarness.scala 229:13]
    end
  end
endmodule
module TestHarness(
  input   clock,
  input   reset,
  output  io_success
);
  wire  lazyNoC_clock; // @[TestHarness.scala 238:19]
  wire  lazyNoC_reset; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_ingress_0_flit_ready; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_ingress_0_flit_valid; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_ingress_0_flit_bits_head; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_ingress_0_flit_bits_tail; // @[TestHarness.scala 238:19]
  wire [63:0] lazyNoC_io_ingress_0_flit_bits_payload; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_ingress_0_flit_bits_egress_id; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_egress_0_flit_valid; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_egress_0_flit_bits_head; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_egress_0_flit_bits_tail; // @[TestHarness.scala 238:19]
  wire [63:0] lazyNoC_io_egress_0_flit_bits_payload; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_egress_0_flit_bits_ingress_id; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_router_clocks_0_clock; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_router_clocks_0_reset; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_router_clocks_1_clock; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_router_clocks_1_reset; // @[TestHarness.scala 238:19]
  wire  noc_tester_clock; // @[TestHarness.scala 269:26]
  wire  noc_tester_reset; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_to_noc_0_flit_ready; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_to_noc_0_flit_valid; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_to_noc_0_flit_bits_head; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_to_noc_0_flit_bits_tail; // @[TestHarness.scala 269:26]
  wire [63:0] noc_tester_io_to_noc_0_flit_bits_payload; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_to_noc_0_flit_bits_egress_id; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_from_noc_0_flit_ready; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_from_noc_0_flit_valid; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_from_noc_0_flit_bits_head; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_from_noc_0_flit_bits_tail; // @[TestHarness.scala 269:26]
  wire [63:0] noc_tester_io_from_noc_0_flit_bits_payload; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_from_noc_0_flit_bits_ingress_id; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_success; // @[TestHarness.scala 269:26]
  NoC lazyNoC ( // @[TestHarness.scala 238:19]
    .clock(lazyNoC_clock),
    .reset(lazyNoC_reset),
    .io_ingress_0_flit_ready(lazyNoC_io_ingress_0_flit_ready),
    .io_ingress_0_flit_valid(lazyNoC_io_ingress_0_flit_valid),
    .io_ingress_0_flit_bits_head(lazyNoC_io_ingress_0_flit_bits_head),
    .io_ingress_0_flit_bits_tail(lazyNoC_io_ingress_0_flit_bits_tail),
    .io_ingress_0_flit_bits_payload(lazyNoC_io_ingress_0_flit_bits_payload),
    .io_ingress_0_flit_bits_egress_id(lazyNoC_io_ingress_0_flit_bits_egress_id),
    .io_egress_0_flit_valid(lazyNoC_io_egress_0_flit_valid),
    .io_egress_0_flit_bits_head(lazyNoC_io_egress_0_flit_bits_head),
    .io_egress_0_flit_bits_tail(lazyNoC_io_egress_0_flit_bits_tail),
    .io_egress_0_flit_bits_payload(lazyNoC_io_egress_0_flit_bits_payload),
    .io_egress_0_flit_bits_ingress_id(lazyNoC_io_egress_0_flit_bits_ingress_id),
    .io_router_clocks_0_clock(lazyNoC_io_router_clocks_0_clock),
    .io_router_clocks_0_reset(lazyNoC_io_router_clocks_0_reset),
    .io_router_clocks_1_clock(lazyNoC_io_router_clocks_1_clock),
    .io_router_clocks_1_reset(lazyNoC_io_router_clocks_1_reset)
  );
  NoCTester noc_tester ( // @[TestHarness.scala 269:26]
    .clock(noc_tester_clock),
    .reset(noc_tester_reset),
    .io_to_noc_0_flit_ready(noc_tester_io_to_noc_0_flit_ready),
    .io_to_noc_0_flit_valid(noc_tester_io_to_noc_0_flit_valid),
    .io_to_noc_0_flit_bits_head(noc_tester_io_to_noc_0_flit_bits_head),
    .io_to_noc_0_flit_bits_tail(noc_tester_io_to_noc_0_flit_bits_tail),
    .io_to_noc_0_flit_bits_payload(noc_tester_io_to_noc_0_flit_bits_payload),
    .io_to_noc_0_flit_bits_egress_id(noc_tester_io_to_noc_0_flit_bits_egress_id),
    .io_from_noc_0_flit_ready(noc_tester_io_from_noc_0_flit_ready),
    .io_from_noc_0_flit_valid(noc_tester_io_from_noc_0_flit_valid),
    .io_from_noc_0_flit_bits_head(noc_tester_io_from_noc_0_flit_bits_head),
    .io_from_noc_0_flit_bits_tail(noc_tester_io_from_noc_0_flit_bits_tail),
    .io_from_noc_0_flit_bits_payload(noc_tester_io_from_noc_0_flit_bits_payload),
    .io_from_noc_0_flit_bits_ingress_id(noc_tester_io_from_noc_0_flit_bits_ingress_id),
    .io_success(noc_tester_io_success)
  );
  assign io_success = noc_tester_io_success; // @[TestHarness.scala 272:14]
  assign lazyNoC_clock = clock;
  assign lazyNoC_reset = reset;
  assign lazyNoC_io_ingress_0_flit_valid = noc_tester_io_to_noc_0_flit_valid; // @[TestHarness.scala 270:18]
  assign lazyNoC_io_ingress_0_flit_bits_head = noc_tester_io_to_noc_0_flit_bits_head; // @[TestHarness.scala 270:18]
  assign lazyNoC_io_ingress_0_flit_bits_tail = noc_tester_io_to_noc_0_flit_bits_tail; // @[TestHarness.scala 270:18]
  assign lazyNoC_io_ingress_0_flit_bits_payload = noc_tester_io_to_noc_0_flit_bits_payload; // @[TestHarness.scala 270:18]
  assign lazyNoC_io_ingress_0_flit_bits_egress_id = noc_tester_io_to_noc_0_flit_bits_egress_id; // @[TestHarness.scala 270:18]
  assign lazyNoC_io_router_clocks_0_clock = clock; // @[TestHarness.scala 239:40]
  assign lazyNoC_io_router_clocks_0_reset = reset; // @[TestHarness.scala 240:40]
  assign lazyNoC_io_router_clocks_1_clock = clock; // @[TestHarness.scala 239:40]
  assign lazyNoC_io_router_clocks_1_reset = reset; // @[TestHarness.scala 240:40]
  assign noc_tester_clock = clock;
  assign noc_tester_reset = reset;
  assign noc_tester_io_to_noc_0_flit_ready = lazyNoC_io_ingress_0_flit_ready; // @[TestHarness.scala 270:18]
  assign noc_tester_io_from_noc_0_flit_valid = lazyNoC_io_egress_0_flit_valid; // @[TestHarness.scala 271:26]
  assign noc_tester_io_from_noc_0_flit_bits_head = lazyNoC_io_egress_0_flit_bits_head; // @[TestHarness.scala 271:26]
  assign noc_tester_io_from_noc_0_flit_bits_tail = lazyNoC_io_egress_0_flit_bits_tail; // @[TestHarness.scala 271:26]
  assign noc_tester_io_from_noc_0_flit_bits_payload = lazyNoC_io_egress_0_flit_bits_payload; // @[TestHarness.scala 271:26]
  assign noc_tester_io_from_noc_0_flit_bits_ingress_id = lazyNoC_io_egress_0_flit_bits_ingress_id; // @[TestHarness.scala 271:26]
endmodule
module NoCChiselTester(
  input   clock,
  input   reset
);
  wire  th_clock; // @[NocTests.scala 11:18]
  wire  th_reset; // @[NocTests.scala 11:18]
  wire  th_io_success; // @[NocTests.scala 11:18]
  TestHarness th ( // @[NocTests.scala 11:18]
    .clock(th_clock),
    .reset(th_reset),
    .io_success(th_io_success)
  );
  assign th_clock = clock;
  assign th_reset = reset;
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (th_io_success & ~reset) begin
          $finish; // @[NocTests.scala 12:30]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
