module SoC #(
    parameter 
)
(
    input           clock,
    input           reset,

);


// VeeR-EH1



endmodule