module NoCMonitor(
  input        clock,
  input        reset,
  input        io_in_flit_0_valid,
  input        io_in_flit_0_bits_head,
  input        io_in_flit_0_bits_tail,
  input  [1:0] io_in_flit_0_bits_flow_ingress_node,
  input  [1:0] io_in_flit_0_bits_flow_egress_node,
  input  [1:0] io_in_flit_0_bits_virt_channel_id
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg  in_flight_0; // @[Monitor.scala 16:26]
  reg  in_flight_1; // @[Monitor.scala 16:26]
  reg  in_flight_2; // @[Monitor.scala 16:26]
  reg  in_flight_3; // @[Monitor.scala 16:26]
  wire  _GEN_0 = 2'h0 == io_in_flit_0_bits_virt_channel_id | in_flight_0; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_1 = 2'h1 == io_in_flit_0_bits_virt_channel_id | in_flight_1; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_2 = 2'h2 == io_in_flit_0_bits_virt_channel_id | in_flight_2; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_3 = 2'h3 == io_in_flit_0_bits_virt_channel_id | in_flight_3; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_5 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? in_flight_1 : in_flight_0; // @[Monitor.scala 22:{17,17}]
  wire  _GEN_6 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? in_flight_2 : _GEN_5; // @[Monitor.scala 22:{17,17}]
  wire  _GEN_7 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? in_flight_3 : _GEN_6; // @[Monitor.scala 22:{17,17}]
  wire  _T_2 = ~reset; // @[Monitor.scala 22:16]
  wire  _GEN_8 = io_in_flit_0_bits_head ? _GEN_0 : in_flight_0; // @[Monitor.scala 16:26 20:29]
  wire  _GEN_9 = io_in_flit_0_bits_head ? _GEN_1 : in_flight_1; // @[Monitor.scala 16:26 20:29]
  wire  _GEN_10 = io_in_flit_0_bits_head ? _GEN_2 : in_flight_2; // @[Monitor.scala 16:26 20:29]
  wire  _GEN_11 = io_in_flit_0_bits_head ? _GEN_3 : in_flight_3; // @[Monitor.scala 16:26 20:29]
  wire  _T_4 = io_in_flit_0_valid & io_in_flit_0_bits_head; // @[Monitor.scala 29:22]
  wire  _T_7 = io_in_flit_0_bits_flow_egress_node == 2'h0; // @[Types.scala 54:21]
  wire  _T_8 = io_in_flit_0_bits_flow_ingress_node == 2'h2 & _T_7; // @[Types.scala 53:39]
  wire  _T_20 = io_in_flit_0_bits_flow_ingress_node == 2'h1 & _T_7; // @[Types.scala 53:39]
  wire  _T_26 = io_in_flit_0_bits_flow_egress_node == 2'h3; // @[Types.scala 54:21]
  wire  _T_27 = io_in_flit_0_bits_flow_ingress_node == 2'h1 & _T_26; // @[Types.scala 53:39]
  wire  _T_40 = _T_20 | _T_27 | _T_8; // @[package.scala 73:59]
  wire  _GEN_29 = _T_4 & ~reset; // @[Monitor.scala 22:16]
  always @(posedge clock) begin
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_0 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h0 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_0 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_0 <= _GEN_8;
        end
      end else begin
        in_flight_0 <= _GEN_8;
      end
    end
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_1 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h1 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_1 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_1 <= _GEN_9;
        end
      end else begin
        in_flight_1 <= _GEN_9;
      end
    end
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_2 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h2 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_2 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_2 <= _GEN_10;
        end
      end else begin
        in_flight_2 <= _GEN_10;
      end
    end
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_3 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h3 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_3 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_3 <= _GEN_11;
        end
      end else begin
        in_flight_3 <= _GEN_11;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4 & ~reset & ~(~_GEN_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed: Flit head/tail sequencing is broken\n    at Monitor.scala:22 assert (!in_flight(flit.bits.virt_channel_id), \"Flit head/tail sequencing is broken\")\n"
            ); // @[Monitor.scala 22:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h0 | _T_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h1 | _T_40)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h2 | _T_40)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h3 | _T_40)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  in_flight_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  in_flight_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  in_flight_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  in_flight_3 = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (_T_4 & ~reset) begin
      assert(~_GEN_7); // @[Monitor.scala 22:16]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h0 | _T_8); // @[Monitor.scala 32:17]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h1 | _T_40); // @[Monitor.scala 32:17]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h2 | _T_40); // @[Monitor.scala 32:17]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h3 | _T_40); // @[Monitor.scala 32:17]
    end
  end
endmodule
module NoCMonitor_1(
  input        clock,
  input        reset,
  input        io_in_flit_0_valid,
  input        io_in_flit_0_bits_head,
  input        io_in_flit_0_bits_tail,
  input  [1:0] io_in_flit_0_bits_flow_ingress_node,
  input  [1:0] io_in_flit_0_bits_flow_egress_node,
  input  [1:0] io_in_flit_0_bits_virt_channel_id
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg  in_flight_0; // @[Monitor.scala 16:26]
  reg  in_flight_1; // @[Monitor.scala 16:26]
  reg  in_flight_2; // @[Monitor.scala 16:26]
  reg  in_flight_3; // @[Monitor.scala 16:26]
  wire  _GEN_0 = 2'h0 == io_in_flit_0_bits_virt_channel_id | in_flight_0; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_1 = 2'h1 == io_in_flit_0_bits_virt_channel_id | in_flight_1; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_2 = 2'h2 == io_in_flit_0_bits_virt_channel_id | in_flight_2; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_3 = 2'h3 == io_in_flit_0_bits_virt_channel_id | in_flight_3; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_5 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? in_flight_1 : in_flight_0; // @[Monitor.scala 22:{17,17}]
  wire  _GEN_6 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? in_flight_2 : _GEN_5; // @[Monitor.scala 22:{17,17}]
  wire  _GEN_7 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? in_flight_3 : _GEN_6; // @[Monitor.scala 22:{17,17}]
  wire  _T_2 = ~reset; // @[Monitor.scala 22:16]
  wire  _GEN_8 = io_in_flit_0_bits_head ? _GEN_0 : in_flight_0; // @[Monitor.scala 16:26 20:29]
  wire  _GEN_9 = io_in_flit_0_bits_head ? _GEN_1 : in_flight_1; // @[Monitor.scala 16:26 20:29]
  wire  _GEN_10 = io_in_flit_0_bits_head ? _GEN_2 : in_flight_2; // @[Monitor.scala 16:26 20:29]
  wire  _GEN_11 = io_in_flit_0_bits_head ? _GEN_3 : in_flight_3; // @[Monitor.scala 16:26 20:29]
  wire  _T_4 = io_in_flit_0_valid & io_in_flit_0_bits_head; // @[Monitor.scala 29:22]
  wire  _T_7 = io_in_flit_0_bits_flow_egress_node == 2'h0; // @[Types.scala 54:21]
  wire  _T_8 = io_in_flit_0_bits_flow_ingress_node == 2'h2 & _T_7; // @[Types.scala 53:39]
  wire  _T_27 = io_in_flit_0_bits_flow_ingress_node == 2'h3 & _T_7; // @[Types.scala 53:39]
  wire  _T_33 = io_in_flit_0_bits_flow_egress_node == 2'h1; // @[Types.scala 54:21]
  wire  _T_34 = io_in_flit_0_bits_flow_ingress_node == 2'h3 & _T_33; // @[Types.scala 53:39]
  wire  _T_40 = _T_8 | _T_27 | _T_34; // @[package.scala 73:59]
  wire  _T_88 = _T_27 | _T_34; // @[package.scala 73:59]
  wire  _GEN_29 = _T_4 & ~reset; // @[Monitor.scala 22:16]
  always @(posedge clock) begin
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_0 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h0 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_0 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_0 <= _GEN_8;
        end
      end else begin
        in_flight_0 <= _GEN_8;
      end
    end
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_1 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h1 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_1 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_1 <= _GEN_9;
        end
      end else begin
        in_flight_1 <= _GEN_9;
      end
    end
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_2 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h2 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_2 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_2 <= _GEN_10;
        end
      end else begin
        in_flight_2 <= _GEN_10;
      end
    end
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_3 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h3 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_3 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_3 <= _GEN_11;
        end
      end else begin
        in_flight_3 <= _GEN_11;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4 & ~reset & ~(~_GEN_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed: Flit head/tail sequencing is broken\n    at Monitor.scala:22 assert (!in_flight(flit.bits.virt_channel_id), \"Flit head/tail sequencing is broken\")\n"
            ); // @[Monitor.scala 22:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h0 | _T_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h1 | _T_40)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h2 | _T_40)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h3 | _T_88)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  in_flight_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  in_flight_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  in_flight_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  in_flight_3 = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (_T_4 & ~reset) begin
      assert(~_GEN_7); // @[Monitor.scala 22:16]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h0 | _T_8); // @[Monitor.scala 32:17]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h1 | _T_40); // @[Monitor.scala 32:17]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h2 | _T_40); // @[Monitor.scala 32:17]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h3 | _T_88); // @[Monitor.scala 32:17]
    end
  end
endmodule
module Queue(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_head,
  input         io_enq_bits_tail,
  input  [63:0] io_enq_bits_payload,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_head,
  output        io_deq_bits_tail,
  output [63:0] io_deq_bits_payload
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg  ram_head [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_head_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_head_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_head_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_tail [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_tail_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_tail_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_tail_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_en; // @[Decoupled.scala 273:95]
  reg [63:0] ram_payload [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_payload_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_payload_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [63:0] ram_payload_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [63:0] ram_payload_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_payload_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_payload_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_payload_MPORT_en; // @[Decoupled.scala 273:95]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 278:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  assign ram_head_io_deq_bits_MPORT_en = 1'h1;
  assign ram_head_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_head_io_deq_bits_MPORT_data = ram_head[ram_head_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_head_MPORT_data = io_enq_bits_head;
  assign ram_head_MPORT_addr = 1'h0;
  assign ram_head_MPORT_mask = 1'h1;
  assign ram_head_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tail_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tail_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tail_io_deq_bits_MPORT_data = ram_tail[ram_tail_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_tail_MPORT_data = io_enq_bits_tail;
  assign ram_tail_MPORT_addr = 1'h0;
  assign ram_tail_MPORT_mask = 1'h1;
  assign ram_tail_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_payload_io_deq_bits_MPORT_en = 1'h1;
  assign ram_payload_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_payload_io_deq_bits_MPORT_data = ram_payload[ram_payload_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_payload_MPORT_data = io_enq_bits_payload;
  assign ram_payload_MPORT_addr = 1'h0;
  assign ram_payload_MPORT_mask = 1'h1;
  assign ram_payload_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = io_deq_ready | empty; // @[Decoupled.scala 303:16 323:{24,39}]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_head = ram_head_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_tail = ram_tail_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_payload = ram_payload_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  always @(posedge clock) begin
    if (ram_head_MPORT_en & ram_head_MPORT_mask) begin
      ram_head[ram_head_MPORT_addr] <= ram_head_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_tail_MPORT_en & ram_tail_MPORT_mask) begin
      ram_tail[ram_tail_MPORT_addr] <= ram_tail_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_payload_MPORT_en & ram_payload_MPORT_mask) begin
      ram_payload[ram_payload_MPORT_addr] <= ram_payload_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_head[initvar] = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tail[initvar] = _RAND_1[0:0];
  _RAND_2 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload[initvar] = _RAND_2[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module InputBuffer(
  input         clock,
  input         reset,
  input         io_enq_0_valid,
  input         io_enq_0_bits_head,
  input         io_enq_0_bits_tail,
  input  [63:0] io_enq_0_bits_payload,
  input  [1:0]  io_enq_0_bits_virt_channel_id,
  input         io_deq_0_ready,
  output        io_deq_0_valid,
  output        io_deq_0_bits_head,
  output        io_deq_0_bits_tail,
  output [63:0] io_deq_0_bits_payload,
  input         io_deq_1_ready,
  output        io_deq_1_valid,
  output        io_deq_1_bits_head,
  output        io_deq_1_bits_tail,
  output [63:0] io_deq_1_bits_payload,
  input         io_deq_2_ready,
  output        io_deq_2_valid,
  output        io_deq_2_bits_head,
  output        io_deq_2_bits_tail,
  output [63:0] io_deq_2_bits_payload,
  input         io_deq_3_ready,
  output        io_deq_3_valid,
  output        io_deq_3_bits_head,
  output        io_deq_3_bits_tail,
  output [63:0] io_deq_3_bits_payload
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_10;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
`endif // RANDOMIZE_REG_INIT
  reg  mem_head [0:19]; // @[InputUnit.scala 85:18]
  wire  mem_head_qs_0_io_enq_bits_MPORT_en; // @[InputUnit.scala 85:18]
  wire [4:0] mem_head_qs_0_io_enq_bits_MPORT_addr; // @[InputUnit.scala 85:18]
  wire  mem_head_qs_0_io_enq_bits_MPORT_data; // @[InputUnit.scala 85:18]
  wire  mem_head_qs_1_io_enq_bits_MPORT_en; // @[InputUnit.scala 85:18]
  wire [4:0] mem_head_qs_1_io_enq_bits_MPORT_addr; // @[InputUnit.scala 85:18]
  wire  mem_head_qs_1_io_enq_bits_MPORT_data; // @[InputUnit.scala 85:18]
  wire  mem_head_qs_2_io_enq_bits_MPORT_en; // @[InputUnit.scala 85:18]
  wire [4:0] mem_head_qs_2_io_enq_bits_MPORT_addr; // @[InputUnit.scala 85:18]
  wire  mem_head_qs_2_io_enq_bits_MPORT_data; // @[InputUnit.scala 85:18]
  wire  mem_head_qs_3_io_enq_bits_MPORT_en; // @[InputUnit.scala 85:18]
  wire [4:0] mem_head_qs_3_io_enq_bits_MPORT_addr; // @[InputUnit.scala 85:18]
  wire  mem_head_qs_3_io_enq_bits_MPORT_data; // @[InputUnit.scala 85:18]
  wire  mem_head_MPORT_data; // @[InputUnit.scala 85:18]
  wire [4:0] mem_head_MPORT_addr; // @[InputUnit.scala 85:18]
  wire  mem_head_MPORT_mask; // @[InputUnit.scala 85:18]
  wire  mem_head_MPORT_en; // @[InputUnit.scala 85:18]
  reg  mem_tail [0:19]; // @[InputUnit.scala 85:18]
  wire  mem_tail_qs_0_io_enq_bits_MPORT_en; // @[InputUnit.scala 85:18]
  wire [4:0] mem_tail_qs_0_io_enq_bits_MPORT_addr; // @[InputUnit.scala 85:18]
  wire  mem_tail_qs_0_io_enq_bits_MPORT_data; // @[InputUnit.scala 85:18]
  wire  mem_tail_qs_1_io_enq_bits_MPORT_en; // @[InputUnit.scala 85:18]
  wire [4:0] mem_tail_qs_1_io_enq_bits_MPORT_addr; // @[InputUnit.scala 85:18]
  wire  mem_tail_qs_1_io_enq_bits_MPORT_data; // @[InputUnit.scala 85:18]
  wire  mem_tail_qs_2_io_enq_bits_MPORT_en; // @[InputUnit.scala 85:18]
  wire [4:0] mem_tail_qs_2_io_enq_bits_MPORT_addr; // @[InputUnit.scala 85:18]
  wire  mem_tail_qs_2_io_enq_bits_MPORT_data; // @[InputUnit.scala 85:18]
  wire  mem_tail_qs_3_io_enq_bits_MPORT_en; // @[InputUnit.scala 85:18]
  wire [4:0] mem_tail_qs_3_io_enq_bits_MPORT_addr; // @[InputUnit.scala 85:18]
  wire  mem_tail_qs_3_io_enq_bits_MPORT_data; // @[InputUnit.scala 85:18]
  wire  mem_tail_MPORT_data; // @[InputUnit.scala 85:18]
  wire [4:0] mem_tail_MPORT_addr; // @[InputUnit.scala 85:18]
  wire  mem_tail_MPORT_mask; // @[InputUnit.scala 85:18]
  wire  mem_tail_MPORT_en; // @[InputUnit.scala 85:18]
  reg [63:0] mem_payload [0:19]; // @[InputUnit.scala 85:18]
  wire  mem_payload_qs_0_io_enq_bits_MPORT_en; // @[InputUnit.scala 85:18]
  wire [4:0] mem_payload_qs_0_io_enq_bits_MPORT_addr; // @[InputUnit.scala 85:18]
  wire [63:0] mem_payload_qs_0_io_enq_bits_MPORT_data; // @[InputUnit.scala 85:18]
  wire  mem_payload_qs_1_io_enq_bits_MPORT_en; // @[InputUnit.scala 85:18]
  wire [4:0] mem_payload_qs_1_io_enq_bits_MPORT_addr; // @[InputUnit.scala 85:18]
  wire [63:0] mem_payload_qs_1_io_enq_bits_MPORT_data; // @[InputUnit.scala 85:18]
  wire  mem_payload_qs_2_io_enq_bits_MPORT_en; // @[InputUnit.scala 85:18]
  wire [4:0] mem_payload_qs_2_io_enq_bits_MPORT_addr; // @[InputUnit.scala 85:18]
  wire [63:0] mem_payload_qs_2_io_enq_bits_MPORT_data; // @[InputUnit.scala 85:18]
  wire  mem_payload_qs_3_io_enq_bits_MPORT_en; // @[InputUnit.scala 85:18]
  wire [4:0] mem_payload_qs_3_io_enq_bits_MPORT_addr; // @[InputUnit.scala 85:18]
  wire [63:0] mem_payload_qs_3_io_enq_bits_MPORT_data; // @[InputUnit.scala 85:18]
  wire [63:0] mem_payload_MPORT_data; // @[InputUnit.scala 85:18]
  wire [4:0] mem_payload_MPORT_addr; // @[InputUnit.scala 85:18]
  wire  mem_payload_MPORT_mask; // @[InputUnit.scala 85:18]
  wire  mem_payload_MPORT_en; // @[InputUnit.scala 85:18]
  wire  qs_0_clock; // @[InputUnit.scala 90:49]
  wire  qs_0_reset; // @[InputUnit.scala 90:49]
  wire  qs_0_io_enq_ready; // @[InputUnit.scala 90:49]
  wire  qs_0_io_enq_valid; // @[InputUnit.scala 90:49]
  wire  qs_0_io_enq_bits_head; // @[InputUnit.scala 90:49]
  wire  qs_0_io_enq_bits_tail; // @[InputUnit.scala 90:49]
  wire [63:0] qs_0_io_enq_bits_payload; // @[InputUnit.scala 90:49]
  wire  qs_0_io_deq_ready; // @[InputUnit.scala 90:49]
  wire  qs_0_io_deq_valid; // @[InputUnit.scala 90:49]
  wire  qs_0_io_deq_bits_head; // @[InputUnit.scala 90:49]
  wire  qs_0_io_deq_bits_tail; // @[InputUnit.scala 90:49]
  wire [63:0] qs_0_io_deq_bits_payload; // @[InputUnit.scala 90:49]
  wire  qs_1_clock; // @[InputUnit.scala 90:49]
  wire  qs_1_reset; // @[InputUnit.scala 90:49]
  wire  qs_1_io_enq_ready; // @[InputUnit.scala 90:49]
  wire  qs_1_io_enq_valid; // @[InputUnit.scala 90:49]
  wire  qs_1_io_enq_bits_head; // @[InputUnit.scala 90:49]
  wire  qs_1_io_enq_bits_tail; // @[InputUnit.scala 90:49]
  wire [63:0] qs_1_io_enq_bits_payload; // @[InputUnit.scala 90:49]
  wire  qs_1_io_deq_ready; // @[InputUnit.scala 90:49]
  wire  qs_1_io_deq_valid; // @[InputUnit.scala 90:49]
  wire  qs_1_io_deq_bits_head; // @[InputUnit.scala 90:49]
  wire  qs_1_io_deq_bits_tail; // @[InputUnit.scala 90:49]
  wire [63:0] qs_1_io_deq_bits_payload; // @[InputUnit.scala 90:49]
  wire  qs_2_clock; // @[InputUnit.scala 90:49]
  wire  qs_2_reset; // @[InputUnit.scala 90:49]
  wire  qs_2_io_enq_ready; // @[InputUnit.scala 90:49]
  wire  qs_2_io_enq_valid; // @[InputUnit.scala 90:49]
  wire  qs_2_io_enq_bits_head; // @[InputUnit.scala 90:49]
  wire  qs_2_io_enq_bits_tail; // @[InputUnit.scala 90:49]
  wire [63:0] qs_2_io_enq_bits_payload; // @[InputUnit.scala 90:49]
  wire  qs_2_io_deq_ready; // @[InputUnit.scala 90:49]
  wire  qs_2_io_deq_valid; // @[InputUnit.scala 90:49]
  wire  qs_2_io_deq_bits_head; // @[InputUnit.scala 90:49]
  wire  qs_2_io_deq_bits_tail; // @[InputUnit.scala 90:49]
  wire [63:0] qs_2_io_deq_bits_payload; // @[InputUnit.scala 90:49]
  wire  qs_3_clock; // @[InputUnit.scala 90:49]
  wire  qs_3_reset; // @[InputUnit.scala 90:49]
  wire  qs_3_io_enq_ready; // @[InputUnit.scala 90:49]
  wire  qs_3_io_enq_valid; // @[InputUnit.scala 90:49]
  wire  qs_3_io_enq_bits_head; // @[InputUnit.scala 90:49]
  wire  qs_3_io_enq_bits_tail; // @[InputUnit.scala 90:49]
  wire [63:0] qs_3_io_enq_bits_payload; // @[InputUnit.scala 90:49]
  wire  qs_3_io_deq_ready; // @[InputUnit.scala 90:49]
  wire  qs_3_io_deq_valid; // @[InputUnit.scala 90:49]
  wire  qs_3_io_deq_bits_head; // @[InputUnit.scala 90:49]
  wire  qs_3_io_deq_bits_tail; // @[InputUnit.scala 90:49]
  wire [63:0] qs_3_io_deq_bits_payload; // @[InputUnit.scala 90:49]
  reg [4:0] heads_0; // @[InputUnit.scala 86:24]
  reg [4:0] heads_1; // @[InputUnit.scala 86:24]
  reg [4:0] heads_2; // @[InputUnit.scala 86:24]
  reg [4:0] heads_3; // @[InputUnit.scala 86:24]
  reg [4:0] tails_0; // @[InputUnit.scala 87:24]
  reg [4:0] tails_1; // @[InputUnit.scala 87:24]
  reg [4:0] tails_2; // @[InputUnit.scala 87:24]
  reg [4:0] tails_3; // @[InputUnit.scala 87:24]
  wire  empty_0 = heads_0 == tails_0; // @[InputUnit.scala 88:49]
  wire  empty_1 = heads_1 == tails_1; // @[InputUnit.scala 88:49]
  wire  empty_2 = heads_2 == tails_2; // @[InputUnit.scala 88:49]
  wire  empty_3 = heads_3 == tails_3; // @[InputUnit.scala 88:49]
  wire [3:0] vc_sel = 4'h1 << io_enq_0_bits_virt_channel_id; // @[OneHot.scala 57:35]
  wire  _direct_to_q_T_10 = vc_sel[0] & qs_0_io_enq_ready | vc_sel[1] & qs_1_io_enq_ready | vc_sel[2] &
    qs_2_io_enq_ready | vc_sel[3] & qs_3_io_enq_ready; // @[Mux.scala 27:73]
  wire  _direct_to_q_T_21 = vc_sel[0] & empty_0 | vc_sel[1] & empty_1 | vc_sel[2] & empty_2 | vc_sel[3] & empty_3; // @[Mux.scala 27:73]
  wire  direct_to_q = _direct_to_q_T_10 & _direct_to_q_T_21; // @[InputUnit.scala 96:62]
  wire  _T = ~direct_to_q; // @[InputUnit.scala 100:30]
  wire [4:0] _GEN_1 = 2'h1 == io_enq_0_bits_virt_channel_id ? tails_1 : tails_0; // @[]
  wire [4:0] _GEN_2 = 2'h2 == io_enq_0_bits_virt_channel_id ? tails_2 : _GEN_1; // @[]
  wire [4:0] _GEN_3 = 2'h3 == io_enq_0_bits_virt_channel_id ? tails_3 : _GEN_2; // @[]
  wire [2:0] _tails_T_4 = vc_sel[0] ? 3'h4 : 3'h0; // @[Mux.scala 27:73]
  wire [3:0] _tails_T_5 = vc_sel[1] ? 4'h9 : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _tails_T_6 = vc_sel[2] ? 4'he : 4'h0; // @[Mux.scala 27:73]
  wire [4:0] _tails_T_7 = vc_sel[3] ? 5'h13 : 5'h0; // @[Mux.scala 27:73]
  wire [3:0] _GEN_131 = {{1'd0}, _tails_T_4}; // @[Mux.scala 27:73]
  wire [3:0] _tails_T_8 = _GEN_131 | _tails_T_5; // @[Mux.scala 27:73]
  wire [3:0] _tails_T_9 = _tails_T_8 | _tails_T_6; // @[Mux.scala 27:73]
  wire [4:0] _GEN_132 = {{1'd0}, _tails_T_9}; // @[Mux.scala 27:73]
  wire [4:0] _tails_T_10 = _GEN_132 | _tails_T_7; // @[Mux.scala 27:73]
  wire  _tails_T_11 = _GEN_3 == _tails_T_10; // @[InputUnit.scala 104:14]
  wire [2:0] _tails_T_17 = vc_sel[1] ? 3'h5 : 3'h0; // @[Mux.scala 27:73]
  wire [3:0] _tails_T_18 = vc_sel[2] ? 4'ha : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _tails_T_19 = vc_sel[3] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _GEN_133 = {{1'd0}, _tails_T_17}; // @[Mux.scala 27:73]
  wire [3:0] _tails_T_21 = _GEN_133 | _tails_T_18; // @[Mux.scala 27:73]
  wire [3:0] _tails_T_22 = _tails_T_21 | _tails_T_19; // @[Mux.scala 27:73]
  wire [4:0] _tails_T_24 = _GEN_3 + 5'h1; // @[InputUnit.scala 106:14]
  wire  _T_3 = io_enq_0_bits_virt_channel_id == 2'h0; // @[InputUnit.scala 109:46]
  wire  _T_4 = io_enq_0_bits_virt_channel_id == 2'h1; // @[InputUnit.scala 109:46]
  wire  _T_5 = io_enq_0_bits_virt_channel_id == 2'h2; // @[InputUnit.scala 109:46]
  wire  _T_6 = io_enq_0_bits_virt_channel_id == 2'h3; // @[InputUnit.scala 109:46]
  wire  _GEN_24 = io_enq_0_valid & direct_to_q & _T_3; // @[InputUnit.scala 107:50 91:31]
  wire  _GEN_28 = io_enq_0_valid & direct_to_q & _T_4; // @[InputUnit.scala 107:50 91:31]
  wire  _GEN_32 = io_enq_0_valid & direct_to_q & _T_5; // @[InputUnit.scala 107:50 91:31]
  wire  _GEN_36 = io_enq_0_valid & direct_to_q & _T_6; // @[InputUnit.scala 107:50 91:31]
  wire  _GEN_51 = io_enq_0_valid & ~direct_to_q ? 1'h0 : _GEN_24; // @[InputUnit.scala 100:44 91:31]
  wire  _GEN_55 = io_enq_0_valid & ~direct_to_q ? 1'h0 : _GEN_28; // @[InputUnit.scala 100:44 91:31]
  wire  _GEN_59 = io_enq_0_valid & ~direct_to_q ? 1'h0 : _GEN_32; // @[InputUnit.scala 100:44 91:31]
  wire  _GEN_63 = io_enq_0_valid & ~direct_to_q ? 1'h0 : _GEN_36; // @[InputUnit.scala 100:44 91:31]
  wire  can_to_q_0 = ~empty_0 & qs_0_io_enq_ready; // @[InputUnit.scala 117:70]
  wire  can_to_q_1 = ~empty_1 & qs_1_io_enq_ready; // @[InputUnit.scala 117:70]
  wire  can_to_q_2 = ~empty_2 & qs_2_io_enq_ready; // @[InputUnit.scala 117:70]
  wire  can_to_q_3 = ~empty_3 & qs_3_io_enq_ready; // @[InputUnit.scala 117:70]
  wire [3:0] _to_q_oh_enc_T = can_to_q_3 ? 4'h8 : 4'h0; // @[Mux.scala 47:70]
  wire [3:0] _to_q_oh_enc_T_1 = can_to_q_2 ? 4'h4 : _to_q_oh_enc_T; // @[Mux.scala 47:70]
  wire [3:0] _to_q_oh_enc_T_2 = can_to_q_1 ? 4'h2 : _to_q_oh_enc_T_1; // @[Mux.scala 47:70]
  wire [3:0] to_q_oh_enc = can_to_q_0 ? 4'h1 : _to_q_oh_enc_T_2; // @[Mux.scala 47:70]
  wire  to_q_oh_0 = to_q_oh_enc[0]; // @[OneHot.scala 82:30]
  wire  to_q_oh_1 = to_q_oh_enc[1]; // @[OneHot.scala 82:30]
  wire  to_q_oh_2 = to_q_oh_enc[2]; // @[OneHot.scala 82:30]
  wire  to_q_oh_3 = to_q_oh_enc[3]; // @[OneHot.scala 82:30]
  wire [3:0] _to_q_T = {to_q_oh_3,to_q_oh_2,to_q_oh_1,to_q_oh_0}; // @[Cat.scala 33:92]
  wire [1:0] to_q_hi_1 = _to_q_T[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] to_q_lo_1 = _to_q_T[1:0]; // @[OneHot.scala 31:18]
  wire  _to_q_T_1 = |to_q_hi_1; // @[OneHot.scala 32:14]
  wire [1:0] _to_q_T_2 = to_q_hi_1 | to_q_lo_1; // @[OneHot.scala 32:28]
  wire [1:0] to_q = {_to_q_T_1,_to_q_T_2[1]}; // @[Cat.scala 33:92]
  wire  _T_9 = can_to_q_0 | can_to_q_1 | can_to_q_2 | can_to_q_3; // @[package.scala 73:59]
  wire [4:0] _head_T = to_q_oh_0 ? heads_0 : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _head_T_1 = to_q_oh_1 ? heads_1 : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _head_T_2 = to_q_oh_2 ? heads_2 : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _head_T_3 = to_q_oh_3 ? heads_3 : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _head_T_4 = _head_T | _head_T_1; // @[Mux.scala 27:73]
  wire [4:0] _head_T_5 = _head_T_4 | _head_T_2; // @[Mux.scala 27:73]
  wire [4:0] head = _head_T_5 | _head_T_3; // @[Mux.scala 27:73]
  wire [2:0] _heads_T = to_q_oh_0 ? 3'h4 : 3'h0; // @[Mux.scala 27:73]
  wire [3:0] _heads_T_1 = to_q_oh_1 ? 4'h9 : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _heads_T_2 = to_q_oh_2 ? 4'he : 4'h0; // @[Mux.scala 27:73]
  wire [4:0] _heads_T_3 = to_q_oh_3 ? 5'h13 : 5'h0; // @[Mux.scala 27:73]
  wire [3:0] _GEN_134 = {{1'd0}, _heads_T}; // @[Mux.scala 27:73]
  wire [3:0] _heads_T_4 = _GEN_134 | _heads_T_1; // @[Mux.scala 27:73]
  wire [3:0] _heads_T_5 = _heads_T_4 | _heads_T_2; // @[Mux.scala 27:73]
  wire [4:0] _GEN_135 = {{1'd0}, _heads_T_5}; // @[Mux.scala 27:73]
  wire [4:0] _heads_T_6 = _GEN_135 | _heads_T_3; // @[Mux.scala 27:73]
  wire  _heads_T_7 = head == _heads_T_6; // @[InputUnit.scala 123:16]
  wire [2:0] _heads_T_9 = to_q_oh_1 ? 3'h5 : 3'h0; // @[Mux.scala 27:73]
  wire [3:0] _heads_T_10 = to_q_oh_2 ? 4'ha : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _heads_T_11 = to_q_oh_3 ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _GEN_136 = {{1'd0}, _heads_T_9}; // @[Mux.scala 27:73]
  wire [3:0] _heads_T_13 = _GEN_136 | _heads_T_10; // @[Mux.scala 27:73]
  wire [3:0] _heads_T_14 = _heads_T_13 | _heads_T_11; // @[Mux.scala 27:73]
  wire [4:0] _heads_T_16 = head + 5'h1; // @[InputUnit.scala 125:16]
  wire  _GEN_71 = to_q_oh_0 | _GEN_51; // @[InputUnit.scala 127:29 128:32]
  wire [63:0] _GEN_75 = to_q_oh_0 ? mem_payload_qs_0_io_enq_bits_MPORT_data : io_enq_0_bits_payload; // @[InputUnit.scala 127:29 129:31]
  wire  _GEN_76 = to_q_oh_0 ? mem_tail_qs_0_io_enq_bits_MPORT_data : io_enq_0_bits_tail; // @[InputUnit.scala 127:29 129:31]
  wire  _GEN_77 = to_q_oh_0 ? mem_head_qs_0_io_enq_bits_MPORT_data : io_enq_0_bits_head; // @[InputUnit.scala 127:29 129:31]
  wire  _GEN_78 = to_q_oh_1 | _GEN_55; // @[InputUnit.scala 127:29 128:32]
  wire [63:0] _GEN_82 = to_q_oh_1 ? mem_payload_qs_1_io_enq_bits_MPORT_data : io_enq_0_bits_payload; // @[InputUnit.scala 127:29 129:31]
  wire  _GEN_83 = to_q_oh_1 ? mem_tail_qs_1_io_enq_bits_MPORT_data : io_enq_0_bits_tail; // @[InputUnit.scala 127:29 129:31]
  wire  _GEN_84 = to_q_oh_1 ? mem_head_qs_1_io_enq_bits_MPORT_data : io_enq_0_bits_head; // @[InputUnit.scala 127:29 129:31]
  wire  _GEN_85 = to_q_oh_2 | _GEN_59; // @[InputUnit.scala 127:29 128:32]
  wire [63:0] _GEN_89 = to_q_oh_2 ? mem_payload_qs_2_io_enq_bits_MPORT_data : io_enq_0_bits_payload; // @[InputUnit.scala 127:29 129:31]
  wire  _GEN_90 = to_q_oh_2 ? mem_tail_qs_2_io_enq_bits_MPORT_data : io_enq_0_bits_tail; // @[InputUnit.scala 127:29 129:31]
  wire  _GEN_91 = to_q_oh_2 ? mem_head_qs_2_io_enq_bits_MPORT_data : io_enq_0_bits_head; // @[InputUnit.scala 127:29 129:31]
  wire  _GEN_92 = to_q_oh_3 | _GEN_63; // @[InputUnit.scala 127:29 128:32]
  wire [63:0] _GEN_96 = to_q_oh_3 ? mem_payload_qs_3_io_enq_bits_MPORT_data : io_enq_0_bits_payload; // @[InputUnit.scala 127:29 129:31]
  wire  _GEN_97 = to_q_oh_3 ? mem_tail_qs_3_io_enq_bits_MPORT_data : io_enq_0_bits_tail; // @[InputUnit.scala 127:29 129:31]
  wire  _GEN_98 = to_q_oh_3 ? mem_head_qs_3_io_enq_bits_MPORT_data : io_enq_0_bits_head; // @[InputUnit.scala 127:29 129:31]
  Queue qs_0 ( // @[InputUnit.scala 90:49]
    .clock(qs_0_clock),
    .reset(qs_0_reset),
    .io_enq_ready(qs_0_io_enq_ready),
    .io_enq_valid(qs_0_io_enq_valid),
    .io_enq_bits_head(qs_0_io_enq_bits_head),
    .io_enq_bits_tail(qs_0_io_enq_bits_tail),
    .io_enq_bits_payload(qs_0_io_enq_bits_payload),
    .io_deq_ready(qs_0_io_deq_ready),
    .io_deq_valid(qs_0_io_deq_valid),
    .io_deq_bits_head(qs_0_io_deq_bits_head),
    .io_deq_bits_tail(qs_0_io_deq_bits_tail),
    .io_deq_bits_payload(qs_0_io_deq_bits_payload)
  );
  Queue qs_1 ( // @[InputUnit.scala 90:49]
    .clock(qs_1_clock),
    .reset(qs_1_reset),
    .io_enq_ready(qs_1_io_enq_ready),
    .io_enq_valid(qs_1_io_enq_valid),
    .io_enq_bits_head(qs_1_io_enq_bits_head),
    .io_enq_bits_tail(qs_1_io_enq_bits_tail),
    .io_enq_bits_payload(qs_1_io_enq_bits_payload),
    .io_deq_ready(qs_1_io_deq_ready),
    .io_deq_valid(qs_1_io_deq_valid),
    .io_deq_bits_head(qs_1_io_deq_bits_head),
    .io_deq_bits_tail(qs_1_io_deq_bits_tail),
    .io_deq_bits_payload(qs_1_io_deq_bits_payload)
  );
  Queue qs_2 ( // @[InputUnit.scala 90:49]
    .clock(qs_2_clock),
    .reset(qs_2_reset),
    .io_enq_ready(qs_2_io_enq_ready),
    .io_enq_valid(qs_2_io_enq_valid),
    .io_enq_bits_head(qs_2_io_enq_bits_head),
    .io_enq_bits_tail(qs_2_io_enq_bits_tail),
    .io_enq_bits_payload(qs_2_io_enq_bits_payload),
    .io_deq_ready(qs_2_io_deq_ready),
    .io_deq_valid(qs_2_io_deq_valid),
    .io_deq_bits_head(qs_2_io_deq_bits_head),
    .io_deq_bits_tail(qs_2_io_deq_bits_tail),
    .io_deq_bits_payload(qs_2_io_deq_bits_payload)
  );
  Queue qs_3 ( // @[InputUnit.scala 90:49]
    .clock(qs_3_clock),
    .reset(qs_3_reset),
    .io_enq_ready(qs_3_io_enq_ready),
    .io_enq_valid(qs_3_io_enq_valid),
    .io_enq_bits_head(qs_3_io_enq_bits_head),
    .io_enq_bits_tail(qs_3_io_enq_bits_tail),
    .io_enq_bits_payload(qs_3_io_enq_bits_payload),
    .io_deq_ready(qs_3_io_deq_ready),
    .io_deq_valid(qs_3_io_deq_valid),
    .io_deq_bits_head(qs_3_io_deq_bits_head),
    .io_deq_bits_tail(qs_3_io_deq_bits_tail),
    .io_deq_bits_payload(qs_3_io_deq_bits_payload)
  );
  assign mem_head_qs_0_io_enq_bits_MPORT_en = _T_9 & to_q_oh_0;
  assign mem_head_qs_0_io_enq_bits_MPORT_addr = _head_T_5 | _head_T_3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_head_qs_0_io_enq_bits_MPORT_data = mem_head[mem_head_qs_0_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `else
  assign mem_head_qs_0_io_enq_bits_MPORT_data = mem_head_qs_0_io_enq_bits_MPORT_addr >= 5'h14 ? _RAND_1[0:0] :
    mem_head[mem_head_qs_0_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_head_qs_1_io_enq_bits_MPORT_en = _T_9 & to_q_oh_1;
  assign mem_head_qs_1_io_enq_bits_MPORT_addr = _head_T_5 | _head_T_3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_head_qs_1_io_enq_bits_MPORT_data = mem_head[mem_head_qs_1_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `else
  assign mem_head_qs_1_io_enq_bits_MPORT_data = mem_head_qs_1_io_enq_bits_MPORT_addr >= 5'h14 ? _RAND_2[0:0] :
    mem_head[mem_head_qs_1_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_head_qs_2_io_enq_bits_MPORT_en = _T_9 & to_q_oh_2;
  assign mem_head_qs_2_io_enq_bits_MPORT_addr = _head_T_5 | _head_T_3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_head_qs_2_io_enq_bits_MPORT_data = mem_head[mem_head_qs_2_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `else
  assign mem_head_qs_2_io_enq_bits_MPORT_data = mem_head_qs_2_io_enq_bits_MPORT_addr >= 5'h14 ? _RAND_3[0:0] :
    mem_head[mem_head_qs_2_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_head_qs_3_io_enq_bits_MPORT_en = _T_9 & to_q_oh_3;
  assign mem_head_qs_3_io_enq_bits_MPORT_addr = _head_T_5 | _head_T_3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_head_qs_3_io_enq_bits_MPORT_data = mem_head[mem_head_qs_3_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `else
  assign mem_head_qs_3_io_enq_bits_MPORT_data = mem_head_qs_3_io_enq_bits_MPORT_addr >= 5'h14 ? _RAND_4[0:0] :
    mem_head[mem_head_qs_3_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_head_MPORT_data = io_enq_0_bits_head;
  assign mem_head_MPORT_addr = 2'h3 == io_enq_0_bits_virt_channel_id ? tails_3 : _GEN_2;
  assign mem_head_MPORT_mask = 1'h1;
  assign mem_head_MPORT_en = io_enq_0_valid & _T;
  assign mem_tail_qs_0_io_enq_bits_MPORT_en = _T_9 & to_q_oh_0;
  assign mem_tail_qs_0_io_enq_bits_MPORT_addr = _head_T_5 | _head_T_3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_tail_qs_0_io_enq_bits_MPORT_data = mem_tail[mem_tail_qs_0_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `else
  assign mem_tail_qs_0_io_enq_bits_MPORT_data = mem_tail_qs_0_io_enq_bits_MPORT_addr >= 5'h14 ? _RAND_6[0:0] :
    mem_tail[mem_tail_qs_0_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_tail_qs_1_io_enq_bits_MPORT_en = _T_9 & to_q_oh_1;
  assign mem_tail_qs_1_io_enq_bits_MPORT_addr = _head_T_5 | _head_T_3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_tail_qs_1_io_enq_bits_MPORT_data = mem_tail[mem_tail_qs_1_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `else
  assign mem_tail_qs_1_io_enq_bits_MPORT_data = mem_tail_qs_1_io_enq_bits_MPORT_addr >= 5'h14 ? _RAND_7[0:0] :
    mem_tail[mem_tail_qs_1_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_tail_qs_2_io_enq_bits_MPORT_en = _T_9 & to_q_oh_2;
  assign mem_tail_qs_2_io_enq_bits_MPORT_addr = _head_T_5 | _head_T_3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_tail_qs_2_io_enq_bits_MPORT_data = mem_tail[mem_tail_qs_2_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `else
  assign mem_tail_qs_2_io_enq_bits_MPORT_data = mem_tail_qs_2_io_enq_bits_MPORT_addr >= 5'h14 ? _RAND_8[0:0] :
    mem_tail[mem_tail_qs_2_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_tail_qs_3_io_enq_bits_MPORT_en = _T_9 & to_q_oh_3;
  assign mem_tail_qs_3_io_enq_bits_MPORT_addr = _head_T_5 | _head_T_3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_tail_qs_3_io_enq_bits_MPORT_data = mem_tail[mem_tail_qs_3_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `else
  assign mem_tail_qs_3_io_enq_bits_MPORT_data = mem_tail_qs_3_io_enq_bits_MPORT_addr >= 5'h14 ? _RAND_9[0:0] :
    mem_tail[mem_tail_qs_3_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_tail_MPORT_data = io_enq_0_bits_tail;
  assign mem_tail_MPORT_addr = 2'h3 == io_enq_0_bits_virt_channel_id ? tails_3 : _GEN_2;
  assign mem_tail_MPORT_mask = 1'h1;
  assign mem_tail_MPORT_en = io_enq_0_valid & _T;
  assign mem_payload_qs_0_io_enq_bits_MPORT_en = _T_9 & to_q_oh_0;
  assign mem_payload_qs_0_io_enq_bits_MPORT_addr = _head_T_5 | _head_T_3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_payload_qs_0_io_enq_bits_MPORT_data = mem_payload[mem_payload_qs_0_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `else
  assign mem_payload_qs_0_io_enq_bits_MPORT_data = mem_payload_qs_0_io_enq_bits_MPORT_addr >= 5'h14 ? _RAND_11[63:0] :
    mem_payload[mem_payload_qs_0_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_payload_qs_1_io_enq_bits_MPORT_en = _T_9 & to_q_oh_1;
  assign mem_payload_qs_1_io_enq_bits_MPORT_addr = _head_T_5 | _head_T_3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_payload_qs_1_io_enq_bits_MPORT_data = mem_payload[mem_payload_qs_1_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `else
  assign mem_payload_qs_1_io_enq_bits_MPORT_data = mem_payload_qs_1_io_enq_bits_MPORT_addr >= 5'h14 ? _RAND_12[63:0] :
    mem_payload[mem_payload_qs_1_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_payload_qs_2_io_enq_bits_MPORT_en = _T_9 & to_q_oh_2;
  assign mem_payload_qs_2_io_enq_bits_MPORT_addr = _head_T_5 | _head_T_3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_payload_qs_2_io_enq_bits_MPORT_data = mem_payload[mem_payload_qs_2_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `else
  assign mem_payload_qs_2_io_enq_bits_MPORT_data = mem_payload_qs_2_io_enq_bits_MPORT_addr >= 5'h14 ? _RAND_13[63:0] :
    mem_payload[mem_payload_qs_2_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_payload_qs_3_io_enq_bits_MPORT_en = _T_9 & to_q_oh_3;
  assign mem_payload_qs_3_io_enq_bits_MPORT_addr = _head_T_5 | _head_T_3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_payload_qs_3_io_enq_bits_MPORT_data = mem_payload[mem_payload_qs_3_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `else
  assign mem_payload_qs_3_io_enq_bits_MPORT_data = mem_payload_qs_3_io_enq_bits_MPORT_addr >= 5'h14 ? _RAND_14[63:0] :
    mem_payload[mem_payload_qs_3_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_payload_MPORT_data = io_enq_0_bits_payload;
  assign mem_payload_MPORT_addr = 2'h3 == io_enq_0_bits_virt_channel_id ? tails_3 : _GEN_2;
  assign mem_payload_MPORT_mask = 1'h1;
  assign mem_payload_MPORT_en = io_enq_0_valid & _T;
  assign io_deq_0_valid = qs_0_io_deq_valid; // @[InputUnit.scala 134:19]
  assign io_deq_0_bits_head = qs_0_io_deq_bits_head; // @[InputUnit.scala 134:19]
  assign io_deq_0_bits_tail = qs_0_io_deq_bits_tail; // @[InputUnit.scala 134:19]
  assign io_deq_0_bits_payload = qs_0_io_deq_bits_payload; // @[InputUnit.scala 134:19]
  assign io_deq_1_valid = qs_1_io_deq_valid; // @[InputUnit.scala 134:19]
  assign io_deq_1_bits_head = qs_1_io_deq_bits_head; // @[InputUnit.scala 134:19]
  assign io_deq_1_bits_tail = qs_1_io_deq_bits_tail; // @[InputUnit.scala 134:19]
  assign io_deq_1_bits_payload = qs_1_io_deq_bits_payload; // @[InputUnit.scala 134:19]
  assign io_deq_2_valid = qs_2_io_deq_valid; // @[InputUnit.scala 134:19]
  assign io_deq_2_bits_head = qs_2_io_deq_bits_head; // @[InputUnit.scala 134:19]
  assign io_deq_2_bits_tail = qs_2_io_deq_bits_tail; // @[InputUnit.scala 134:19]
  assign io_deq_2_bits_payload = qs_2_io_deq_bits_payload; // @[InputUnit.scala 134:19]
  assign io_deq_3_valid = qs_3_io_deq_valid; // @[InputUnit.scala 134:19]
  assign io_deq_3_bits_head = qs_3_io_deq_bits_head; // @[InputUnit.scala 134:19]
  assign io_deq_3_bits_tail = qs_3_io_deq_bits_tail; // @[InputUnit.scala 134:19]
  assign io_deq_3_bits_payload = qs_3_io_deq_bits_payload; // @[InputUnit.scala 134:19]
  assign qs_0_clock = clock;
  assign qs_0_reset = reset;
  assign qs_0_io_enq_valid = _T_9 ? _GEN_71 : _GEN_51; // @[InputUnit.scala 120:27]
  assign qs_0_io_enq_bits_head = _T_9 ? _GEN_77 : io_enq_0_bits_head; // @[InputUnit.scala 120:27]
  assign qs_0_io_enq_bits_tail = _T_9 ? _GEN_76 : io_enq_0_bits_tail; // @[InputUnit.scala 120:27]
  assign qs_0_io_enq_bits_payload = _T_9 ? _GEN_75 : io_enq_0_bits_payload; // @[InputUnit.scala 120:27]
  assign qs_0_io_deq_ready = io_deq_0_ready; // @[InputUnit.scala 134:19]
  assign qs_1_clock = clock;
  assign qs_1_reset = reset;
  assign qs_1_io_enq_valid = _T_9 ? _GEN_78 : _GEN_55; // @[InputUnit.scala 120:27]
  assign qs_1_io_enq_bits_head = _T_9 ? _GEN_84 : io_enq_0_bits_head; // @[InputUnit.scala 120:27]
  assign qs_1_io_enq_bits_tail = _T_9 ? _GEN_83 : io_enq_0_bits_tail; // @[InputUnit.scala 120:27]
  assign qs_1_io_enq_bits_payload = _T_9 ? _GEN_82 : io_enq_0_bits_payload; // @[InputUnit.scala 120:27]
  assign qs_1_io_deq_ready = io_deq_1_ready; // @[InputUnit.scala 134:19]
  assign qs_2_clock = clock;
  assign qs_2_reset = reset;
  assign qs_2_io_enq_valid = _T_9 ? _GEN_85 : _GEN_59; // @[InputUnit.scala 120:27]
  assign qs_2_io_enq_bits_head = _T_9 ? _GEN_91 : io_enq_0_bits_head; // @[InputUnit.scala 120:27]
  assign qs_2_io_enq_bits_tail = _T_9 ? _GEN_90 : io_enq_0_bits_tail; // @[InputUnit.scala 120:27]
  assign qs_2_io_enq_bits_payload = _T_9 ? _GEN_89 : io_enq_0_bits_payload; // @[InputUnit.scala 120:27]
  assign qs_2_io_deq_ready = io_deq_2_ready; // @[InputUnit.scala 134:19]
  assign qs_3_clock = clock;
  assign qs_3_reset = reset;
  assign qs_3_io_enq_valid = _T_9 ? _GEN_92 : _GEN_63; // @[InputUnit.scala 120:27]
  assign qs_3_io_enq_bits_head = _T_9 ? _GEN_98 : io_enq_0_bits_head; // @[InputUnit.scala 120:27]
  assign qs_3_io_enq_bits_tail = _T_9 ? _GEN_97 : io_enq_0_bits_tail; // @[InputUnit.scala 120:27]
  assign qs_3_io_enq_bits_payload = _T_9 ? _GEN_96 : io_enq_0_bits_payload; // @[InputUnit.scala 120:27]
  assign qs_3_io_deq_ready = io_deq_3_ready; // @[InputUnit.scala 134:19]
  always @(posedge clock) begin
    if (mem_head_MPORT_en & mem_head_MPORT_mask) begin
      mem_head[mem_head_MPORT_addr] <= mem_head_MPORT_data; // @[InputUnit.scala 85:18]
    end
    if (mem_tail_MPORT_en & mem_tail_MPORT_mask) begin
      mem_tail[mem_tail_MPORT_addr] <= mem_tail_MPORT_data; // @[InputUnit.scala 85:18]
    end
    if (mem_payload_MPORT_en & mem_payload_MPORT_mask) begin
      mem_payload[mem_payload_MPORT_addr] <= mem_payload_MPORT_data; // @[InputUnit.scala 85:18]
    end
    if (reset) begin // @[InputUnit.scala 86:24]
      heads_0 <= 5'h0; // @[InputUnit.scala 86:24]
    end else if (_T_9) begin // @[InputUnit.scala 120:27]
      if (2'h0 == to_q) begin // @[InputUnit.scala 122:21]
        if (_heads_T_7) begin // @[InputUnit.scala 122:27]
          heads_0 <= {{1'd0}, _heads_T_14};
        end else begin
          heads_0 <= _heads_T_16;
        end
      end
    end
    if (reset) begin // @[InputUnit.scala 86:24]
      heads_1 <= 5'h5; // @[InputUnit.scala 86:24]
    end else if (_T_9) begin // @[InputUnit.scala 120:27]
      if (2'h1 == to_q) begin // @[InputUnit.scala 122:21]
        if (_heads_T_7) begin // @[InputUnit.scala 122:27]
          heads_1 <= {{1'd0}, _heads_T_14};
        end else begin
          heads_1 <= _heads_T_16;
        end
      end
    end
    if (reset) begin // @[InputUnit.scala 86:24]
      heads_2 <= 5'ha; // @[InputUnit.scala 86:24]
    end else if (_T_9) begin // @[InputUnit.scala 120:27]
      if (2'h2 == to_q) begin // @[InputUnit.scala 122:21]
        if (_heads_T_7) begin // @[InputUnit.scala 122:27]
          heads_2 <= {{1'd0}, _heads_T_14};
        end else begin
          heads_2 <= _heads_T_16;
        end
      end
    end
    if (reset) begin // @[InputUnit.scala 86:24]
      heads_3 <= 5'hf; // @[InputUnit.scala 86:24]
    end else if (_T_9) begin // @[InputUnit.scala 120:27]
      if (2'h3 == to_q) begin // @[InputUnit.scala 122:21]
        if (_heads_T_7) begin // @[InputUnit.scala 122:27]
          heads_3 <= {{1'd0}, _heads_T_14};
        end else begin
          heads_3 <= _heads_T_16;
        end
      end
    end
    if (reset) begin // @[InputUnit.scala 87:24]
      tails_0 <= 5'h0; // @[InputUnit.scala 87:24]
    end else if (io_enq_0_valid & ~direct_to_q) begin // @[InputUnit.scala 100:44]
      if (2'h0 == io_enq_0_bits_virt_channel_id) begin // @[InputUnit.scala 103:45]
        if (_tails_T_11) begin // @[InputUnit.scala 103:51]
          tails_0 <= {{1'd0}, _tails_T_22};
        end else begin
          tails_0 <= _tails_T_24;
        end
      end
    end
    if (reset) begin // @[InputUnit.scala 87:24]
      tails_1 <= 5'h5; // @[InputUnit.scala 87:24]
    end else if (io_enq_0_valid & ~direct_to_q) begin // @[InputUnit.scala 100:44]
      if (2'h1 == io_enq_0_bits_virt_channel_id) begin // @[InputUnit.scala 103:45]
        if (_tails_T_11) begin // @[InputUnit.scala 103:51]
          tails_1 <= {{1'd0}, _tails_T_22};
        end else begin
          tails_1 <= _tails_T_24;
        end
      end
    end
    if (reset) begin // @[InputUnit.scala 87:24]
      tails_2 <= 5'ha; // @[InputUnit.scala 87:24]
    end else if (io_enq_0_valid & ~direct_to_q) begin // @[InputUnit.scala 100:44]
      if (2'h2 == io_enq_0_bits_virt_channel_id) begin // @[InputUnit.scala 103:45]
        if (_tails_T_11) begin // @[InputUnit.scala 103:51]
          tails_2 <= {{1'd0}, _tails_T_22};
        end else begin
          tails_2 <= _tails_T_24;
        end
      end
    end
    if (reset) begin // @[InputUnit.scala 87:24]
      tails_3 <= 5'hf; // @[InputUnit.scala 87:24]
    end else if (io_enq_0_valid & ~direct_to_q) begin // @[InputUnit.scala 100:44]
      if (2'h3 == io_enq_0_bits_virt_channel_id) begin // @[InputUnit.scala 103:45]
        if (_tails_T_11) begin // @[InputUnit.scala 103:51]
          tails_3 <= {{1'd0}, _tails_T_22};
        end else begin
          tails_3 <= _tails_T_24;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {1{`RANDOM}};
  _RAND_2 = {1{`RANDOM}};
  _RAND_3 = {1{`RANDOM}};
  _RAND_4 = {1{`RANDOM}};
  _RAND_6 = {1{`RANDOM}};
  _RAND_7 = {1{`RANDOM}};
  _RAND_8 = {1{`RANDOM}};
  _RAND_9 = {1{`RANDOM}};
  _RAND_11 = {2{`RANDOM}};
  _RAND_12 = {2{`RANDOM}};
  _RAND_13 = {2{`RANDOM}};
  _RAND_14 = {2{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 20; initvar = initvar+1)
    mem_head[initvar] = _RAND_0[0:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 20; initvar = initvar+1)
    mem_tail[initvar] = _RAND_5[0:0];
  _RAND_10 = {2{`RANDOM}};
  for (initvar = 0; initvar < 20; initvar = initvar+1)
    mem_payload[initvar] = _RAND_10[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  heads_0 = _RAND_15[4:0];
  _RAND_16 = {1{`RANDOM}};
  heads_1 = _RAND_16[4:0];
  _RAND_17 = {1{`RANDOM}};
  heads_2 = _RAND_17[4:0];
  _RAND_18 = {1{`RANDOM}};
  heads_3 = _RAND_18[4:0];
  _RAND_19 = {1{`RANDOM}};
  tails_0 = _RAND_19[4:0];
  _RAND_20 = {1{`RANDOM}};
  tails_1 = _RAND_20[4:0];
  _RAND_21 = {1{`RANDOM}};
  tails_2 = _RAND_21[4:0];
  _RAND_22 = {1{`RANDOM}};
  tails_3 = _RAND_22[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Arbiter(
  input        io_in_0_valid,
  input  [1:0] io_in_0_bits_flow_ingress_node,
  input  [1:0] io_in_0_bits_flow_egress_node,
  output       io_in_1_ready,
  input        io_in_1_valid,
  input  [1:0] io_in_1_bits_flow_ingress_node,
  input  [1:0] io_in_1_bits_flow_egress_node,
  output       io_in_2_ready,
  input        io_in_2_valid,
  input  [1:0] io_in_2_bits_flow_ingress_node,
  input  [1:0] io_in_2_bits_flow_egress_node,
  output       io_in_3_ready,
  input        io_in_3_valid,
  input  [1:0] io_in_3_bits_flow_ingress_node,
  input  [1:0] io_in_3_bits_flow_egress_node,
  output       io_out_valid,
  output [1:0] io_out_bits_src_virt_id,
  output [1:0] io_out_bits_flow_ingress_node,
  output [1:0] io_out_bits_flow_egress_node
);
  wire [1:0] _GEN_0 = io_in_2_valid ? 2'h2 : 2'h3; // @[Arbiter.scala 135:13 138:26 139:17]
  wire [1:0] _GEN_3 = io_in_2_valid ? io_in_2_bits_flow_ingress_node : io_in_3_bits_flow_ingress_node; // @[Arbiter.scala 136:15 138:26 140:19]
  wire [1:0] _GEN_5 = io_in_2_valid ? io_in_2_bits_flow_egress_node : io_in_3_bits_flow_egress_node; // @[Arbiter.scala 136:15 138:26 140:19]
  wire [1:0] _GEN_7 = io_in_1_valid ? 2'h1 : _GEN_0; // @[Arbiter.scala 138:26 139:17]
  wire [1:0] _GEN_10 = io_in_1_valid ? io_in_1_bits_flow_ingress_node : _GEN_3; // @[Arbiter.scala 138:26 140:19]
  wire [1:0] _GEN_12 = io_in_1_valid ? io_in_1_bits_flow_egress_node : _GEN_5; // @[Arbiter.scala 138:26 140:19]
  wire  grant_3 = ~(io_in_0_valid | io_in_1_valid | io_in_2_valid); // @[Arbiter.scala 45:78]
  assign io_in_1_ready = ~io_in_0_valid; // @[Arbiter.scala 45:78]
  assign io_in_2_ready = ~(io_in_0_valid | io_in_1_valid); // @[Arbiter.scala 45:78]
  assign io_in_3_ready = ~(io_in_0_valid | io_in_1_valid | io_in_2_valid); // @[Arbiter.scala 45:78]
  assign io_out_valid = ~grant_3 | io_in_3_valid; // @[Arbiter.scala 147:31]
  assign io_out_bits_src_virt_id = io_in_0_valid ? 2'h0 : _GEN_7; // @[Arbiter.scala 138:26 140:19]
  assign io_out_bits_flow_ingress_node = io_in_0_valid ? io_in_0_bits_flow_ingress_node : _GEN_10; // @[Arbiter.scala 138:26 140:19]
  assign io_out_bits_flow_egress_node = io_in_0_valid ? io_in_0_bits_flow_egress_node : _GEN_12; // @[Arbiter.scala 138:26 140:19]
endmodule
module SwitchArbiter(
  input        clock,
  input        reset,
  output       io_in_0_ready,
  input        io_in_0_valid,
  input        io_in_0_bits_vc_sel_2_0,
  input        io_in_0_bits_vc_sel_1_0,
  input        io_in_0_bits_vc_sel_0_0,
  input        io_in_0_bits_tail,
  output       io_in_1_ready,
  input        io_in_1_valid,
  input        io_in_1_bits_vc_sel_2_0,
  input        io_in_1_bits_vc_sel_1_0,
  input        io_in_1_bits_vc_sel_1_1,
  input        io_in_1_bits_vc_sel_0_0,
  input        io_in_1_bits_vc_sel_0_1,
  input        io_in_1_bits_tail,
  output       io_in_2_ready,
  input        io_in_2_valid,
  input        io_in_2_bits_vc_sel_2_0,
  input        io_in_2_bits_vc_sel_1_0,
  input        io_in_2_bits_vc_sel_1_1,
  input        io_in_2_bits_vc_sel_1_2,
  input        io_in_2_bits_vc_sel_0_0,
  input        io_in_2_bits_vc_sel_0_1,
  input        io_in_2_bits_vc_sel_0_2,
  input        io_in_2_bits_tail,
  output       io_in_3_ready,
  input        io_in_3_valid,
  input        io_in_3_bits_vc_sel_2_0,
  input        io_in_3_bits_vc_sel_1_0,
  input        io_in_3_bits_vc_sel_1_1,
  input        io_in_3_bits_vc_sel_1_2,
  input        io_in_3_bits_vc_sel_1_3,
  input        io_in_3_bits_vc_sel_0_0,
  input        io_in_3_bits_vc_sel_0_1,
  input        io_in_3_bits_vc_sel_0_2,
  input        io_in_3_bits_vc_sel_0_3,
  input        io_in_3_bits_tail,
  input        io_out_0_ready,
  output       io_out_0_valid,
  output       io_out_0_bits_vc_sel_2_0,
  output       io_out_0_bits_vc_sel_1_0,
  output       io_out_0_bits_vc_sel_1_1,
  output       io_out_0_bits_vc_sel_1_2,
  output       io_out_0_bits_vc_sel_1_3,
  output       io_out_0_bits_vc_sel_0_0,
  output       io_out_0_bits_vc_sel_0_1,
  output       io_out_0_bits_vc_sel_0_2,
  output       io_out_0_bits_vc_sel_0_3,
  output       io_out_0_bits_tail,
  output [3:0] io_chosen_oh_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] lock_0; // @[SwitchAllocator.scala 24:38]
  wire [3:0] _unassigned_T = {io_in_3_valid,io_in_2_valid,io_in_1_valid,io_in_0_valid}; // @[Cat.scala 33:92]
  wire [3:0] _unassigned_T_1 = ~lock_0; // @[SwitchAllocator.scala 25:54]
  wire [3:0] unassigned = _unassigned_T & _unassigned_T_1; // @[SwitchAllocator.scala 25:52]
  reg [3:0] mask; // @[SwitchAllocator.scala 27:21]
  wire [3:0] _GEN_6 = {{3'd0}, mask == 4'h0}; // @[SwitchAllocator.scala 30:58]
  wire [3:0] _sel_T_1 = unassigned & _GEN_6; // @[SwitchAllocator.scala 30:58]
  wire [7:0] _sel_T_2 = {unassigned,_sel_T_1}; // @[Cat.scala 33:92]
  wire [7:0] _sel_T_11 = _sel_T_2[7] ? 8'h80 : 8'h0; // @[Mux.scala 47:70]
  wire [7:0] _sel_T_12 = _sel_T_2[6] ? 8'h40 : _sel_T_11; // @[Mux.scala 47:70]
  wire [7:0] _sel_T_13 = _sel_T_2[5] ? 8'h20 : _sel_T_12; // @[Mux.scala 47:70]
  wire [7:0] _sel_T_14 = _sel_T_2[4] ? 8'h10 : _sel_T_13; // @[Mux.scala 47:70]
  wire [7:0] _sel_T_15 = _sel_T_2[3] ? 8'h8 : _sel_T_14; // @[Mux.scala 47:70]
  wire [7:0] _sel_T_16 = _sel_T_2[2] ? 8'h4 : _sel_T_15; // @[Mux.scala 47:70]
  wire [7:0] _sel_T_17 = _sel_T_2[1] ? 8'h2 : _sel_T_16; // @[Mux.scala 47:70]
  wire [7:0] sel = _sel_T_2[0] ? 8'h1 : _sel_T_17; // @[Mux.scala 47:70]
  wire [7:0] _GEN_7 = {{4'd0}, sel[7:4]}; // @[SwitchAllocator.scala 32:23]
  wire [7:0] _choices_0_T_1 = sel | _GEN_7; // @[SwitchAllocator.scala 32:23]
  wire [3:0] choices_0 = _choices_0_T_1[3:0]; // @[SwitchAllocator.scala 28:21 32:16]
  wire [3:0] in_tails = {io_in_3_bits_tail,io_in_2_bits_tail,io_in_1_bits_tail,io_in_0_bits_tail}; // @[Cat.scala 33:92]
  wire [3:0] _chosen_T = _unassigned_T & lock_0; // @[SwitchAllocator.scala 42:33]
  wire [3:0] chosen = |_chosen_T ? lock_0 : choices_0; // @[SwitchAllocator.scala 42:21]
  wire [3:0] _io_out_0_valid_T = _unassigned_T & chosen; // @[SwitchAllocator.scala 44:35]
  wire  _T_17 = io_out_0_ready & io_out_0_valid; // @[Decoupled.scala 51:35]
  wire [3:0] _lock_0_T = ~in_tails; // @[SwitchAllocator.scala 53:27]
  wire [3:0] _lock_0_T_1 = chosen & _lock_0_T; // @[SwitchAllocator.scala 53:25]
  wire [3:0] _GEN_8 = {{1'd0}, io_chosen_oh_0[3:1]}; // @[SwitchAllocator.scala 58:71]
  wire [3:0] _mask_T_4 = io_chosen_oh_0 | _GEN_8; // @[SwitchAllocator.scala 58:71]
  wire [3:0] _GEN_9 = {{2'd0}, io_chosen_oh_0[3:2]}; // @[SwitchAllocator.scala 58:71]
  wire [3:0] _mask_T_5 = _mask_T_4 | _GEN_9; // @[SwitchAllocator.scala 58:71]
  wire [3:0] _GEN_10 = {{3'd0}, io_chosen_oh_0[3]}; // @[SwitchAllocator.scala 58:71]
  wire [3:0] _mask_T_6 = _mask_T_5 | _GEN_10; // @[SwitchAllocator.scala 58:71]
  wire [3:0] _mask_T_7 = ~mask; // @[SwitchAllocator.scala 60:17]
  wire [4:0] _mask_T_9 = {mask, 1'h0}; // @[SwitchAllocator.scala 60:43]
  wire [4:0] _mask_T_10 = _mask_T_9 | 5'h1; // @[SwitchAllocator.scala 60:49]
  wire [4:0] _mask_T_11 = _mask_T_7 == 4'h0 ? 5'h0 : _mask_T_10; // @[SwitchAllocator.scala 60:16]
  wire [4:0] _GEN_5 = _T_17 ? {{1'd0}, _mask_T_6} : _mask_T_11; // @[SwitchAllocator.scala 57:27 58:10 60:10]
  wire [4:0] _GEN_11 = reset ? 5'h0 : _GEN_5; // @[SwitchAllocator.scala 27:{21,21}]
  assign io_in_0_ready = chosen[0] & io_out_0_ready; // @[SwitchAllocator.scala 47:23]
  assign io_in_1_ready = chosen[1] & io_out_0_ready; // @[SwitchAllocator.scala 47:23]
  assign io_in_2_ready = chosen[2] & io_out_0_ready; // @[SwitchAllocator.scala 47:23]
  assign io_in_3_ready = chosen[3] & io_out_0_ready; // @[SwitchAllocator.scala 47:23]
  assign io_out_0_valid = |_io_out_0_valid_T; // @[SwitchAllocator.scala 44:45]
  assign io_out_0_bits_vc_sel_2_0 = chosen[0] & io_in_0_bits_vc_sel_2_0 | chosen[1] & io_in_1_bits_vc_sel_2_0 | chosen[2
    ] & io_in_2_bits_vc_sel_2_0 | chosen[3] & io_in_3_bits_vc_sel_2_0; // @[Mux.scala 27:73]
  assign io_out_0_bits_vc_sel_1_0 = chosen[0] & io_in_0_bits_vc_sel_1_0 | chosen[1] & io_in_1_bits_vc_sel_1_0 | chosen[2
    ] & io_in_2_bits_vc_sel_1_0 | chosen[3] & io_in_3_bits_vc_sel_1_0; // @[Mux.scala 27:73]
  assign io_out_0_bits_vc_sel_1_1 = chosen[1] & io_in_1_bits_vc_sel_1_1 | chosen[2] & io_in_2_bits_vc_sel_1_1 | chosen[3
    ] & io_in_3_bits_vc_sel_1_1; // @[Mux.scala 27:73]
  assign io_out_0_bits_vc_sel_1_2 = chosen[2] & io_in_2_bits_vc_sel_1_2 | chosen[3] & io_in_3_bits_vc_sel_1_2; // @[Mux.scala 27:73]
  assign io_out_0_bits_vc_sel_1_3 = chosen[3] & io_in_3_bits_vc_sel_1_3; // @[Mux.scala 27:73]
  assign io_out_0_bits_vc_sel_0_0 = chosen[0] & io_in_0_bits_vc_sel_0_0 | chosen[1] & io_in_1_bits_vc_sel_0_0 | chosen[2
    ] & io_in_2_bits_vc_sel_0_0 | chosen[3] & io_in_3_bits_vc_sel_0_0; // @[Mux.scala 27:73]
  assign io_out_0_bits_vc_sel_0_1 = chosen[1] & io_in_1_bits_vc_sel_0_1 | chosen[2] & io_in_2_bits_vc_sel_0_1 | chosen[3
    ] & io_in_3_bits_vc_sel_0_1; // @[Mux.scala 27:73]
  assign io_out_0_bits_vc_sel_0_2 = chosen[2] & io_in_2_bits_vc_sel_0_2 | chosen[3] & io_in_3_bits_vc_sel_0_2; // @[Mux.scala 27:73]
  assign io_out_0_bits_vc_sel_0_3 = chosen[3] & io_in_3_bits_vc_sel_0_3; // @[Mux.scala 27:73]
  assign io_out_0_bits_tail = chosen[0] & io_in_0_bits_tail | chosen[1] & io_in_1_bits_tail | chosen[2] &
    io_in_2_bits_tail | chosen[3] & io_in_3_bits_tail; // @[Mux.scala 27:73]
  assign io_chosen_oh_0 = |_chosen_T ? lock_0 : choices_0; // @[SwitchAllocator.scala 42:21]
  always @(posedge clock) begin
    if (reset) begin // @[SwitchAllocator.scala 24:38]
      lock_0 <= 4'h0; // @[SwitchAllocator.scala 24:38]
    end else if (_T_17) begin // @[SwitchAllocator.scala 52:29]
      lock_0 <= _lock_0_T_1; // @[SwitchAllocator.scala 53:15]
    end
    mask <= _GEN_11[3:0]; // @[SwitchAllocator.scala 27:{21,21}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lock_0 = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  mask = _RAND_1[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module InputUnit(
  input         clock,
  input         reset,
  output        io_router_req_valid,
  output [1:0]  io_router_req_bits_src_virt_id,
  output [1:0]  io_router_req_bits_flow_ingress_node,
  output [1:0]  io_router_req_bits_flow_egress_node,
  input         io_router_resp_vc_sel_1_0,
  input         io_router_resp_vc_sel_1_1,
  input         io_router_resp_vc_sel_1_2,
  input         io_router_resp_vc_sel_0_0,
  input         io_router_resp_vc_sel_0_1,
  input         io_router_resp_vc_sel_0_2,
  input         io_router_resp_vc_sel_0_3,
  input         io_vcalloc_req_ready,
  output        io_vcalloc_req_valid,
  output        io_vcalloc_req_bits_vc_sel_2_0,
  output        io_vcalloc_req_bits_vc_sel_1_0,
  output        io_vcalloc_req_bits_vc_sel_1_1,
  output        io_vcalloc_req_bits_vc_sel_1_2,
  output        io_vcalloc_req_bits_vc_sel_0_0,
  output        io_vcalloc_req_bits_vc_sel_0_1,
  output        io_vcalloc_req_bits_vc_sel_0_2,
  output        io_vcalloc_req_bits_vc_sel_0_3,
  input         io_vcalloc_resp_vc_sel_2_0,
  input         io_vcalloc_resp_vc_sel_1_0,
  input         io_vcalloc_resp_vc_sel_1_1,
  input         io_vcalloc_resp_vc_sel_1_2,
  input         io_vcalloc_resp_vc_sel_0_0,
  input         io_vcalloc_resp_vc_sel_0_1,
  input         io_vcalloc_resp_vc_sel_0_2,
  input         io_vcalloc_resp_vc_sel_0_3,
  input         io_out_credit_available_2_0,
  input         io_out_credit_available_1_0,
  input         io_out_credit_available_1_1,
  input         io_out_credit_available_1_2,
  input         io_out_credit_available_1_3,
  input         io_out_credit_available_0_0,
  input         io_out_credit_available_0_1,
  input         io_out_credit_available_0_2,
  input         io_out_credit_available_0_3,
  input         io_salloc_req_0_ready,
  output        io_salloc_req_0_valid,
  output        io_salloc_req_0_bits_vc_sel_2_0,
  output        io_salloc_req_0_bits_vc_sel_1_0,
  output        io_salloc_req_0_bits_vc_sel_1_1,
  output        io_salloc_req_0_bits_vc_sel_1_2,
  output        io_salloc_req_0_bits_vc_sel_1_3,
  output        io_salloc_req_0_bits_vc_sel_0_0,
  output        io_salloc_req_0_bits_vc_sel_0_1,
  output        io_salloc_req_0_bits_vc_sel_0_2,
  output        io_salloc_req_0_bits_vc_sel_0_3,
  output        io_salloc_req_0_bits_tail,
  output        io_out_0_valid,
  output        io_out_0_bits_flit_head,
  output        io_out_0_bits_flit_tail,
  output [63:0] io_out_0_bits_flit_payload,
  output [1:0]  io_out_0_bits_flit_flow_ingress_node,
  output [1:0]  io_out_0_bits_flit_flow_egress_node,
  output [1:0]  io_out_0_bits_out_virt_channel,
  output [1:0]  io_debug_va_stall,
  output [1:0]  io_debug_sa_stall,
  input         io_in_flit_0_valid,
  input         io_in_flit_0_bits_head,
  input         io_in_flit_0_bits_tail,
  input  [63:0] io_in_flit_0_bits_payload,
  input  [1:0]  io_in_flit_0_bits_flow_ingress_node,
  input  [1:0]  io_in_flit_0_bits_flow_egress_node,
  input  [1:0]  io_in_flit_0_bits_virt_channel_id,
  output [3:0]  io_in_credit_return,
  output [3:0]  io_in_vc_free
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
`endif // RANDOMIZE_REG_INIT
  wire  input_buffer_clock; // @[InputUnit.scala 180:28]
  wire  input_buffer_reset; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_enq_0_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_enq_0_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_enq_0_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_enq_0_bits_payload; // @[InputUnit.scala 180:28]
  wire [1:0] input_buffer_io_enq_0_bits_virt_channel_id; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_0_ready; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_0_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_0_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_0_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_deq_0_bits_payload; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_ready; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_deq_1_bits_payload; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_ready; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_deq_2_bits_payload; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_3_ready; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_3_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_3_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_3_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_deq_3_bits_payload; // @[InputUnit.scala 180:28]
  wire  route_arbiter_io_in_0_valid; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_0_bits_flow_ingress_node; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_0_bits_flow_egress_node; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_1_ready; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_1_valid; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_1_bits_flow_ingress_node; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_1_bits_flow_egress_node; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_2_ready; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_2_valid; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_2_bits_flow_ingress_node; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_2_bits_flow_egress_node; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_3_ready; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_3_valid; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_3_bits_flow_ingress_node; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_3_bits_flow_egress_node; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_out_valid; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_out_bits_src_virt_id; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_out_bits_flow_ingress_node; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_out_bits_flow_egress_node; // @[InputUnit.scala 186:29]
  wire  salloc_arb_clock; // @[InputUnit.scala 279:26]
  wire  salloc_arb_reset; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_bits_vc_sel_2_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_bits_vc_sel_1_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_bits_tail; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_vc_sel_2_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_vc_sel_1_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_vc_sel_1_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_vc_sel_0_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_tail; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_2_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_1_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_1_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_1_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_0_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_0_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_tail; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_2_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_1_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_1_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_1_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_1_3; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_0_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_0_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_0_3; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_tail; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_2_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_1_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_1_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_1_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_1_3; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_0_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_0_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_0_3; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_tail; // @[InputUnit.scala 279:26]
  wire [3:0] salloc_arb_io_chosen_oh_0; // @[InputUnit.scala 279:26]
  reg [2:0] states_0_g; // @[InputUnit.scala 191:19]
  reg  states_0_vc_sel_2_0; // @[InputUnit.scala 191:19]
  reg  states_0_vc_sel_1_0; // @[InputUnit.scala 191:19]
  reg  states_0_vc_sel_0_0; // @[InputUnit.scala 191:19]
  reg [1:0] states_0_flow_ingress_node; // @[InputUnit.scala 191:19]
  reg [1:0] states_0_flow_egress_node; // @[InputUnit.scala 191:19]
  reg [2:0] states_1_g; // @[InputUnit.scala 191:19]
  reg  states_1_vc_sel_2_0; // @[InputUnit.scala 191:19]
  reg  states_1_vc_sel_1_0; // @[InputUnit.scala 191:19]
  reg  states_1_vc_sel_0_1; // @[InputUnit.scala 191:19]
  reg [1:0] states_1_flow_ingress_node; // @[InputUnit.scala 191:19]
  reg [1:0] states_1_flow_egress_node; // @[InputUnit.scala 191:19]
  reg [2:0] states_2_g; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_2_0; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_1_0; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_1_1; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_0_1; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_0_2; // @[InputUnit.scala 191:19]
  reg [1:0] states_2_flow_ingress_node; // @[InputUnit.scala 191:19]
  reg [1:0] states_2_flow_egress_node; // @[InputUnit.scala 191:19]
  reg [2:0] states_3_g; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_2_0; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_1_0; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_1_1; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_1_2; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_0_1; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_0_2; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_0_3; // @[InputUnit.scala 191:19]
  reg [1:0] states_3_flow_ingress_node; // @[InputUnit.scala 191:19]
  reg [1:0] states_3_flow_egress_node; // @[InputUnit.scala 191:19]
  wire  _T = io_in_flit_0_valid & io_in_flit_0_bits_head; // @[InputUnit.scala 194:32]
  wire  _T_3 = ~reset; // @[InputUnit.scala 196:13]
  wire [2:0] _GEN_1 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? states_1_g : states_0_g; // @[InputUnit.scala 197:{27,27}]
  wire [2:0] _GEN_2 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? states_2_g : _GEN_1; // @[InputUnit.scala 197:{27,27}]
  wire [2:0] _GEN_3 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? states_3_g : _GEN_2; // @[InputUnit.scala 197:{27,27}]
  wire  at_dest = io_in_flit_0_bits_flow_egress_node == 2'h0; // @[InputUnit.scala 198:57]
  wire [2:0] _states_g_T = at_dest ? 3'h2 : 3'h1; // @[InputUnit.scala 199:26]
  wire [2:0] _GEN_4 = 2'h0 == io_in_flit_0_bits_virt_channel_id ? _states_g_T : states_0_g; // @[InputUnit.scala 191:19 199:{20,20}]
  wire [2:0] _GEN_5 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? _states_g_T : states_1_g; // @[InputUnit.scala 191:19 199:{20,20}]
  wire [2:0] _GEN_6 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? _states_g_T : states_2_g; // @[InputUnit.scala 191:19 199:{20,20}]
  wire [2:0] _GEN_7 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? _states_g_T : states_3_g; // @[InputUnit.scala 191:19 199:{20,20}]
  wire  _GEN_8 = 2'h0 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_0_vc_sel_0_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_13 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_1_vc_sel_0_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_14 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_0_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_15 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_0_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_18 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_0_2; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_19 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_0_2; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_23 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_0_3; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_24 = 2'h0 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_0_vc_sel_1_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_25 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_1_vc_sel_1_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_26 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_1_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_27 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_1_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_30 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_1_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_31 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_1_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_35 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_1_2; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_40 = 2'h0 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_0_vc_sel_2_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_41 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_1_vc_sel_2_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_42 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_2_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_43 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_2_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_44 = 2'h0 == io_in_flit_0_bits_virt_channel_id | _GEN_40; // @[InputUnit.scala 203:{44,44}]
  wire  _GEN_45 = 2'h1 == io_in_flit_0_bits_virt_channel_id | _GEN_41; // @[InputUnit.scala 203:{44,44}]
  wire  _GEN_46 = 2'h2 == io_in_flit_0_bits_virt_channel_id | _GEN_42; // @[InputUnit.scala 203:{44,44}]
  wire  _GEN_47 = 2'h3 == io_in_flit_0_bits_virt_channel_id | _GEN_43; // @[InputUnit.scala 203:{44,44}]
  wire [2:0] _GEN_72 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_4 : states_0_g; // @[InputUnit.scala 191:19 194:60]
  wire [2:0] _GEN_73 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_5 : states_1_g; // @[InputUnit.scala 191:19 194:60]
  wire [2:0] _GEN_74 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_6 : states_2_g; // @[InputUnit.scala 191:19 194:60]
  wire [2:0] _GEN_75 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_7 : states_3_g; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_76 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_8 : states_0_vc_sel_0_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_81 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_13 : states_1_vc_sel_0_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_82 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_14 : states_2_vc_sel_0_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_83 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_15 : states_3_vc_sel_0_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_86 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_18 : states_2_vc_sel_0_2; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_87 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_19 : states_3_vc_sel_0_2; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_91 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_23 : states_3_vc_sel_0_3; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_92 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_24 : states_0_vc_sel_1_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_93 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_25 : states_1_vc_sel_1_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_94 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_26 : states_2_vc_sel_1_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_95 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_27 : states_3_vc_sel_1_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_98 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_30 : states_2_vc_sel_1_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_99 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_31 : states_3_vc_sel_1_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_103 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_35 : states_3_vc_sel_1_2; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_108 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_44 : states_0_vc_sel_2_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_109 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_45 : states_1_vc_sel_2_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_110 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_46 : states_2_vc_sel_2_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_111 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_47 : states_3_vc_sel_2_0; // @[InputUnit.scala 191:19 194:60]
  wire  _T_10 = route_arbiter_io_in_0_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_132 = _T_10 ? 3'h2 : _GEN_72; // @[InputUnit.scala 215:{23,29}]
  wire  _T_11 = route_arbiter_io_in_1_ready & route_arbiter_io_in_1_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_133 = _T_11 ? 3'h2 : _GEN_73; // @[InputUnit.scala 215:{23,29}]
  wire  _T_12 = route_arbiter_io_in_2_ready & route_arbiter_io_in_2_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_134 = _T_12 ? 3'h2 : _GEN_74; // @[InputUnit.scala 215:{23,29}]
  wire  _T_13 = route_arbiter_io_in_3_ready & route_arbiter_io_in_3_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_135 = _T_13 ? 3'h2 : _GEN_75; // @[InputUnit.scala 215:{23,29}]
  wire [2:0] _GEN_137 = 2'h1 == io_router_req_bits_src_virt_id ? states_1_g : states_0_g; // @[InputUnit.scala 224:{25,25}]
  wire [2:0] _GEN_138 = 2'h2 == io_router_req_bits_src_virt_id ? states_2_g : _GEN_137; // @[InputUnit.scala 224:{25,25}]
  wire [2:0] _GEN_139 = 2'h3 == io_router_req_bits_src_virt_id ? states_3_g : _GEN_138; // @[InputUnit.scala 224:{25,25}]
  wire [2:0] _GEN_140 = 2'h0 == io_router_req_bits_src_virt_id ? 3'h2 : _GEN_132; // @[InputUnit.scala 225:{18,18}]
  wire [2:0] _GEN_141 = 2'h1 == io_router_req_bits_src_virt_id ? 3'h2 : _GEN_133; // @[InputUnit.scala 225:{18,18}]
  wire [2:0] _GEN_142 = 2'h2 == io_router_req_bits_src_virt_id ? 3'h2 : _GEN_134; // @[InputUnit.scala 225:{18,18}]
  wire [2:0] _GEN_143 = 2'h3 == io_router_req_bits_src_virt_id ? 3'h2 : _GEN_135; // @[InputUnit.scala 225:{18,18}]
  wire  _GEN_144 = 2'h0 == io_router_req_bits_src_virt_id ? 1'h0 : _GEN_108; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_145 = 2'h0 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_0 : _GEN_92; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_149 = 2'h0 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_0 : _GEN_76; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_153 = 2'h1 == io_router_req_bits_src_virt_id ? 1'h0 : _GEN_109; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_154 = 2'h1 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_0 : _GEN_93; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_159 = 2'h1 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_1 : _GEN_81; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_162 = 2'h2 == io_router_req_bits_src_virt_id ? 1'h0 : _GEN_110; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_163 = 2'h2 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_0 : _GEN_94; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_164 = 2'h2 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_1 : _GEN_98; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_168 = 2'h2 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_1 : _GEN_82; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_169 = 2'h2 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_2 : _GEN_86; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_171 = 2'h3 == io_router_req_bits_src_virt_id ? 1'h0 : _GEN_111; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_172 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_0 : _GEN_95; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_173 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_1 : _GEN_99; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_174 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_2 : _GEN_103; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_177 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_1 : _GEN_83; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_178 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_2 : _GEN_87; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_179 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_3 : _GEN_91; // @[InputUnit.scala 227:25 228:26]
  wire [2:0] _GEN_180 = io_router_req_valid ? _GEN_140 : _GEN_132; // @[InputUnit.scala 222:31]
  wire [2:0] _GEN_181 = io_router_req_valid ? _GEN_141 : _GEN_133; // @[InputUnit.scala 222:31]
  wire [2:0] _GEN_182 = io_router_req_valid ? _GEN_142 : _GEN_134; // @[InputUnit.scala 222:31]
  wire [2:0] _GEN_183 = io_router_req_valid ? _GEN_143 : _GEN_135; // @[InputUnit.scala 222:31]
  wire  _GEN_184 = io_router_req_valid ? _GEN_144 : _GEN_108; // @[InputUnit.scala 222:31]
  wire  _GEN_185 = io_router_req_valid ? _GEN_145 : _GEN_92; // @[InputUnit.scala 222:31]
  wire  _GEN_189 = io_router_req_valid ? _GEN_149 : _GEN_76; // @[InputUnit.scala 222:31]
  wire  _GEN_193 = io_router_req_valid ? _GEN_153 : _GEN_109; // @[InputUnit.scala 222:31]
  wire  _GEN_194 = io_router_req_valid ? _GEN_154 : _GEN_93; // @[InputUnit.scala 222:31]
  wire  _GEN_199 = io_router_req_valid ? _GEN_159 : _GEN_81; // @[InputUnit.scala 222:31]
  wire  _GEN_202 = io_router_req_valid ? _GEN_162 : _GEN_110; // @[InputUnit.scala 222:31]
  wire  _GEN_203 = io_router_req_valid ? _GEN_163 : _GEN_94; // @[InputUnit.scala 222:31]
  wire  _GEN_204 = io_router_req_valid ? _GEN_164 : _GEN_98; // @[InputUnit.scala 222:31]
  wire  _GEN_208 = io_router_req_valid ? _GEN_168 : _GEN_82; // @[InputUnit.scala 222:31]
  wire  _GEN_209 = io_router_req_valid ? _GEN_169 : _GEN_86; // @[InputUnit.scala 222:31]
  wire  _GEN_211 = io_router_req_valid ? _GEN_171 : _GEN_111; // @[InputUnit.scala 222:31]
  wire  _GEN_212 = io_router_req_valid ? _GEN_172 : _GEN_95; // @[InputUnit.scala 222:31]
  wire  _GEN_213 = io_router_req_valid ? _GEN_173 : _GEN_99; // @[InputUnit.scala 222:31]
  wire  _GEN_214 = io_router_req_valid ? _GEN_174 : _GEN_103; // @[InputUnit.scala 222:31]
  wire  _GEN_217 = io_router_req_valid ? _GEN_177 : _GEN_83; // @[InputUnit.scala 222:31]
  wire  _GEN_218 = io_router_req_valid ? _GEN_178 : _GEN_87; // @[InputUnit.scala 222:31]
  wire  _GEN_219 = io_router_req_valid ? _GEN_179 : _GEN_91; // @[InputUnit.scala 222:31]
  reg [3:0] mask; // @[InputUnit.scala 233:21]
  wire  vcalloc_vals_1 = states_1_g == 3'h2; // @[InputUnit.scala 249:32]
  wire  vcalloc_vals_0 = states_0_g == 3'h2; // @[InputUnit.scala 249:32]
  wire  vcalloc_vals_3 = states_3_g == 3'h2; // @[InputUnit.scala 249:32]
  wire  vcalloc_vals_2 = states_2_g == 3'h2; // @[InputUnit.scala 249:32]
  wire [3:0] _vcalloc_filter_T = {vcalloc_vals_3,vcalloc_vals_2,vcalloc_vals_1,vcalloc_vals_0}; // @[InputUnit.scala 236:59]
  wire [3:0] _vcalloc_filter_T_2 = ~mask; // @[InputUnit.scala 236:89]
  wire [3:0] _vcalloc_filter_T_3 = _vcalloc_filter_T & _vcalloc_filter_T_2; // @[InputUnit.scala 236:87]
  wire [7:0] _vcalloc_filter_T_4 = {vcalloc_vals_3,vcalloc_vals_2,vcalloc_vals_1,vcalloc_vals_0,_vcalloc_filter_T_3}; // @[Cat.scala 33:92]
  wire [7:0] _vcalloc_filter_T_13 = _vcalloc_filter_T_4[7] ? 8'h80 : 8'h0; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_14 = _vcalloc_filter_T_4[6] ? 8'h40 : _vcalloc_filter_T_13; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_15 = _vcalloc_filter_T_4[5] ? 8'h20 : _vcalloc_filter_T_14; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_16 = _vcalloc_filter_T_4[4] ? 8'h10 : _vcalloc_filter_T_15; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_17 = _vcalloc_filter_T_4[3] ? 8'h8 : _vcalloc_filter_T_16; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_18 = _vcalloc_filter_T_4[2] ? 8'h4 : _vcalloc_filter_T_17; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_19 = _vcalloc_filter_T_4[1] ? 8'h2 : _vcalloc_filter_T_18; // @[Mux.scala 47:70]
  wire [7:0] vcalloc_filter = _vcalloc_filter_T_4[0] ? 8'h1 : _vcalloc_filter_T_19; // @[Mux.scala 47:70]
  wire [3:0] vcalloc_sel = vcalloc_filter[3:0] | vcalloc_filter[7:4]; // @[InputUnit.scala 237:58]
  wire [3:0] _mask_T = 4'h1 << io_router_req_bits_src_virt_id; // @[InputUnit.scala 240:18]
  wire [3:0] _mask_T_2 = _mask_T - 4'h1; // @[InputUnit.scala 240:53]
  wire  _T_26 = vcalloc_vals_0 | vcalloc_vals_1 | vcalloc_vals_2 | vcalloc_vals_3; // @[package.scala 73:59]
  wire [1:0] _mask_T_12 = vcalloc_sel[1] ? 2'h3 : 2'h0; // @[Mux.scala 27:73]
  wire [2:0] _mask_T_13 = vcalloc_sel[2] ? 3'h7 : 3'h0; // @[Mux.scala 27:73]
  wire [3:0] _mask_T_14 = vcalloc_sel[3] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [1:0] _GEN_60 = {{1'd0}, vcalloc_sel[0]}; // @[Mux.scala 27:73]
  wire [1:0] _mask_T_15 = _GEN_60 | _mask_T_12; // @[Mux.scala 27:73]
  wire [2:0] _GEN_61 = {{1'd0}, _mask_T_15}; // @[Mux.scala 27:73]
  wire [2:0] _mask_T_16 = _GEN_61 | _mask_T_13; // @[Mux.scala 27:73]
  wire [3:0] _GEN_62 = {{1'd0}, _mask_T_16}; // @[Mux.scala 27:73]
  wire [3:0] _mask_T_17 = _GEN_62 | _mask_T_14; // @[Mux.scala 27:73]
  wire [2:0] _GEN_222 = vcalloc_vals_0 & vcalloc_sel[0] & io_vcalloc_req_ready ? 3'h3 : _GEN_180; // @[InputUnit.scala 253:{76,82}]
  wire [2:0] _GEN_223 = vcalloc_vals_1 & vcalloc_sel[1] & io_vcalloc_req_ready ? 3'h3 : _GEN_181; // @[InputUnit.scala 253:{76,82}]
  wire [2:0] _GEN_224 = vcalloc_vals_2 & vcalloc_sel[2] & io_vcalloc_req_ready ? 3'h3 : _GEN_182; // @[InputUnit.scala 253:{76,82}]
  wire [2:0] _GEN_225 = vcalloc_vals_3 & vcalloc_sel[3] & io_vcalloc_req_ready ? 3'h3 : _GEN_183; // @[InputUnit.scala 253:{76,82}]
  wire [1:0] _io_debug_va_stall_T = vcalloc_vals_0 + vcalloc_vals_1; // @[Bitwise.scala 51:90]
  wire [1:0] _io_debug_va_stall_T_2 = vcalloc_vals_2 + vcalloc_vals_3; // @[Bitwise.scala 51:90]
  wire [2:0] _io_debug_va_stall_T_4 = _io_debug_va_stall_T + _io_debug_va_stall_T_2; // @[Bitwise.scala 51:90]
  wire [2:0] _GEN_63 = {{2'd0}, io_vcalloc_req_ready}; // @[InputUnit.scala 266:47]
  wire [2:0] _io_debug_va_stall_T_7 = _io_debug_va_stall_T_4 - _GEN_63; // @[InputUnit.scala 266:47]
  wire  _T_39 = io_vcalloc_req_ready & io_vcalloc_req_valid; // @[Decoupled.scala 51:35]
  wire [8:0] _credit_available_T = {states_0_vc_sel_2_0,1'h0,1'h0,1'h0,states_0_vc_sel_1_0,2'h0,1'h0,states_0_vc_sel_0_0
    }; // @[InputUnit.scala 287:40]
  wire [8:0] _credit_available_T_1 = {io_out_credit_available_2_0,io_out_credit_available_1_3,
    io_out_credit_available_1_2,io_out_credit_available_1_1,io_out_credit_available_1_0,io_out_credit_available_0_3,
    io_out_credit_available_0_2,io_out_credit_available_0_1,io_out_credit_available_0_0}; // @[InputUnit.scala 287:73]
  wire [8:0] _credit_available_T_2 = _credit_available_T & _credit_available_T_1; // @[InputUnit.scala 287:47]
  wire  credit_available = _credit_available_T_2 != 9'h0; // @[InputUnit.scala 287:81]
  wire  _T_60 = salloc_arb_io_in_0_ready & salloc_arb_io_in_0_valid; // @[Decoupled.scala 51:35]
  wire [8:0] _credit_available_T_3 = {states_1_vc_sel_2_0,1'h0,1'h0,1'h0,states_1_vc_sel_1_0,2'h0,states_1_vc_sel_0_1,1'h0
    }; // @[InputUnit.scala 287:40]
  wire [8:0] _credit_available_T_5 = _credit_available_T_3 & _credit_available_T_1; // @[InputUnit.scala 287:47]
  wire  credit_available_1 = _credit_available_T_5 != 9'h0; // @[InputUnit.scala 287:81]
  wire  _T_62 = salloc_arb_io_in_1_ready & salloc_arb_io_in_1_valid; // @[Decoupled.scala 51:35]
  wire [8:0] _credit_available_T_6 = {states_2_vc_sel_2_0,1'h0,1'h0,states_2_vc_sel_1_1,states_2_vc_sel_1_0,1'h0,
    states_2_vc_sel_0_2,states_2_vc_sel_0_1,1'h0}; // @[InputUnit.scala 287:40]
  wire [8:0] _credit_available_T_8 = _credit_available_T_6 & _credit_available_T_1; // @[InputUnit.scala 287:47]
  wire  credit_available_2 = _credit_available_T_8 != 9'h0; // @[InputUnit.scala 287:81]
  wire  _T_64 = salloc_arb_io_in_2_ready & salloc_arb_io_in_2_valid; // @[Decoupled.scala 51:35]
  wire [8:0] _credit_available_T_9 = {states_3_vc_sel_2_0,1'h0,states_3_vc_sel_1_2,states_3_vc_sel_1_1,
    states_3_vc_sel_1_0,states_3_vc_sel_0_3,states_3_vc_sel_0_2,states_3_vc_sel_0_1,1'h0}; // @[InputUnit.scala 287:40]
  wire [8:0] _credit_available_T_11 = _credit_available_T_9 & _credit_available_T_1; // @[InputUnit.scala 287:47]
  wire  credit_available_3 = _credit_available_T_11 != 9'h0; // @[InputUnit.scala 287:81]
  wire  _T_66 = salloc_arb_io_in_3_ready & salloc_arb_io_in_3_valid; // @[Decoupled.scala 51:35]
  wire  _io_debug_sa_stall_T_1 = salloc_arb_io_in_0_valid & ~salloc_arb_io_in_0_ready; // @[InputUnit.scala 301:67]
  wire  _io_debug_sa_stall_T_3 = salloc_arb_io_in_1_valid & ~salloc_arb_io_in_1_ready; // @[InputUnit.scala 301:67]
  wire  _io_debug_sa_stall_T_5 = salloc_arb_io_in_2_valid & ~salloc_arb_io_in_2_ready; // @[InputUnit.scala 301:67]
  wire  _io_debug_sa_stall_T_7 = salloc_arb_io_in_3_valid & ~salloc_arb_io_in_3_ready; // @[InputUnit.scala 301:67]
  wire [1:0] _io_debug_sa_stall_T_8 = _io_debug_sa_stall_T_1 + _io_debug_sa_stall_T_3; // @[Bitwise.scala 51:90]
  wire [1:0] _io_debug_sa_stall_T_10 = _io_debug_sa_stall_T_5 + _io_debug_sa_stall_T_7; // @[Bitwise.scala 51:90]
  wire [2:0] _io_debug_sa_stall_T_12 = _io_debug_sa_stall_T_8 + _io_debug_sa_stall_T_10; // @[Bitwise.scala 51:90]
  reg  salloc_outs_0_valid; // @[InputUnit.scala 318:8]
  reg [1:0] salloc_outs_0_out_vid; // @[InputUnit.scala 318:8]
  reg  salloc_outs_0_flit_head; // @[InputUnit.scala 318:8]
  reg  salloc_outs_0_flit_tail; // @[InputUnit.scala 318:8]
  reg [63:0] salloc_outs_0_flit_payload; // @[InputUnit.scala 318:8]
  reg [1:0] salloc_outs_0_flit_flow_ingress_node; // @[InputUnit.scala 318:8]
  reg [1:0] salloc_outs_0_flit_flow_egress_node; // @[InputUnit.scala 318:8]
  wire  _io_in_credit_return_T = salloc_arb_io_out_0_ready & salloc_arb_io_out_0_valid; // @[Decoupled.scala 51:35]
  wire  _io_in_vc_free_T_11 = salloc_arb_io_chosen_oh_0[0] & input_buffer_io_deq_0_bits_tail | salloc_arb_io_chosen_oh_0
    [1] & input_buffer_io_deq_1_bits_tail | salloc_arb_io_chosen_oh_0[2] & input_buffer_io_deq_2_bits_tail |
    salloc_arb_io_chosen_oh_0[3] & input_buffer_io_deq_3_bits_tail; // @[Mux.scala 27:73]
  wire  vc_sel_0_0 = salloc_arb_io_chosen_oh_0[0] & states_0_vc_sel_0_0; // @[Mux.scala 27:73]
  wire  vc_sel_0_1 = salloc_arb_io_chosen_oh_0[1] & states_1_vc_sel_0_1 | salloc_arb_io_chosen_oh_0[2] &
    states_2_vc_sel_0_1 | salloc_arb_io_chosen_oh_0[3] & states_3_vc_sel_0_1; // @[Mux.scala 27:73]
  wire  vc_sel_0_2 = salloc_arb_io_chosen_oh_0[2] & states_2_vc_sel_0_2 | salloc_arb_io_chosen_oh_0[3] &
    states_3_vc_sel_0_2; // @[Mux.scala 27:73]
  wire  vc_sel_0_3 = salloc_arb_io_chosen_oh_0[3] & states_3_vc_sel_0_3; // @[Mux.scala 27:73]
  wire  vc_sel_1_0 = salloc_arb_io_chosen_oh_0[0] & states_0_vc_sel_1_0 | salloc_arb_io_chosen_oh_0[1] &
    states_1_vc_sel_1_0 | salloc_arb_io_chosen_oh_0[2] & states_2_vc_sel_1_0 | salloc_arb_io_chosen_oh_0[3] &
    states_3_vc_sel_1_0; // @[Mux.scala 27:73]
  wire  vc_sel_1_1 = salloc_arb_io_chosen_oh_0[2] & states_2_vc_sel_1_1 | salloc_arb_io_chosen_oh_0[3] &
    states_3_vc_sel_1_1; // @[Mux.scala 27:73]
  wire  vc_sel_1_2 = salloc_arb_io_chosen_oh_0[3] & states_3_vc_sel_1_2; // @[Mux.scala 27:73]
  wire  channel_oh_0 = vc_sel_0_0 | vc_sel_0_1 | vc_sel_0_2 | vc_sel_0_3; // @[InputUnit.scala 334:43]
  wire  channel_oh_1 = vc_sel_1_0 | vc_sel_1_1 | vc_sel_1_2; // @[InputUnit.scala 334:43]
  wire [3:0] _virt_channel_T = {vc_sel_0_3,vc_sel_0_2,vc_sel_0_1,vc_sel_0_0}; // @[OneHot.scala 22:45]
  wire [1:0] virt_channel_hi_1 = _virt_channel_T[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] virt_channel_lo_1 = _virt_channel_T[1:0]; // @[OneHot.scala 31:18]
  wire  _virt_channel_T_1 = |virt_channel_hi_1; // @[OneHot.scala 32:14]
  wire [1:0] _virt_channel_T_2 = virt_channel_hi_1 | virt_channel_lo_1; // @[OneHot.scala 32:28]
  wire [1:0] _virt_channel_T_4 = {_virt_channel_T_1,_virt_channel_T_2[1]}; // @[Cat.scala 33:92]
  wire [3:0] _virt_channel_T_5 = {1'h0,vc_sel_1_2,vc_sel_1_1,vc_sel_1_0}; // @[OneHot.scala 22:45]
  wire [1:0] virt_channel_hi_3 = _virt_channel_T_5[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] virt_channel_lo_3 = _virt_channel_T_5[1:0]; // @[OneHot.scala 31:18]
  wire  _virt_channel_T_6 = |virt_channel_hi_3; // @[OneHot.scala 32:14]
  wire [1:0] _virt_channel_T_7 = virt_channel_hi_3 | virt_channel_lo_3; // @[OneHot.scala 32:28]
  wire [1:0] _virt_channel_T_9 = {_virt_channel_T_6,_virt_channel_T_7[1]}; // @[Cat.scala 33:92]
  wire [1:0] _virt_channel_T_10 = channel_oh_0 ? _virt_channel_T_4 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _virt_channel_T_11 = channel_oh_1 ? _virt_channel_T_9 : 2'h0; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_4 = salloc_arb_io_chosen_oh_0[0] ? input_buffer_io_deq_0_bits_payload : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_5 = salloc_arb_io_chosen_oh_0[1] ? input_buffer_io_deq_1_bits_payload : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_6 = salloc_arb_io_chosen_oh_0[2] ? input_buffer_io_deq_2_bits_payload : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_7 = salloc_arb_io_chosen_oh_0[3] ? input_buffer_io_deq_3_bits_payload : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_8 = _salloc_outs_0_flit_payload_T_4 | _salloc_outs_0_flit_payload_T_5; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_9 = _salloc_outs_0_flit_payload_T_8 | _salloc_outs_0_flit_payload_T_6; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_11 = salloc_arb_io_chosen_oh_0[0] ? states_0_flow_egress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_12 = salloc_arb_io_chosen_oh_0[1] ? states_1_flow_egress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_13 = salloc_arb_io_chosen_oh_0[2] ? states_2_flow_egress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_14 = salloc_arb_io_chosen_oh_0[3] ? states_3_flow_egress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_15 = _salloc_outs_0_flit_flow_T_11 | _salloc_outs_0_flit_flow_T_12; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_16 = _salloc_outs_0_flit_flow_T_15 | _salloc_outs_0_flit_flow_T_13; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_25 = salloc_arb_io_chosen_oh_0[0] ? states_0_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_26 = salloc_arb_io_chosen_oh_0[1] ? states_1_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_27 = salloc_arb_io_chosen_oh_0[2] ? states_2_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_28 = salloc_arb_io_chosen_oh_0[3] ? states_3_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_29 = _salloc_outs_0_flit_flow_T_25 | _salloc_outs_0_flit_flow_T_26; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_30 = _salloc_outs_0_flit_flow_T_29 | _salloc_outs_0_flit_flow_T_27; // @[Mux.scala 27:73]
  InputBuffer input_buffer ( // @[InputUnit.scala 180:28]
    .clock(input_buffer_clock),
    .reset(input_buffer_reset),
    .io_enq_0_valid(input_buffer_io_enq_0_valid),
    .io_enq_0_bits_head(input_buffer_io_enq_0_bits_head),
    .io_enq_0_bits_tail(input_buffer_io_enq_0_bits_tail),
    .io_enq_0_bits_payload(input_buffer_io_enq_0_bits_payload),
    .io_enq_0_bits_virt_channel_id(input_buffer_io_enq_0_bits_virt_channel_id),
    .io_deq_0_ready(input_buffer_io_deq_0_ready),
    .io_deq_0_valid(input_buffer_io_deq_0_valid),
    .io_deq_0_bits_head(input_buffer_io_deq_0_bits_head),
    .io_deq_0_bits_tail(input_buffer_io_deq_0_bits_tail),
    .io_deq_0_bits_payload(input_buffer_io_deq_0_bits_payload),
    .io_deq_1_ready(input_buffer_io_deq_1_ready),
    .io_deq_1_valid(input_buffer_io_deq_1_valid),
    .io_deq_1_bits_head(input_buffer_io_deq_1_bits_head),
    .io_deq_1_bits_tail(input_buffer_io_deq_1_bits_tail),
    .io_deq_1_bits_payload(input_buffer_io_deq_1_bits_payload),
    .io_deq_2_ready(input_buffer_io_deq_2_ready),
    .io_deq_2_valid(input_buffer_io_deq_2_valid),
    .io_deq_2_bits_head(input_buffer_io_deq_2_bits_head),
    .io_deq_2_bits_tail(input_buffer_io_deq_2_bits_tail),
    .io_deq_2_bits_payload(input_buffer_io_deq_2_bits_payload),
    .io_deq_3_ready(input_buffer_io_deq_3_ready),
    .io_deq_3_valid(input_buffer_io_deq_3_valid),
    .io_deq_3_bits_head(input_buffer_io_deq_3_bits_head),
    .io_deq_3_bits_tail(input_buffer_io_deq_3_bits_tail),
    .io_deq_3_bits_payload(input_buffer_io_deq_3_bits_payload)
  );
  Arbiter route_arbiter ( // @[InputUnit.scala 186:29]
    .io_in_0_valid(route_arbiter_io_in_0_valid),
    .io_in_0_bits_flow_ingress_node(route_arbiter_io_in_0_bits_flow_ingress_node),
    .io_in_0_bits_flow_egress_node(route_arbiter_io_in_0_bits_flow_egress_node),
    .io_in_1_ready(route_arbiter_io_in_1_ready),
    .io_in_1_valid(route_arbiter_io_in_1_valid),
    .io_in_1_bits_flow_ingress_node(route_arbiter_io_in_1_bits_flow_ingress_node),
    .io_in_1_bits_flow_egress_node(route_arbiter_io_in_1_bits_flow_egress_node),
    .io_in_2_ready(route_arbiter_io_in_2_ready),
    .io_in_2_valid(route_arbiter_io_in_2_valid),
    .io_in_2_bits_flow_ingress_node(route_arbiter_io_in_2_bits_flow_ingress_node),
    .io_in_2_bits_flow_egress_node(route_arbiter_io_in_2_bits_flow_egress_node),
    .io_in_3_ready(route_arbiter_io_in_3_ready),
    .io_in_3_valid(route_arbiter_io_in_3_valid),
    .io_in_3_bits_flow_ingress_node(route_arbiter_io_in_3_bits_flow_ingress_node),
    .io_in_3_bits_flow_egress_node(route_arbiter_io_in_3_bits_flow_egress_node),
    .io_out_valid(route_arbiter_io_out_valid),
    .io_out_bits_src_virt_id(route_arbiter_io_out_bits_src_virt_id),
    .io_out_bits_flow_ingress_node(route_arbiter_io_out_bits_flow_ingress_node),
    .io_out_bits_flow_egress_node(route_arbiter_io_out_bits_flow_egress_node)
  );
  SwitchArbiter salloc_arb ( // @[InputUnit.scala 279:26]
    .clock(salloc_arb_clock),
    .reset(salloc_arb_reset),
    .io_in_0_ready(salloc_arb_io_in_0_ready),
    .io_in_0_valid(salloc_arb_io_in_0_valid),
    .io_in_0_bits_vc_sel_2_0(salloc_arb_io_in_0_bits_vc_sel_2_0),
    .io_in_0_bits_vc_sel_1_0(salloc_arb_io_in_0_bits_vc_sel_1_0),
    .io_in_0_bits_vc_sel_0_0(salloc_arb_io_in_0_bits_vc_sel_0_0),
    .io_in_0_bits_tail(salloc_arb_io_in_0_bits_tail),
    .io_in_1_ready(salloc_arb_io_in_1_ready),
    .io_in_1_valid(salloc_arb_io_in_1_valid),
    .io_in_1_bits_vc_sel_2_0(salloc_arb_io_in_1_bits_vc_sel_2_0),
    .io_in_1_bits_vc_sel_1_0(salloc_arb_io_in_1_bits_vc_sel_1_0),
    .io_in_1_bits_vc_sel_1_1(salloc_arb_io_in_1_bits_vc_sel_1_1),
    .io_in_1_bits_vc_sel_0_0(salloc_arb_io_in_1_bits_vc_sel_0_0),
    .io_in_1_bits_vc_sel_0_1(salloc_arb_io_in_1_bits_vc_sel_0_1),
    .io_in_1_bits_tail(salloc_arb_io_in_1_bits_tail),
    .io_in_2_ready(salloc_arb_io_in_2_ready),
    .io_in_2_valid(salloc_arb_io_in_2_valid),
    .io_in_2_bits_vc_sel_2_0(salloc_arb_io_in_2_bits_vc_sel_2_0),
    .io_in_2_bits_vc_sel_1_0(salloc_arb_io_in_2_bits_vc_sel_1_0),
    .io_in_2_bits_vc_sel_1_1(salloc_arb_io_in_2_bits_vc_sel_1_1),
    .io_in_2_bits_vc_sel_1_2(salloc_arb_io_in_2_bits_vc_sel_1_2),
    .io_in_2_bits_vc_sel_0_0(salloc_arb_io_in_2_bits_vc_sel_0_0),
    .io_in_2_bits_vc_sel_0_1(salloc_arb_io_in_2_bits_vc_sel_0_1),
    .io_in_2_bits_vc_sel_0_2(salloc_arb_io_in_2_bits_vc_sel_0_2),
    .io_in_2_bits_tail(salloc_arb_io_in_2_bits_tail),
    .io_in_3_ready(salloc_arb_io_in_3_ready),
    .io_in_3_valid(salloc_arb_io_in_3_valid),
    .io_in_3_bits_vc_sel_2_0(salloc_arb_io_in_3_bits_vc_sel_2_0),
    .io_in_3_bits_vc_sel_1_0(salloc_arb_io_in_3_bits_vc_sel_1_0),
    .io_in_3_bits_vc_sel_1_1(salloc_arb_io_in_3_bits_vc_sel_1_1),
    .io_in_3_bits_vc_sel_1_2(salloc_arb_io_in_3_bits_vc_sel_1_2),
    .io_in_3_bits_vc_sel_1_3(salloc_arb_io_in_3_bits_vc_sel_1_3),
    .io_in_3_bits_vc_sel_0_0(salloc_arb_io_in_3_bits_vc_sel_0_0),
    .io_in_3_bits_vc_sel_0_1(salloc_arb_io_in_3_bits_vc_sel_0_1),
    .io_in_3_bits_vc_sel_0_2(salloc_arb_io_in_3_bits_vc_sel_0_2),
    .io_in_3_bits_vc_sel_0_3(salloc_arb_io_in_3_bits_vc_sel_0_3),
    .io_in_3_bits_tail(salloc_arb_io_in_3_bits_tail),
    .io_out_0_ready(salloc_arb_io_out_0_ready),
    .io_out_0_valid(salloc_arb_io_out_0_valid),
    .io_out_0_bits_vc_sel_2_0(salloc_arb_io_out_0_bits_vc_sel_2_0),
    .io_out_0_bits_vc_sel_1_0(salloc_arb_io_out_0_bits_vc_sel_1_0),
    .io_out_0_bits_vc_sel_1_1(salloc_arb_io_out_0_bits_vc_sel_1_1),
    .io_out_0_bits_vc_sel_1_2(salloc_arb_io_out_0_bits_vc_sel_1_2),
    .io_out_0_bits_vc_sel_1_3(salloc_arb_io_out_0_bits_vc_sel_1_3),
    .io_out_0_bits_vc_sel_0_0(salloc_arb_io_out_0_bits_vc_sel_0_0),
    .io_out_0_bits_vc_sel_0_1(salloc_arb_io_out_0_bits_vc_sel_0_1),
    .io_out_0_bits_vc_sel_0_2(salloc_arb_io_out_0_bits_vc_sel_0_2),
    .io_out_0_bits_vc_sel_0_3(salloc_arb_io_out_0_bits_vc_sel_0_3),
    .io_out_0_bits_tail(salloc_arb_io_out_0_bits_tail),
    .io_chosen_oh_0(salloc_arb_io_chosen_oh_0)
  );
  assign io_router_req_valid = route_arbiter_io_out_valid; // @[InputUnit.scala 189:17]
  assign io_router_req_bits_src_virt_id = route_arbiter_io_out_bits_src_virt_id; // @[InputUnit.scala 189:17]
  assign io_router_req_bits_flow_ingress_node = route_arbiter_io_out_bits_flow_ingress_node; // @[InputUnit.scala 189:17]
  assign io_router_req_bits_flow_egress_node = route_arbiter_io_out_bits_flow_egress_node; // @[InputUnit.scala 189:17]
  assign io_vcalloc_req_valid = vcalloc_vals_0 | vcalloc_vals_1 | vcalloc_vals_2 | vcalloc_vals_3; // @[package.scala 73:59]
  assign io_vcalloc_req_bits_vc_sel_2_0 = vcalloc_sel[0] & states_0_vc_sel_2_0 | vcalloc_sel[1] & states_1_vc_sel_2_0 |
    vcalloc_sel[2] & states_2_vc_sel_2_0 | vcalloc_sel[3] & states_3_vc_sel_2_0; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_1_0 = vcalloc_sel[0] & states_0_vc_sel_1_0 | vcalloc_sel[1] & states_1_vc_sel_1_0 |
    vcalloc_sel[2] & states_2_vc_sel_1_0 | vcalloc_sel[3] & states_3_vc_sel_1_0; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_1_1 = vcalloc_sel[2] & states_2_vc_sel_1_1 | vcalloc_sel[3] & states_3_vc_sel_1_1; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_1_2 = vcalloc_sel[3] & states_3_vc_sel_1_2; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_0_0 = vcalloc_sel[0] & states_0_vc_sel_0_0; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_0_1 = vcalloc_sel[1] & states_1_vc_sel_0_1 | vcalloc_sel[2] & states_2_vc_sel_0_1 |
    vcalloc_sel[3] & states_3_vc_sel_0_1; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_0_2 = vcalloc_sel[2] & states_2_vc_sel_0_2 | vcalloc_sel[3] & states_3_vc_sel_0_2; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_0_3 = vcalloc_sel[3] & states_3_vc_sel_0_3; // @[Mux.scala 27:73]
  assign io_salloc_req_0_valid = salloc_arb_io_out_0_valid; // @[InputUnit.scala 302:17 303:19 305:35]
  assign io_salloc_req_0_bits_vc_sel_2_0 = salloc_arb_io_out_0_bits_vc_sel_2_0; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_1_0 = salloc_arb_io_out_0_bits_vc_sel_1_0; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_1_1 = salloc_arb_io_out_0_bits_vc_sel_1_1; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_1_2 = salloc_arb_io_out_0_bits_vc_sel_1_2; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_1_3 = salloc_arb_io_out_0_bits_vc_sel_1_3; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_0_0 = salloc_arb_io_out_0_bits_vc_sel_0_0; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_0_1 = salloc_arb_io_out_0_bits_vc_sel_0_1; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_0_2 = salloc_arb_io_out_0_bits_vc_sel_0_2; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_0_3 = salloc_arb_io_out_0_bits_vc_sel_0_3; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_tail = salloc_arb_io_out_0_bits_tail; // @[InputUnit.scala 302:17]
  assign io_out_0_valid = salloc_outs_0_valid; // @[InputUnit.scala 349:21]
  assign io_out_0_bits_flit_head = salloc_outs_0_flit_head; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_flit_tail = salloc_outs_0_flit_tail; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_flit_payload = salloc_outs_0_flit_payload; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_flit_flow_ingress_node = salloc_outs_0_flit_flow_ingress_node; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_flit_flow_egress_node = salloc_outs_0_flit_flow_egress_node; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_out_virt_channel = salloc_outs_0_out_vid; // @[InputUnit.scala 351:37]
  assign io_debug_va_stall = _io_debug_va_stall_T_7[1:0]; // @[InputUnit.scala 266:21]
  assign io_debug_sa_stall = _io_debug_sa_stall_T_12[1:0]; // @[InputUnit.scala 301:21]
  assign io_in_credit_return = _io_in_credit_return_T ? salloc_arb_io_chosen_oh_0 : 4'h0; // @[InputUnit.scala 322:8]
  assign io_in_vc_free = _io_in_credit_return_T & _io_in_vc_free_T_11 ? salloc_arb_io_chosen_oh_0 : 4'h0; // @[InputUnit.scala 325:8]
  assign input_buffer_clock = clock;
  assign input_buffer_reset = reset;
  assign input_buffer_io_enq_0_valid = io_in_flit_0_valid; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_head = io_in_flit_0_bits_head; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_tail = io_in_flit_0_bits_tail; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_payload = io_in_flit_0_bits_payload; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_virt_channel_id = io_in_flit_0_bits_virt_channel_id; // @[InputUnit.scala 182:28]
  assign input_buffer_io_deq_0_ready = salloc_arb_io_in_0_ready; // @[InputUnit.scala 295:36]
  assign input_buffer_io_deq_1_ready = salloc_arb_io_in_1_ready; // @[InputUnit.scala 295:36]
  assign input_buffer_io_deq_2_ready = salloc_arb_io_in_2_ready; // @[InputUnit.scala 295:36]
  assign input_buffer_io_deq_3_ready = salloc_arb_io_in_3_ready; // @[InputUnit.scala 295:36]
  assign route_arbiter_io_in_0_valid = states_0_g == 3'h1; // @[InputUnit.scala 212:22]
  assign route_arbiter_io_in_0_bits_flow_ingress_node = states_0_flow_ingress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_0_bits_flow_egress_node = states_0_flow_egress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_1_valid = states_1_g == 3'h1; // @[InputUnit.scala 212:22]
  assign route_arbiter_io_in_1_bits_flow_ingress_node = states_1_flow_ingress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_1_bits_flow_egress_node = states_1_flow_egress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_2_valid = states_2_g == 3'h1; // @[InputUnit.scala 212:22]
  assign route_arbiter_io_in_2_bits_flow_ingress_node = states_2_flow_ingress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_2_bits_flow_egress_node = states_2_flow_egress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_3_valid = states_3_g == 3'h1; // @[InputUnit.scala 212:22]
  assign route_arbiter_io_in_3_bits_flow_ingress_node = states_3_flow_ingress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_3_bits_flow_egress_node = states_3_flow_egress_node; // @[InputUnit.scala 213:19]
  assign salloc_arb_clock = clock;
  assign salloc_arb_reset = reset;
  assign salloc_arb_io_in_0_valid = states_0_g == 3'h3 & credit_available & input_buffer_io_deq_0_valid; // @[InputUnit.scala 288:50]
  assign salloc_arb_io_in_0_bits_vc_sel_2_0 = states_0_vc_sel_2_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_0_bits_vc_sel_1_0 = states_0_vc_sel_1_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_0_bits_vc_sel_0_0 = states_0_vc_sel_0_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_0_bits_tail = input_buffer_io_deq_0_bits_tail; // @[InputUnit.scala 291:19]
  assign salloc_arb_io_in_1_valid = states_1_g == 3'h3 & credit_available_1 & input_buffer_io_deq_1_valid; // @[InputUnit.scala 288:50]
  assign salloc_arb_io_in_1_bits_vc_sel_2_0 = states_1_vc_sel_2_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_1_bits_vc_sel_1_0 = states_1_vc_sel_1_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_1_bits_vc_sel_1_1 = 1'h0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_1_bits_vc_sel_0_0 = 1'h0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_1_bits_vc_sel_0_1 = states_1_vc_sel_0_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_1_bits_tail = input_buffer_io_deq_1_bits_tail; // @[InputUnit.scala 291:19]
  assign salloc_arb_io_in_2_valid = states_2_g == 3'h3 & credit_available_2 & input_buffer_io_deq_2_valid; // @[InputUnit.scala 288:50]
  assign salloc_arb_io_in_2_bits_vc_sel_2_0 = states_2_vc_sel_2_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_1_0 = states_2_vc_sel_1_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_1_1 = states_2_vc_sel_1_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_1_2 = 1'h0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_0_0 = 1'h0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_0_1 = states_2_vc_sel_0_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_0_2 = states_2_vc_sel_0_2; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_tail = input_buffer_io_deq_2_bits_tail; // @[InputUnit.scala 291:19]
  assign salloc_arb_io_in_3_valid = states_3_g == 3'h3 & credit_available_3 & input_buffer_io_deq_3_valid; // @[InputUnit.scala 288:50]
  assign salloc_arb_io_in_3_bits_vc_sel_2_0 = states_3_vc_sel_2_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_1_0 = states_3_vc_sel_1_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_1_1 = states_3_vc_sel_1_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_1_2 = states_3_vc_sel_1_2; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_1_3 = 1'h0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_0_0 = 1'h0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_0_1 = states_3_vc_sel_0_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_0_2 = states_3_vc_sel_0_2; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_0_3 = states_3_vc_sel_0_3; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_tail = input_buffer_io_deq_3_bits_tail; // @[InputUnit.scala 291:19]
  assign salloc_arb_io_out_0_ready = io_salloc_req_0_ready; // @[InputUnit.scala 302:17 303:19 304:39]
  always @(posedge clock) begin
    if (reset) begin // @[InputUnit.scala 377:23]
      states_0_g <= 3'h0; // @[InputUnit.scala 378:24]
    end else if (_T_60 & input_buffer_io_deq_0_bits_tail) begin // @[InputUnit.scala 292:35]
      states_0_g <= 3'h0; // @[InputUnit.scala 293:13]
    end else if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[0]) begin // @[InputUnit.scala 270:29]
        states_0_g <= 3'h3; // @[InputUnit.scala 272:21]
      end else begin
        states_0_g <= _GEN_222;
      end
    end else begin
      states_0_g <= _GEN_222;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[0]) begin // @[InputUnit.scala 270:29]
        states_0_vc_sel_2_0 <= io_vcalloc_resp_vc_sel_2_0; // @[InputUnit.scala 271:26]
      end else begin
        states_0_vc_sel_2_0 <= _GEN_184;
      end
    end else begin
      states_0_vc_sel_2_0 <= _GEN_184;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[0]) begin // @[InputUnit.scala 270:29]
        states_0_vc_sel_1_0 <= io_vcalloc_resp_vc_sel_1_0; // @[InputUnit.scala 271:26]
      end else begin
        states_0_vc_sel_1_0 <= _GEN_185;
      end
    end else begin
      states_0_vc_sel_1_0 <= _GEN_185;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[0]) begin // @[InputUnit.scala 270:29]
        states_0_vc_sel_0_0 <= io_vcalloc_resp_vc_sel_0_0; // @[InputUnit.scala 271:26]
      end else begin
        states_0_vc_sel_0_0 <= _GEN_189;
      end
    end else begin
      states_0_vc_sel_0_0 <= _GEN_189;
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h0 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_0_flow_ingress_node <= io_in_flit_0_bits_flow_ingress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h0 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_0_flow_egress_node <= io_in_flit_0_bits_flow_egress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (reset) begin // @[InputUnit.scala 377:23]
      states_1_g <= 3'h0; // @[InputUnit.scala 378:24]
    end else if (_T_62 & input_buffer_io_deq_1_bits_tail) begin // @[InputUnit.scala 292:35]
      states_1_g <= 3'h0; // @[InputUnit.scala 293:13]
    end else if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_g <= 3'h3; // @[InputUnit.scala 272:21]
      end else begin
        states_1_g <= _GEN_223;
      end
    end else begin
      states_1_g <= _GEN_223;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_vc_sel_2_0 <= io_vcalloc_resp_vc_sel_2_0; // @[InputUnit.scala 271:26]
      end else begin
        states_1_vc_sel_2_0 <= _GEN_193;
      end
    end else begin
      states_1_vc_sel_2_0 <= _GEN_193;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_vc_sel_1_0 <= io_vcalloc_resp_vc_sel_1_0; // @[InputUnit.scala 271:26]
      end else begin
        states_1_vc_sel_1_0 <= _GEN_194;
      end
    end else begin
      states_1_vc_sel_1_0 <= _GEN_194;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_vc_sel_0_1 <= io_vcalloc_resp_vc_sel_0_1; // @[InputUnit.scala 271:26]
      end else begin
        states_1_vc_sel_0_1 <= _GEN_199;
      end
    end else begin
      states_1_vc_sel_0_1 <= _GEN_199;
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h1 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_1_flow_ingress_node <= io_in_flit_0_bits_flow_ingress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h1 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_1_flow_egress_node <= io_in_flit_0_bits_flow_egress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (reset) begin // @[InputUnit.scala 377:23]
      states_2_g <= 3'h0; // @[InputUnit.scala 378:24]
    end else if (_T_64 & input_buffer_io_deq_2_bits_tail) begin // @[InputUnit.scala 292:35]
      states_2_g <= 3'h0; // @[InputUnit.scala 293:13]
    end else if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_g <= 3'h3; // @[InputUnit.scala 272:21]
      end else begin
        states_2_g <= _GEN_224;
      end
    end else begin
      states_2_g <= _GEN_224;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_2_0 <= io_vcalloc_resp_vc_sel_2_0; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_2_0 <= _GEN_202;
      end
    end else begin
      states_2_vc_sel_2_0 <= _GEN_202;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_1_0 <= io_vcalloc_resp_vc_sel_1_0; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_1_0 <= _GEN_203;
      end
    end else begin
      states_2_vc_sel_1_0 <= _GEN_203;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_1_1 <= io_vcalloc_resp_vc_sel_1_1; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_1_1 <= _GEN_204;
      end
    end else begin
      states_2_vc_sel_1_1 <= _GEN_204;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_0_1 <= io_vcalloc_resp_vc_sel_0_1; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_0_1 <= _GEN_208;
      end
    end else begin
      states_2_vc_sel_0_1 <= _GEN_208;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_0_2 <= io_vcalloc_resp_vc_sel_0_2; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_0_2 <= _GEN_209;
      end
    end else begin
      states_2_vc_sel_0_2 <= _GEN_209;
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h2 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_2_flow_ingress_node <= io_in_flit_0_bits_flow_ingress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h2 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_2_flow_egress_node <= io_in_flit_0_bits_flow_egress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (reset) begin // @[InputUnit.scala 377:23]
      states_3_g <= 3'h0; // @[InputUnit.scala 378:24]
    end else if (_T_66 & input_buffer_io_deq_3_bits_tail) begin // @[InputUnit.scala 292:35]
      states_3_g <= 3'h0; // @[InputUnit.scala 293:13]
    end else if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_g <= 3'h3; // @[InputUnit.scala 272:21]
      end else begin
        states_3_g <= _GEN_225;
      end
    end else begin
      states_3_g <= _GEN_225;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_2_0 <= io_vcalloc_resp_vc_sel_2_0; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_2_0 <= _GEN_211;
      end
    end else begin
      states_3_vc_sel_2_0 <= _GEN_211;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_1_0 <= io_vcalloc_resp_vc_sel_1_0; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_1_0 <= _GEN_212;
      end
    end else begin
      states_3_vc_sel_1_0 <= _GEN_212;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_1_1 <= io_vcalloc_resp_vc_sel_1_1; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_1_1 <= _GEN_213;
      end
    end else begin
      states_3_vc_sel_1_1 <= _GEN_213;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_1_2 <= io_vcalloc_resp_vc_sel_1_2; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_1_2 <= _GEN_214;
      end
    end else begin
      states_3_vc_sel_1_2 <= _GEN_214;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_0_1 <= io_vcalloc_resp_vc_sel_0_1; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_0_1 <= _GEN_217;
      end
    end else begin
      states_3_vc_sel_0_1 <= _GEN_217;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_0_2 <= io_vcalloc_resp_vc_sel_0_2; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_0_2 <= _GEN_218;
      end
    end else begin
      states_3_vc_sel_0_2 <= _GEN_218;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_0_3 <= io_vcalloc_resp_vc_sel_0_3; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_0_3 <= _GEN_219;
      end
    end else begin
      states_3_vc_sel_0_3 <= _GEN_219;
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h3 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_3_flow_ingress_node <= io_in_flit_0_bits_flow_ingress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h3 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_3_flow_egress_node <= io_in_flit_0_bits_flow_egress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (reset) begin // @[InputUnit.scala 233:21]
      mask <= 4'h0; // @[InputUnit.scala 233:21]
    end else if (io_router_req_valid) begin // @[InputUnit.scala 239:31]
      mask <= _mask_T_2; // @[InputUnit.scala 240:10]
    end else if (_T_26) begin // @[InputUnit.scala 241:34]
      mask <= _mask_T_17; // @[InputUnit.scala 242:10]
    end
    salloc_outs_0_valid <= salloc_arb_io_out_0_ready & salloc_arb_io_out_0_valid; // @[Decoupled.scala 51:35]
    salloc_outs_0_out_vid <= _virt_channel_T_10 | _virt_channel_T_11; // @[Mux.scala 27:73]
    salloc_outs_0_flit_head <= salloc_arb_io_chosen_oh_0[0] & input_buffer_io_deq_0_bits_head |
      salloc_arb_io_chosen_oh_0[1] & input_buffer_io_deq_1_bits_head | salloc_arb_io_chosen_oh_0[2] &
      input_buffer_io_deq_2_bits_head | salloc_arb_io_chosen_oh_0[3] & input_buffer_io_deq_3_bits_head; // @[Mux.scala 27:73]
    salloc_outs_0_flit_tail <= salloc_arb_io_chosen_oh_0[0] & input_buffer_io_deq_0_bits_tail |
      salloc_arb_io_chosen_oh_0[1] & input_buffer_io_deq_1_bits_tail | salloc_arb_io_chosen_oh_0[2] &
      input_buffer_io_deq_2_bits_tail | salloc_arb_io_chosen_oh_0[3] & input_buffer_io_deq_3_bits_tail; // @[Mux.scala 27:73]
    salloc_outs_0_flit_payload <= _salloc_outs_0_flit_payload_T_9 | _salloc_outs_0_flit_payload_T_7; // @[Mux.scala 27:73]
    salloc_outs_0_flit_flow_ingress_node <= _salloc_outs_0_flit_flow_T_30 | _salloc_outs_0_flit_flow_T_28; // @[Mux.scala 27:73]
    salloc_outs_0_flit_flow_egress_node <= _salloc_outs_0_flit_flow_T_16 | _salloc_outs_0_flit_flow_T_14; // @[Mux.scala 27:73]
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T & _T_3 & ~(_GEN_3 == 3'h0)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:197 assert(states(id).g === g_i)\n"); // @[InputUnit.scala 197:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_router_req_valid & _T_3 & ~(_GEN_139 == 3'h1)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:224 assert(states(id).g === g_r)\n"); // @[InputUnit.scala 224:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_39 & vcalloc_sel[0] & _T_3 & ~vcalloc_vals_0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:274 assert(states(i).g === g_v)\n"); // @[InputUnit.scala 274:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_39 & vcalloc_sel[1] & _T_3 & ~vcalloc_vals_1) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:274 assert(states(i).g === g_v)\n"); // @[InputUnit.scala 274:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_39 & vcalloc_sel[2] & _T_3 & ~vcalloc_vals_2) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:274 assert(states(i).g === g_v)\n"); // @[InputUnit.scala 274:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_39 & vcalloc_sel[3] & _T_3 & ~vcalloc_vals_3) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:274 assert(states(i).g === g_v)\n"); // @[InputUnit.scala 274:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  states_0_g = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  states_0_vc_sel_2_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  states_0_vc_sel_1_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  states_0_vc_sel_0_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  states_0_flow_ingress_node = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  states_0_flow_egress_node = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  states_1_g = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  states_1_vc_sel_2_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  states_1_vc_sel_1_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  states_1_vc_sel_0_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  states_1_flow_ingress_node = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  states_1_flow_egress_node = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  states_2_g = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  states_2_vc_sel_2_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  states_2_vc_sel_1_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  states_2_vc_sel_1_1 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  states_2_vc_sel_0_1 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  states_2_vc_sel_0_2 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  states_2_flow_ingress_node = _RAND_18[1:0];
  _RAND_19 = {1{`RANDOM}};
  states_2_flow_egress_node = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  states_3_g = _RAND_20[2:0];
  _RAND_21 = {1{`RANDOM}};
  states_3_vc_sel_2_0 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  states_3_vc_sel_1_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  states_3_vc_sel_1_1 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  states_3_vc_sel_1_2 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  states_3_vc_sel_0_1 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  states_3_vc_sel_0_2 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  states_3_vc_sel_0_3 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  states_3_flow_ingress_node = _RAND_28[1:0];
  _RAND_29 = {1{`RANDOM}};
  states_3_flow_egress_node = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  mask = _RAND_30[3:0];
  _RAND_31 = {1{`RANDOM}};
  salloc_outs_0_valid = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  salloc_outs_0_out_vid = _RAND_32[1:0];
  _RAND_33 = {1{`RANDOM}};
  salloc_outs_0_flit_head = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  salloc_outs_0_flit_tail = _RAND_34[0:0];
  _RAND_35 = {2{`RANDOM}};
  salloc_outs_0_flit_payload = _RAND_35[63:0];
  _RAND_36 = {1{`RANDOM}};
  salloc_outs_0_flit_flow_ingress_node = _RAND_36[1:0];
  _RAND_37 = {1{`RANDOM}};
  salloc_outs_0_flit_flow_egress_node = _RAND_37[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (_T & ~reset) begin
      assert(1'h1); // @[InputUnit.scala 196:13]
    end
    //
    if (_T & _T_3) begin
      assert(_GEN_3 == 3'h0); // @[InputUnit.scala 197:13]
    end
    //
    if (io_router_req_valid & _T_3) begin
      assert(_GEN_139 == 3'h1); // @[InputUnit.scala 224:11]
    end
    //
    if (_T_39 & vcalloc_sel[0] & _T_3) begin
      assert(vcalloc_vals_0); // @[InputUnit.scala 274:17]
    end
    //
    if (_T_39 & vcalloc_sel[1] & _T_3) begin
      assert(vcalloc_vals_1); // @[InputUnit.scala 274:17]
    end
    //
    if (_T_39 & vcalloc_sel[2] & _T_3) begin
      assert(vcalloc_vals_2); // @[InputUnit.scala 274:17]
    end
    //
    if (_T_39 & vcalloc_sel[3] & _T_3) begin
      assert(vcalloc_vals_3); // @[InputUnit.scala 274:17]
    end
  end
endmodule
module InputUnit_1(
  input         clock,
  input         reset,
  output        io_router_req_valid,
  output [1:0]  io_router_req_bits_src_virt_id,
  output [1:0]  io_router_req_bits_flow_ingress_node,
  output [1:0]  io_router_req_bits_flow_egress_node,
  input         io_router_resp_vc_sel_1_0,
  input         io_router_resp_vc_sel_1_1,
  input         io_router_resp_vc_sel_1_2,
  input         io_router_resp_vc_sel_0_0,
  input         io_router_resp_vc_sel_0_1,
  input         io_router_resp_vc_sel_0_2,
  input         io_router_resp_vc_sel_0_3,
  input         io_vcalloc_req_ready,
  output        io_vcalloc_req_valid,
  output        io_vcalloc_req_bits_vc_sel_2_0,
  output        io_vcalloc_req_bits_vc_sel_1_0,
  output        io_vcalloc_req_bits_vc_sel_1_1,
  output        io_vcalloc_req_bits_vc_sel_1_2,
  output        io_vcalloc_req_bits_vc_sel_0_0,
  output        io_vcalloc_req_bits_vc_sel_0_1,
  output        io_vcalloc_req_bits_vc_sel_0_2,
  output        io_vcalloc_req_bits_vc_sel_0_3,
  input         io_vcalloc_resp_vc_sel_2_0,
  input         io_vcalloc_resp_vc_sel_1_0,
  input         io_vcalloc_resp_vc_sel_1_1,
  input         io_vcalloc_resp_vc_sel_1_2,
  input         io_vcalloc_resp_vc_sel_0_0,
  input         io_vcalloc_resp_vc_sel_0_1,
  input         io_vcalloc_resp_vc_sel_0_2,
  input         io_vcalloc_resp_vc_sel_0_3,
  input         io_out_credit_available_2_0,
  input         io_out_credit_available_1_0,
  input         io_out_credit_available_1_1,
  input         io_out_credit_available_1_2,
  input         io_out_credit_available_1_3,
  input         io_out_credit_available_0_0,
  input         io_out_credit_available_0_1,
  input         io_out_credit_available_0_2,
  input         io_out_credit_available_0_3,
  input         io_salloc_req_0_ready,
  output        io_salloc_req_0_valid,
  output        io_salloc_req_0_bits_vc_sel_2_0,
  output        io_salloc_req_0_bits_vc_sel_1_0,
  output        io_salloc_req_0_bits_vc_sel_1_1,
  output        io_salloc_req_0_bits_vc_sel_1_2,
  output        io_salloc_req_0_bits_vc_sel_1_3,
  output        io_salloc_req_0_bits_vc_sel_0_0,
  output        io_salloc_req_0_bits_vc_sel_0_1,
  output        io_salloc_req_0_bits_vc_sel_0_2,
  output        io_salloc_req_0_bits_vc_sel_0_3,
  output        io_salloc_req_0_bits_tail,
  output        io_out_0_valid,
  output        io_out_0_bits_flit_head,
  output        io_out_0_bits_flit_tail,
  output [63:0] io_out_0_bits_flit_payload,
  output [1:0]  io_out_0_bits_flit_flow_ingress_node,
  output [1:0]  io_out_0_bits_flit_flow_egress_node,
  output [1:0]  io_out_0_bits_out_virt_channel,
  output [1:0]  io_debug_va_stall,
  output [1:0]  io_debug_sa_stall,
  input         io_in_flit_0_valid,
  input         io_in_flit_0_bits_head,
  input         io_in_flit_0_bits_tail,
  input  [63:0] io_in_flit_0_bits_payload,
  input  [1:0]  io_in_flit_0_bits_flow_ingress_node,
  input  [1:0]  io_in_flit_0_bits_flow_egress_node,
  input  [1:0]  io_in_flit_0_bits_virt_channel_id,
  output [3:0]  io_in_credit_return,
  output [3:0]  io_in_vc_free
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
`endif // RANDOMIZE_REG_INIT
  wire  input_buffer_clock; // @[InputUnit.scala 180:28]
  wire  input_buffer_reset; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_enq_0_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_enq_0_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_enq_0_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_enq_0_bits_payload; // @[InputUnit.scala 180:28]
  wire [1:0] input_buffer_io_enq_0_bits_virt_channel_id; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_0_ready; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_0_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_0_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_0_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_deq_0_bits_payload; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_ready; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_deq_1_bits_payload; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_ready; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_deq_2_bits_payload; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_3_ready; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_3_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_3_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_3_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_deq_3_bits_payload; // @[InputUnit.scala 180:28]
  wire  route_arbiter_io_in_0_valid; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_0_bits_flow_ingress_node; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_0_bits_flow_egress_node; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_1_ready; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_1_valid; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_1_bits_flow_ingress_node; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_1_bits_flow_egress_node; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_2_ready; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_2_valid; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_2_bits_flow_ingress_node; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_2_bits_flow_egress_node; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_3_ready; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_3_valid; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_3_bits_flow_ingress_node; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_3_bits_flow_egress_node; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_out_valid; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_out_bits_src_virt_id; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_out_bits_flow_ingress_node; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_out_bits_flow_egress_node; // @[InputUnit.scala 186:29]
  wire  salloc_arb_clock; // @[InputUnit.scala 279:26]
  wire  salloc_arb_reset; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_bits_vc_sel_2_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_bits_vc_sel_1_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_bits_tail; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_vc_sel_2_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_vc_sel_1_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_vc_sel_1_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_vc_sel_0_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_tail; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_2_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_1_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_1_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_1_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_0_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_0_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_tail; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_2_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_1_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_1_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_1_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_1_3; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_0_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_0_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_0_3; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_tail; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_2_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_1_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_1_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_1_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_1_3; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_0_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_0_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_0_3; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_tail; // @[InputUnit.scala 279:26]
  wire [3:0] salloc_arb_io_chosen_oh_0; // @[InputUnit.scala 279:26]
  reg [2:0] states_0_g; // @[InputUnit.scala 191:19]
  reg  states_0_vc_sel_2_0; // @[InputUnit.scala 191:19]
  reg  states_0_vc_sel_1_0; // @[InputUnit.scala 191:19]
  reg  states_0_vc_sel_0_0; // @[InputUnit.scala 191:19]
  reg [1:0] states_0_flow_ingress_node; // @[InputUnit.scala 191:19]
  reg [1:0] states_0_flow_egress_node; // @[InputUnit.scala 191:19]
  reg [2:0] states_1_g; // @[InputUnit.scala 191:19]
  reg  states_1_vc_sel_2_0; // @[InputUnit.scala 191:19]
  reg  states_1_vc_sel_1_0; // @[InputUnit.scala 191:19]
  reg  states_1_vc_sel_0_0; // @[InputUnit.scala 191:19]
  reg  states_1_vc_sel_0_1; // @[InputUnit.scala 191:19]
  reg [1:0] states_1_flow_ingress_node; // @[InputUnit.scala 191:19]
  reg [1:0] states_1_flow_egress_node; // @[InputUnit.scala 191:19]
  reg [2:0] states_2_g; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_2_0; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_1_0; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_1_1; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_0_0; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_0_1; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_0_2; // @[InputUnit.scala 191:19]
  reg [1:0] states_2_flow_ingress_node; // @[InputUnit.scala 191:19]
  reg [1:0] states_2_flow_egress_node; // @[InputUnit.scala 191:19]
  reg [2:0] states_3_g; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_2_0; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_1_0; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_1_1; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_1_2; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_0_0; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_0_1; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_0_2; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_0_3; // @[InputUnit.scala 191:19]
  reg [1:0] states_3_flow_ingress_node; // @[InputUnit.scala 191:19]
  reg [1:0] states_3_flow_egress_node; // @[InputUnit.scala 191:19]
  wire  _T = io_in_flit_0_valid & io_in_flit_0_bits_head; // @[InputUnit.scala 194:32]
  wire  _T_3 = ~reset; // @[InputUnit.scala 196:13]
  wire [2:0] _GEN_1 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? states_1_g : states_0_g; // @[InputUnit.scala 197:{27,27}]
  wire [2:0] _GEN_2 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? states_2_g : _GEN_1; // @[InputUnit.scala 197:{27,27}]
  wire [2:0] _GEN_3 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? states_3_g : _GEN_2; // @[InputUnit.scala 197:{27,27}]
  wire  at_dest = io_in_flit_0_bits_flow_egress_node == 2'h0; // @[InputUnit.scala 198:57]
  wire [2:0] _states_g_T = at_dest ? 3'h2 : 3'h1; // @[InputUnit.scala 199:26]
  wire [2:0] _GEN_4 = 2'h0 == io_in_flit_0_bits_virt_channel_id ? _states_g_T : states_0_g; // @[InputUnit.scala 191:19 199:{20,20}]
  wire [2:0] _GEN_5 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? _states_g_T : states_1_g; // @[InputUnit.scala 191:19 199:{20,20}]
  wire [2:0] _GEN_6 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? _states_g_T : states_2_g; // @[InputUnit.scala 191:19 199:{20,20}]
  wire [2:0] _GEN_7 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? _states_g_T : states_3_g; // @[InputUnit.scala 191:19 199:{20,20}]
  wire  _GEN_8 = 2'h0 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_0_vc_sel_0_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_9 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_1_vc_sel_0_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_10 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_0_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_11 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_0_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_13 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_1_vc_sel_0_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_14 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_0_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_15 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_0_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_18 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_0_2; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_19 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_0_2; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_23 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_0_3; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_24 = 2'h0 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_0_vc_sel_1_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_25 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_1_vc_sel_1_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_26 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_1_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_27 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_1_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_30 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_1_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_31 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_1_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_35 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_1_2; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_40 = 2'h0 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_0_vc_sel_2_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_41 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_1_vc_sel_2_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_42 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_2_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_43 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_2_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_44 = 2'h0 == io_in_flit_0_bits_virt_channel_id | _GEN_40; // @[InputUnit.scala 203:{44,44}]
  wire  _GEN_45 = 2'h1 == io_in_flit_0_bits_virt_channel_id | _GEN_41; // @[InputUnit.scala 203:{44,44}]
  wire  _GEN_46 = 2'h2 == io_in_flit_0_bits_virt_channel_id | _GEN_42; // @[InputUnit.scala 203:{44,44}]
  wire  _GEN_47 = 2'h3 == io_in_flit_0_bits_virt_channel_id | _GEN_43; // @[InputUnit.scala 203:{44,44}]
  wire [2:0] _GEN_72 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_4 : states_0_g; // @[InputUnit.scala 191:19 194:60]
  wire [2:0] _GEN_73 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_5 : states_1_g; // @[InputUnit.scala 191:19 194:60]
  wire [2:0] _GEN_74 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_6 : states_2_g; // @[InputUnit.scala 191:19 194:60]
  wire [2:0] _GEN_75 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_7 : states_3_g; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_76 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_8 : states_0_vc_sel_0_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_77 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_9 : states_1_vc_sel_0_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_78 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_10 : states_2_vc_sel_0_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_79 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_11 : states_3_vc_sel_0_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_81 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_13 : states_1_vc_sel_0_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_82 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_14 : states_2_vc_sel_0_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_83 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_15 : states_3_vc_sel_0_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_86 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_18 : states_2_vc_sel_0_2; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_87 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_19 : states_3_vc_sel_0_2; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_91 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_23 : states_3_vc_sel_0_3; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_92 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_24 : states_0_vc_sel_1_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_93 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_25 : states_1_vc_sel_1_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_94 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_26 : states_2_vc_sel_1_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_95 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_27 : states_3_vc_sel_1_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_98 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_30 : states_2_vc_sel_1_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_99 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_31 : states_3_vc_sel_1_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_103 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_35 : states_3_vc_sel_1_2; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_108 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_44 : states_0_vc_sel_2_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_109 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_45 : states_1_vc_sel_2_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_110 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_46 : states_2_vc_sel_2_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_111 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_47 : states_3_vc_sel_2_0; // @[InputUnit.scala 191:19 194:60]
  wire  _T_10 = route_arbiter_io_in_0_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_132 = _T_10 ? 3'h2 : _GEN_72; // @[InputUnit.scala 215:{23,29}]
  wire  _T_11 = route_arbiter_io_in_1_ready & route_arbiter_io_in_1_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_133 = _T_11 ? 3'h2 : _GEN_73; // @[InputUnit.scala 215:{23,29}]
  wire  _T_12 = route_arbiter_io_in_2_ready & route_arbiter_io_in_2_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_134 = _T_12 ? 3'h2 : _GEN_74; // @[InputUnit.scala 215:{23,29}]
  wire  _T_13 = route_arbiter_io_in_3_ready & route_arbiter_io_in_3_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_135 = _T_13 ? 3'h2 : _GEN_75; // @[InputUnit.scala 215:{23,29}]
  wire [2:0] _GEN_137 = 2'h1 == io_router_req_bits_src_virt_id ? states_1_g : states_0_g; // @[InputUnit.scala 224:{25,25}]
  wire [2:0] _GEN_138 = 2'h2 == io_router_req_bits_src_virt_id ? states_2_g : _GEN_137; // @[InputUnit.scala 224:{25,25}]
  wire [2:0] _GEN_139 = 2'h3 == io_router_req_bits_src_virt_id ? states_3_g : _GEN_138; // @[InputUnit.scala 224:{25,25}]
  wire [2:0] _GEN_140 = 2'h0 == io_router_req_bits_src_virt_id ? 3'h2 : _GEN_132; // @[InputUnit.scala 225:{18,18}]
  wire [2:0] _GEN_141 = 2'h1 == io_router_req_bits_src_virt_id ? 3'h2 : _GEN_133; // @[InputUnit.scala 225:{18,18}]
  wire [2:0] _GEN_142 = 2'h2 == io_router_req_bits_src_virt_id ? 3'h2 : _GEN_134; // @[InputUnit.scala 225:{18,18}]
  wire [2:0] _GEN_143 = 2'h3 == io_router_req_bits_src_virt_id ? 3'h2 : _GEN_135; // @[InputUnit.scala 225:{18,18}]
  wire  _GEN_144 = 2'h0 == io_router_req_bits_src_virt_id ? 1'h0 : _GEN_108; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_145 = 2'h0 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_0 : _GEN_92; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_149 = 2'h0 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_0 : _GEN_76; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_153 = 2'h1 == io_router_req_bits_src_virt_id ? 1'h0 : _GEN_109; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_154 = 2'h1 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_0 : _GEN_93; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_158 = 2'h1 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_0 : _GEN_77; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_159 = 2'h1 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_1 : _GEN_81; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_162 = 2'h2 == io_router_req_bits_src_virt_id ? 1'h0 : _GEN_110; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_163 = 2'h2 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_0 : _GEN_94; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_164 = 2'h2 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_1 : _GEN_98; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_167 = 2'h2 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_0 : _GEN_78; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_168 = 2'h2 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_1 : _GEN_82; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_169 = 2'h2 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_2 : _GEN_86; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_171 = 2'h3 == io_router_req_bits_src_virt_id ? 1'h0 : _GEN_111; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_172 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_0 : _GEN_95; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_173 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_1 : _GEN_99; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_174 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_2 : _GEN_103; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_176 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_0 : _GEN_79; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_177 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_1 : _GEN_83; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_178 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_2 : _GEN_87; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_179 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_3 : _GEN_91; // @[InputUnit.scala 227:25 228:26]
  wire [2:0] _GEN_180 = io_router_req_valid ? _GEN_140 : _GEN_132; // @[InputUnit.scala 222:31]
  wire [2:0] _GEN_181 = io_router_req_valid ? _GEN_141 : _GEN_133; // @[InputUnit.scala 222:31]
  wire [2:0] _GEN_182 = io_router_req_valid ? _GEN_142 : _GEN_134; // @[InputUnit.scala 222:31]
  wire [2:0] _GEN_183 = io_router_req_valid ? _GEN_143 : _GEN_135; // @[InputUnit.scala 222:31]
  wire  _GEN_184 = io_router_req_valid ? _GEN_144 : _GEN_108; // @[InputUnit.scala 222:31]
  wire  _GEN_185 = io_router_req_valid ? _GEN_145 : _GEN_92; // @[InputUnit.scala 222:31]
  wire  _GEN_189 = io_router_req_valid ? _GEN_149 : _GEN_76; // @[InputUnit.scala 222:31]
  wire  _GEN_193 = io_router_req_valid ? _GEN_153 : _GEN_109; // @[InputUnit.scala 222:31]
  wire  _GEN_194 = io_router_req_valid ? _GEN_154 : _GEN_93; // @[InputUnit.scala 222:31]
  wire  _GEN_198 = io_router_req_valid ? _GEN_158 : _GEN_77; // @[InputUnit.scala 222:31]
  wire  _GEN_199 = io_router_req_valid ? _GEN_159 : _GEN_81; // @[InputUnit.scala 222:31]
  wire  _GEN_202 = io_router_req_valid ? _GEN_162 : _GEN_110; // @[InputUnit.scala 222:31]
  wire  _GEN_203 = io_router_req_valid ? _GEN_163 : _GEN_94; // @[InputUnit.scala 222:31]
  wire  _GEN_204 = io_router_req_valid ? _GEN_164 : _GEN_98; // @[InputUnit.scala 222:31]
  wire  _GEN_207 = io_router_req_valid ? _GEN_167 : _GEN_78; // @[InputUnit.scala 222:31]
  wire  _GEN_208 = io_router_req_valid ? _GEN_168 : _GEN_82; // @[InputUnit.scala 222:31]
  wire  _GEN_209 = io_router_req_valid ? _GEN_169 : _GEN_86; // @[InputUnit.scala 222:31]
  wire  _GEN_211 = io_router_req_valid ? _GEN_171 : _GEN_111; // @[InputUnit.scala 222:31]
  wire  _GEN_212 = io_router_req_valid ? _GEN_172 : _GEN_95; // @[InputUnit.scala 222:31]
  wire  _GEN_213 = io_router_req_valid ? _GEN_173 : _GEN_99; // @[InputUnit.scala 222:31]
  wire  _GEN_214 = io_router_req_valid ? _GEN_174 : _GEN_103; // @[InputUnit.scala 222:31]
  wire  _GEN_216 = io_router_req_valid ? _GEN_176 : _GEN_79; // @[InputUnit.scala 222:31]
  wire  _GEN_217 = io_router_req_valid ? _GEN_177 : _GEN_83; // @[InputUnit.scala 222:31]
  wire  _GEN_218 = io_router_req_valid ? _GEN_178 : _GEN_87; // @[InputUnit.scala 222:31]
  wire  _GEN_219 = io_router_req_valid ? _GEN_179 : _GEN_91; // @[InputUnit.scala 222:31]
  reg [3:0] mask; // @[InputUnit.scala 233:21]
  wire  vcalloc_vals_1 = states_1_g == 3'h2; // @[InputUnit.scala 249:32]
  wire  vcalloc_vals_0 = states_0_g == 3'h2; // @[InputUnit.scala 249:32]
  wire  vcalloc_vals_3 = states_3_g == 3'h2; // @[InputUnit.scala 249:32]
  wire  vcalloc_vals_2 = states_2_g == 3'h2; // @[InputUnit.scala 249:32]
  wire [3:0] _vcalloc_filter_T = {vcalloc_vals_3,vcalloc_vals_2,vcalloc_vals_1,vcalloc_vals_0}; // @[InputUnit.scala 236:59]
  wire [3:0] _vcalloc_filter_T_2 = ~mask; // @[InputUnit.scala 236:89]
  wire [3:0] _vcalloc_filter_T_3 = _vcalloc_filter_T & _vcalloc_filter_T_2; // @[InputUnit.scala 236:87]
  wire [7:0] _vcalloc_filter_T_4 = {vcalloc_vals_3,vcalloc_vals_2,vcalloc_vals_1,vcalloc_vals_0,_vcalloc_filter_T_3}; // @[Cat.scala 33:92]
  wire [7:0] _vcalloc_filter_T_13 = _vcalloc_filter_T_4[7] ? 8'h80 : 8'h0; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_14 = _vcalloc_filter_T_4[6] ? 8'h40 : _vcalloc_filter_T_13; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_15 = _vcalloc_filter_T_4[5] ? 8'h20 : _vcalloc_filter_T_14; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_16 = _vcalloc_filter_T_4[4] ? 8'h10 : _vcalloc_filter_T_15; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_17 = _vcalloc_filter_T_4[3] ? 8'h8 : _vcalloc_filter_T_16; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_18 = _vcalloc_filter_T_4[2] ? 8'h4 : _vcalloc_filter_T_17; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_19 = _vcalloc_filter_T_4[1] ? 8'h2 : _vcalloc_filter_T_18; // @[Mux.scala 47:70]
  wire [7:0] vcalloc_filter = _vcalloc_filter_T_4[0] ? 8'h1 : _vcalloc_filter_T_19; // @[Mux.scala 47:70]
  wire [3:0] vcalloc_sel = vcalloc_filter[3:0] | vcalloc_filter[7:4]; // @[InputUnit.scala 237:58]
  wire [3:0] _mask_T = 4'h1 << io_router_req_bits_src_virt_id; // @[InputUnit.scala 240:18]
  wire [3:0] _mask_T_2 = _mask_T - 4'h1; // @[InputUnit.scala 240:53]
  wire  _T_26 = vcalloc_vals_0 | vcalloc_vals_1 | vcalloc_vals_2 | vcalloc_vals_3; // @[package.scala 73:59]
  wire [1:0] _mask_T_12 = vcalloc_sel[1] ? 2'h3 : 2'h0; // @[Mux.scala 27:73]
  wire [2:0] _mask_T_13 = vcalloc_sel[2] ? 3'h7 : 3'h0; // @[Mux.scala 27:73]
  wire [3:0] _mask_T_14 = vcalloc_sel[3] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [1:0] _GEN_60 = {{1'd0}, vcalloc_sel[0]}; // @[Mux.scala 27:73]
  wire [1:0] _mask_T_15 = _GEN_60 | _mask_T_12; // @[Mux.scala 27:73]
  wire [2:0] _GEN_61 = {{1'd0}, _mask_T_15}; // @[Mux.scala 27:73]
  wire [2:0] _mask_T_16 = _GEN_61 | _mask_T_13; // @[Mux.scala 27:73]
  wire [3:0] _GEN_62 = {{1'd0}, _mask_T_16}; // @[Mux.scala 27:73]
  wire [3:0] _mask_T_17 = _GEN_62 | _mask_T_14; // @[Mux.scala 27:73]
  wire [2:0] _GEN_222 = vcalloc_vals_0 & vcalloc_sel[0] & io_vcalloc_req_ready ? 3'h3 : _GEN_180; // @[InputUnit.scala 253:{76,82}]
  wire [2:0] _GEN_223 = vcalloc_vals_1 & vcalloc_sel[1] & io_vcalloc_req_ready ? 3'h3 : _GEN_181; // @[InputUnit.scala 253:{76,82}]
  wire [2:0] _GEN_224 = vcalloc_vals_2 & vcalloc_sel[2] & io_vcalloc_req_ready ? 3'h3 : _GEN_182; // @[InputUnit.scala 253:{76,82}]
  wire [2:0] _GEN_225 = vcalloc_vals_3 & vcalloc_sel[3] & io_vcalloc_req_ready ? 3'h3 : _GEN_183; // @[InputUnit.scala 253:{76,82}]
  wire [1:0] _io_debug_va_stall_T = vcalloc_vals_0 + vcalloc_vals_1; // @[Bitwise.scala 51:90]
  wire [1:0] _io_debug_va_stall_T_2 = vcalloc_vals_2 + vcalloc_vals_3; // @[Bitwise.scala 51:90]
  wire [2:0] _io_debug_va_stall_T_4 = _io_debug_va_stall_T + _io_debug_va_stall_T_2; // @[Bitwise.scala 51:90]
  wire [2:0] _GEN_63 = {{2'd0}, io_vcalloc_req_ready}; // @[InputUnit.scala 266:47]
  wire [2:0] _io_debug_va_stall_T_7 = _io_debug_va_stall_T_4 - _GEN_63; // @[InputUnit.scala 266:47]
  wire  _T_39 = io_vcalloc_req_ready & io_vcalloc_req_valid; // @[Decoupled.scala 51:35]
  wire [8:0] _credit_available_T = {states_0_vc_sel_2_0,1'h0,1'h0,1'h0,states_0_vc_sel_1_0,2'h0,1'h0,states_0_vc_sel_0_0
    }; // @[InputUnit.scala 287:40]
  wire [8:0] _credit_available_T_1 = {io_out_credit_available_2_0,io_out_credit_available_1_3,
    io_out_credit_available_1_2,io_out_credit_available_1_1,io_out_credit_available_1_0,io_out_credit_available_0_3,
    io_out_credit_available_0_2,io_out_credit_available_0_1,io_out_credit_available_0_0}; // @[InputUnit.scala 287:73]
  wire [8:0] _credit_available_T_2 = _credit_available_T & _credit_available_T_1; // @[InputUnit.scala 287:47]
  wire  credit_available = _credit_available_T_2 != 9'h0; // @[InputUnit.scala 287:81]
  wire  _T_60 = salloc_arb_io_in_0_ready & salloc_arb_io_in_0_valid; // @[Decoupled.scala 51:35]
  wire [8:0] _credit_available_T_3 = {states_1_vc_sel_2_0,1'h0,1'h0,1'h0,states_1_vc_sel_1_0,2'h0,states_1_vc_sel_0_1,
    states_1_vc_sel_0_0}; // @[InputUnit.scala 287:40]
  wire [8:0] _credit_available_T_5 = _credit_available_T_3 & _credit_available_T_1; // @[InputUnit.scala 287:47]
  wire  credit_available_1 = _credit_available_T_5 != 9'h0; // @[InputUnit.scala 287:81]
  wire  _T_62 = salloc_arb_io_in_1_ready & salloc_arb_io_in_1_valid; // @[Decoupled.scala 51:35]
  wire [8:0] _credit_available_T_6 = {states_2_vc_sel_2_0,1'h0,1'h0,states_2_vc_sel_1_1,states_2_vc_sel_1_0,1'h0,
    states_2_vc_sel_0_2,states_2_vc_sel_0_1,states_2_vc_sel_0_0}; // @[InputUnit.scala 287:40]
  wire [8:0] _credit_available_T_8 = _credit_available_T_6 & _credit_available_T_1; // @[InputUnit.scala 287:47]
  wire  credit_available_2 = _credit_available_T_8 != 9'h0; // @[InputUnit.scala 287:81]
  wire  _T_64 = salloc_arb_io_in_2_ready & salloc_arb_io_in_2_valid; // @[Decoupled.scala 51:35]
  wire [8:0] _credit_available_T_9 = {states_3_vc_sel_2_0,1'h0,states_3_vc_sel_1_2,states_3_vc_sel_1_1,
    states_3_vc_sel_1_0,states_3_vc_sel_0_3,states_3_vc_sel_0_2,states_3_vc_sel_0_1,states_3_vc_sel_0_0}; // @[InputUnit.scala 287:40]
  wire [8:0] _credit_available_T_11 = _credit_available_T_9 & _credit_available_T_1; // @[InputUnit.scala 287:47]
  wire  credit_available_3 = _credit_available_T_11 != 9'h0; // @[InputUnit.scala 287:81]
  wire  _T_66 = salloc_arb_io_in_3_ready & salloc_arb_io_in_3_valid; // @[Decoupled.scala 51:35]
  wire  _io_debug_sa_stall_T_1 = salloc_arb_io_in_0_valid & ~salloc_arb_io_in_0_ready; // @[InputUnit.scala 301:67]
  wire  _io_debug_sa_stall_T_3 = salloc_arb_io_in_1_valid & ~salloc_arb_io_in_1_ready; // @[InputUnit.scala 301:67]
  wire  _io_debug_sa_stall_T_5 = salloc_arb_io_in_2_valid & ~salloc_arb_io_in_2_ready; // @[InputUnit.scala 301:67]
  wire  _io_debug_sa_stall_T_7 = salloc_arb_io_in_3_valid & ~salloc_arb_io_in_3_ready; // @[InputUnit.scala 301:67]
  wire [1:0] _io_debug_sa_stall_T_8 = _io_debug_sa_stall_T_1 + _io_debug_sa_stall_T_3; // @[Bitwise.scala 51:90]
  wire [1:0] _io_debug_sa_stall_T_10 = _io_debug_sa_stall_T_5 + _io_debug_sa_stall_T_7; // @[Bitwise.scala 51:90]
  wire [2:0] _io_debug_sa_stall_T_12 = _io_debug_sa_stall_T_8 + _io_debug_sa_stall_T_10; // @[Bitwise.scala 51:90]
  reg  salloc_outs_0_valid; // @[InputUnit.scala 318:8]
  reg [1:0] salloc_outs_0_out_vid; // @[InputUnit.scala 318:8]
  reg  salloc_outs_0_flit_head; // @[InputUnit.scala 318:8]
  reg  salloc_outs_0_flit_tail; // @[InputUnit.scala 318:8]
  reg [63:0] salloc_outs_0_flit_payload; // @[InputUnit.scala 318:8]
  reg [1:0] salloc_outs_0_flit_flow_ingress_node; // @[InputUnit.scala 318:8]
  reg [1:0] salloc_outs_0_flit_flow_egress_node; // @[InputUnit.scala 318:8]
  wire  _io_in_credit_return_T = salloc_arb_io_out_0_ready & salloc_arb_io_out_0_valid; // @[Decoupled.scala 51:35]
  wire  _io_in_vc_free_T_11 = salloc_arb_io_chosen_oh_0[0] & input_buffer_io_deq_0_bits_tail | salloc_arb_io_chosen_oh_0
    [1] & input_buffer_io_deq_1_bits_tail | salloc_arb_io_chosen_oh_0[2] & input_buffer_io_deq_2_bits_tail |
    salloc_arb_io_chosen_oh_0[3] & input_buffer_io_deq_3_bits_tail; // @[Mux.scala 27:73]
  wire  vc_sel_0_0 = salloc_arb_io_chosen_oh_0[0] & states_0_vc_sel_0_0 | salloc_arb_io_chosen_oh_0[1] &
    states_1_vc_sel_0_0 | salloc_arb_io_chosen_oh_0[2] & states_2_vc_sel_0_0 | salloc_arb_io_chosen_oh_0[3] &
    states_3_vc_sel_0_0; // @[Mux.scala 27:73]
  wire  vc_sel_0_1 = salloc_arb_io_chosen_oh_0[1] & states_1_vc_sel_0_1 | salloc_arb_io_chosen_oh_0[2] &
    states_2_vc_sel_0_1 | salloc_arb_io_chosen_oh_0[3] & states_3_vc_sel_0_1; // @[Mux.scala 27:73]
  wire  vc_sel_0_2 = salloc_arb_io_chosen_oh_0[2] & states_2_vc_sel_0_2 | salloc_arb_io_chosen_oh_0[3] &
    states_3_vc_sel_0_2; // @[Mux.scala 27:73]
  wire  vc_sel_0_3 = salloc_arb_io_chosen_oh_0[3] & states_3_vc_sel_0_3; // @[Mux.scala 27:73]
  wire  vc_sel_1_0 = salloc_arb_io_chosen_oh_0[0] & states_0_vc_sel_1_0 | salloc_arb_io_chosen_oh_0[1] &
    states_1_vc_sel_1_0 | salloc_arb_io_chosen_oh_0[2] & states_2_vc_sel_1_0 | salloc_arb_io_chosen_oh_0[3] &
    states_3_vc_sel_1_0; // @[Mux.scala 27:73]
  wire  vc_sel_1_1 = salloc_arb_io_chosen_oh_0[2] & states_2_vc_sel_1_1 | salloc_arb_io_chosen_oh_0[3] &
    states_3_vc_sel_1_1; // @[Mux.scala 27:73]
  wire  vc_sel_1_2 = salloc_arb_io_chosen_oh_0[3] & states_3_vc_sel_1_2; // @[Mux.scala 27:73]
  wire  channel_oh_0 = vc_sel_0_0 | vc_sel_0_1 | vc_sel_0_2 | vc_sel_0_3; // @[InputUnit.scala 334:43]
  wire  channel_oh_1 = vc_sel_1_0 | vc_sel_1_1 | vc_sel_1_2; // @[InputUnit.scala 334:43]
  wire [3:0] _virt_channel_T = {vc_sel_0_3,vc_sel_0_2,vc_sel_0_1,vc_sel_0_0}; // @[OneHot.scala 22:45]
  wire [1:0] virt_channel_hi_1 = _virt_channel_T[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] virt_channel_lo_1 = _virt_channel_T[1:0]; // @[OneHot.scala 31:18]
  wire  _virt_channel_T_1 = |virt_channel_hi_1; // @[OneHot.scala 32:14]
  wire [1:0] _virt_channel_T_2 = virt_channel_hi_1 | virt_channel_lo_1; // @[OneHot.scala 32:28]
  wire [1:0] _virt_channel_T_4 = {_virt_channel_T_1,_virt_channel_T_2[1]}; // @[Cat.scala 33:92]
  wire [3:0] _virt_channel_T_5 = {1'h0,vc_sel_1_2,vc_sel_1_1,vc_sel_1_0}; // @[OneHot.scala 22:45]
  wire [1:0] virt_channel_hi_3 = _virt_channel_T_5[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] virt_channel_lo_3 = _virt_channel_T_5[1:0]; // @[OneHot.scala 31:18]
  wire  _virt_channel_T_6 = |virt_channel_hi_3; // @[OneHot.scala 32:14]
  wire [1:0] _virt_channel_T_7 = virt_channel_hi_3 | virt_channel_lo_3; // @[OneHot.scala 32:28]
  wire [1:0] _virt_channel_T_9 = {_virt_channel_T_6,_virt_channel_T_7[1]}; // @[Cat.scala 33:92]
  wire [1:0] _virt_channel_T_10 = channel_oh_0 ? _virt_channel_T_4 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _virt_channel_T_11 = channel_oh_1 ? _virt_channel_T_9 : 2'h0; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_4 = salloc_arb_io_chosen_oh_0[0] ? input_buffer_io_deq_0_bits_payload : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_5 = salloc_arb_io_chosen_oh_0[1] ? input_buffer_io_deq_1_bits_payload : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_6 = salloc_arb_io_chosen_oh_0[2] ? input_buffer_io_deq_2_bits_payload : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_7 = salloc_arb_io_chosen_oh_0[3] ? input_buffer_io_deq_3_bits_payload : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_8 = _salloc_outs_0_flit_payload_T_4 | _salloc_outs_0_flit_payload_T_5; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_9 = _salloc_outs_0_flit_payload_T_8 | _salloc_outs_0_flit_payload_T_6; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_11 = salloc_arb_io_chosen_oh_0[0] ? states_0_flow_egress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_12 = salloc_arb_io_chosen_oh_0[1] ? states_1_flow_egress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_13 = salloc_arb_io_chosen_oh_0[2] ? states_2_flow_egress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_14 = salloc_arb_io_chosen_oh_0[3] ? states_3_flow_egress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_15 = _salloc_outs_0_flit_flow_T_11 | _salloc_outs_0_flit_flow_T_12; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_16 = _salloc_outs_0_flit_flow_T_15 | _salloc_outs_0_flit_flow_T_13; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_25 = salloc_arb_io_chosen_oh_0[0] ? states_0_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_26 = salloc_arb_io_chosen_oh_0[1] ? states_1_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_27 = salloc_arb_io_chosen_oh_0[2] ? states_2_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_28 = salloc_arb_io_chosen_oh_0[3] ? states_3_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_29 = _salloc_outs_0_flit_flow_T_25 | _salloc_outs_0_flit_flow_T_26; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_30 = _salloc_outs_0_flit_flow_T_29 | _salloc_outs_0_flit_flow_T_27; // @[Mux.scala 27:73]
  InputBuffer input_buffer ( // @[InputUnit.scala 180:28]
    .clock(input_buffer_clock),
    .reset(input_buffer_reset),
    .io_enq_0_valid(input_buffer_io_enq_0_valid),
    .io_enq_0_bits_head(input_buffer_io_enq_0_bits_head),
    .io_enq_0_bits_tail(input_buffer_io_enq_0_bits_tail),
    .io_enq_0_bits_payload(input_buffer_io_enq_0_bits_payload),
    .io_enq_0_bits_virt_channel_id(input_buffer_io_enq_0_bits_virt_channel_id),
    .io_deq_0_ready(input_buffer_io_deq_0_ready),
    .io_deq_0_valid(input_buffer_io_deq_0_valid),
    .io_deq_0_bits_head(input_buffer_io_deq_0_bits_head),
    .io_deq_0_bits_tail(input_buffer_io_deq_0_bits_tail),
    .io_deq_0_bits_payload(input_buffer_io_deq_0_bits_payload),
    .io_deq_1_ready(input_buffer_io_deq_1_ready),
    .io_deq_1_valid(input_buffer_io_deq_1_valid),
    .io_deq_1_bits_head(input_buffer_io_deq_1_bits_head),
    .io_deq_1_bits_tail(input_buffer_io_deq_1_bits_tail),
    .io_deq_1_bits_payload(input_buffer_io_deq_1_bits_payload),
    .io_deq_2_ready(input_buffer_io_deq_2_ready),
    .io_deq_2_valid(input_buffer_io_deq_2_valid),
    .io_deq_2_bits_head(input_buffer_io_deq_2_bits_head),
    .io_deq_2_bits_tail(input_buffer_io_deq_2_bits_tail),
    .io_deq_2_bits_payload(input_buffer_io_deq_2_bits_payload),
    .io_deq_3_ready(input_buffer_io_deq_3_ready),
    .io_deq_3_valid(input_buffer_io_deq_3_valid),
    .io_deq_3_bits_head(input_buffer_io_deq_3_bits_head),
    .io_deq_3_bits_tail(input_buffer_io_deq_3_bits_tail),
    .io_deq_3_bits_payload(input_buffer_io_deq_3_bits_payload)
  );
  Arbiter route_arbiter ( // @[InputUnit.scala 186:29]
    .io_in_0_valid(route_arbiter_io_in_0_valid),
    .io_in_0_bits_flow_ingress_node(route_arbiter_io_in_0_bits_flow_ingress_node),
    .io_in_0_bits_flow_egress_node(route_arbiter_io_in_0_bits_flow_egress_node),
    .io_in_1_ready(route_arbiter_io_in_1_ready),
    .io_in_1_valid(route_arbiter_io_in_1_valid),
    .io_in_1_bits_flow_ingress_node(route_arbiter_io_in_1_bits_flow_ingress_node),
    .io_in_1_bits_flow_egress_node(route_arbiter_io_in_1_bits_flow_egress_node),
    .io_in_2_ready(route_arbiter_io_in_2_ready),
    .io_in_2_valid(route_arbiter_io_in_2_valid),
    .io_in_2_bits_flow_ingress_node(route_arbiter_io_in_2_bits_flow_ingress_node),
    .io_in_2_bits_flow_egress_node(route_arbiter_io_in_2_bits_flow_egress_node),
    .io_in_3_ready(route_arbiter_io_in_3_ready),
    .io_in_3_valid(route_arbiter_io_in_3_valid),
    .io_in_3_bits_flow_ingress_node(route_arbiter_io_in_3_bits_flow_ingress_node),
    .io_in_3_bits_flow_egress_node(route_arbiter_io_in_3_bits_flow_egress_node),
    .io_out_valid(route_arbiter_io_out_valid),
    .io_out_bits_src_virt_id(route_arbiter_io_out_bits_src_virt_id),
    .io_out_bits_flow_ingress_node(route_arbiter_io_out_bits_flow_ingress_node),
    .io_out_bits_flow_egress_node(route_arbiter_io_out_bits_flow_egress_node)
  );
  SwitchArbiter salloc_arb ( // @[InputUnit.scala 279:26]
    .clock(salloc_arb_clock),
    .reset(salloc_arb_reset),
    .io_in_0_ready(salloc_arb_io_in_0_ready),
    .io_in_0_valid(salloc_arb_io_in_0_valid),
    .io_in_0_bits_vc_sel_2_0(salloc_arb_io_in_0_bits_vc_sel_2_0),
    .io_in_0_bits_vc_sel_1_0(salloc_arb_io_in_0_bits_vc_sel_1_0),
    .io_in_0_bits_vc_sel_0_0(salloc_arb_io_in_0_bits_vc_sel_0_0),
    .io_in_0_bits_tail(salloc_arb_io_in_0_bits_tail),
    .io_in_1_ready(salloc_arb_io_in_1_ready),
    .io_in_1_valid(salloc_arb_io_in_1_valid),
    .io_in_1_bits_vc_sel_2_0(salloc_arb_io_in_1_bits_vc_sel_2_0),
    .io_in_1_bits_vc_sel_1_0(salloc_arb_io_in_1_bits_vc_sel_1_0),
    .io_in_1_bits_vc_sel_1_1(salloc_arb_io_in_1_bits_vc_sel_1_1),
    .io_in_1_bits_vc_sel_0_0(salloc_arb_io_in_1_bits_vc_sel_0_0),
    .io_in_1_bits_vc_sel_0_1(salloc_arb_io_in_1_bits_vc_sel_0_1),
    .io_in_1_bits_tail(salloc_arb_io_in_1_bits_tail),
    .io_in_2_ready(salloc_arb_io_in_2_ready),
    .io_in_2_valid(salloc_arb_io_in_2_valid),
    .io_in_2_bits_vc_sel_2_0(salloc_arb_io_in_2_bits_vc_sel_2_0),
    .io_in_2_bits_vc_sel_1_0(salloc_arb_io_in_2_bits_vc_sel_1_0),
    .io_in_2_bits_vc_sel_1_1(salloc_arb_io_in_2_bits_vc_sel_1_1),
    .io_in_2_bits_vc_sel_1_2(salloc_arb_io_in_2_bits_vc_sel_1_2),
    .io_in_2_bits_vc_sel_0_0(salloc_arb_io_in_2_bits_vc_sel_0_0),
    .io_in_2_bits_vc_sel_0_1(salloc_arb_io_in_2_bits_vc_sel_0_1),
    .io_in_2_bits_vc_sel_0_2(salloc_arb_io_in_2_bits_vc_sel_0_2),
    .io_in_2_bits_tail(salloc_arb_io_in_2_bits_tail),
    .io_in_3_ready(salloc_arb_io_in_3_ready),
    .io_in_3_valid(salloc_arb_io_in_3_valid),
    .io_in_3_bits_vc_sel_2_0(salloc_arb_io_in_3_bits_vc_sel_2_0),
    .io_in_3_bits_vc_sel_1_0(salloc_arb_io_in_3_bits_vc_sel_1_0),
    .io_in_3_bits_vc_sel_1_1(salloc_arb_io_in_3_bits_vc_sel_1_1),
    .io_in_3_bits_vc_sel_1_2(salloc_arb_io_in_3_bits_vc_sel_1_2),
    .io_in_3_bits_vc_sel_1_3(salloc_arb_io_in_3_bits_vc_sel_1_3),
    .io_in_3_bits_vc_sel_0_0(salloc_arb_io_in_3_bits_vc_sel_0_0),
    .io_in_3_bits_vc_sel_0_1(salloc_arb_io_in_3_bits_vc_sel_0_1),
    .io_in_3_bits_vc_sel_0_2(salloc_arb_io_in_3_bits_vc_sel_0_2),
    .io_in_3_bits_vc_sel_0_3(salloc_arb_io_in_3_bits_vc_sel_0_3),
    .io_in_3_bits_tail(salloc_arb_io_in_3_bits_tail),
    .io_out_0_ready(salloc_arb_io_out_0_ready),
    .io_out_0_valid(salloc_arb_io_out_0_valid),
    .io_out_0_bits_vc_sel_2_0(salloc_arb_io_out_0_bits_vc_sel_2_0),
    .io_out_0_bits_vc_sel_1_0(salloc_arb_io_out_0_bits_vc_sel_1_0),
    .io_out_0_bits_vc_sel_1_1(salloc_arb_io_out_0_bits_vc_sel_1_1),
    .io_out_0_bits_vc_sel_1_2(salloc_arb_io_out_0_bits_vc_sel_1_2),
    .io_out_0_bits_vc_sel_1_3(salloc_arb_io_out_0_bits_vc_sel_1_3),
    .io_out_0_bits_vc_sel_0_0(salloc_arb_io_out_0_bits_vc_sel_0_0),
    .io_out_0_bits_vc_sel_0_1(salloc_arb_io_out_0_bits_vc_sel_0_1),
    .io_out_0_bits_vc_sel_0_2(salloc_arb_io_out_0_bits_vc_sel_0_2),
    .io_out_0_bits_vc_sel_0_3(salloc_arb_io_out_0_bits_vc_sel_0_3),
    .io_out_0_bits_tail(salloc_arb_io_out_0_bits_tail),
    .io_chosen_oh_0(salloc_arb_io_chosen_oh_0)
  );
  assign io_router_req_valid = route_arbiter_io_out_valid; // @[InputUnit.scala 189:17]
  assign io_router_req_bits_src_virt_id = route_arbiter_io_out_bits_src_virt_id; // @[InputUnit.scala 189:17]
  assign io_router_req_bits_flow_ingress_node = route_arbiter_io_out_bits_flow_ingress_node; // @[InputUnit.scala 189:17]
  assign io_router_req_bits_flow_egress_node = route_arbiter_io_out_bits_flow_egress_node; // @[InputUnit.scala 189:17]
  assign io_vcalloc_req_valid = vcalloc_vals_0 | vcalloc_vals_1 | vcalloc_vals_2 | vcalloc_vals_3; // @[package.scala 73:59]
  assign io_vcalloc_req_bits_vc_sel_2_0 = vcalloc_sel[0] & states_0_vc_sel_2_0 | vcalloc_sel[1] & states_1_vc_sel_2_0 |
    vcalloc_sel[2] & states_2_vc_sel_2_0 | vcalloc_sel[3] & states_3_vc_sel_2_0; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_1_0 = vcalloc_sel[0] & states_0_vc_sel_1_0 | vcalloc_sel[1] & states_1_vc_sel_1_0 |
    vcalloc_sel[2] & states_2_vc_sel_1_0 | vcalloc_sel[3] & states_3_vc_sel_1_0; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_1_1 = vcalloc_sel[2] & states_2_vc_sel_1_1 | vcalloc_sel[3] & states_3_vc_sel_1_1; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_1_2 = vcalloc_sel[3] & states_3_vc_sel_1_2; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_0_0 = vcalloc_sel[0] & states_0_vc_sel_0_0 | vcalloc_sel[1] & states_1_vc_sel_0_0 |
    vcalloc_sel[2] & states_2_vc_sel_0_0 | vcalloc_sel[3] & states_3_vc_sel_0_0; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_0_1 = vcalloc_sel[1] & states_1_vc_sel_0_1 | vcalloc_sel[2] & states_2_vc_sel_0_1 |
    vcalloc_sel[3] & states_3_vc_sel_0_1; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_0_2 = vcalloc_sel[2] & states_2_vc_sel_0_2 | vcalloc_sel[3] & states_3_vc_sel_0_2; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_0_3 = vcalloc_sel[3] & states_3_vc_sel_0_3; // @[Mux.scala 27:73]
  assign io_salloc_req_0_valid = salloc_arb_io_out_0_valid; // @[InputUnit.scala 302:17 303:19 305:35]
  assign io_salloc_req_0_bits_vc_sel_2_0 = salloc_arb_io_out_0_bits_vc_sel_2_0; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_1_0 = salloc_arb_io_out_0_bits_vc_sel_1_0; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_1_1 = salloc_arb_io_out_0_bits_vc_sel_1_1; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_1_2 = salloc_arb_io_out_0_bits_vc_sel_1_2; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_1_3 = salloc_arb_io_out_0_bits_vc_sel_1_3; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_0_0 = salloc_arb_io_out_0_bits_vc_sel_0_0; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_0_1 = salloc_arb_io_out_0_bits_vc_sel_0_1; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_0_2 = salloc_arb_io_out_0_bits_vc_sel_0_2; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_0_3 = salloc_arb_io_out_0_bits_vc_sel_0_3; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_tail = salloc_arb_io_out_0_bits_tail; // @[InputUnit.scala 302:17]
  assign io_out_0_valid = salloc_outs_0_valid; // @[InputUnit.scala 349:21]
  assign io_out_0_bits_flit_head = salloc_outs_0_flit_head; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_flit_tail = salloc_outs_0_flit_tail; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_flit_payload = salloc_outs_0_flit_payload; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_flit_flow_ingress_node = salloc_outs_0_flit_flow_ingress_node; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_flit_flow_egress_node = salloc_outs_0_flit_flow_egress_node; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_out_virt_channel = salloc_outs_0_out_vid; // @[InputUnit.scala 351:37]
  assign io_debug_va_stall = _io_debug_va_stall_T_7[1:0]; // @[InputUnit.scala 266:21]
  assign io_debug_sa_stall = _io_debug_sa_stall_T_12[1:0]; // @[InputUnit.scala 301:21]
  assign io_in_credit_return = _io_in_credit_return_T ? salloc_arb_io_chosen_oh_0 : 4'h0; // @[InputUnit.scala 322:8]
  assign io_in_vc_free = _io_in_credit_return_T & _io_in_vc_free_T_11 ? salloc_arb_io_chosen_oh_0 : 4'h0; // @[InputUnit.scala 325:8]
  assign input_buffer_clock = clock;
  assign input_buffer_reset = reset;
  assign input_buffer_io_enq_0_valid = io_in_flit_0_valid; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_head = io_in_flit_0_bits_head; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_tail = io_in_flit_0_bits_tail; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_payload = io_in_flit_0_bits_payload; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_virt_channel_id = io_in_flit_0_bits_virt_channel_id; // @[InputUnit.scala 182:28]
  assign input_buffer_io_deq_0_ready = salloc_arb_io_in_0_ready; // @[InputUnit.scala 295:36]
  assign input_buffer_io_deq_1_ready = salloc_arb_io_in_1_ready; // @[InputUnit.scala 295:36]
  assign input_buffer_io_deq_2_ready = salloc_arb_io_in_2_ready; // @[InputUnit.scala 295:36]
  assign input_buffer_io_deq_3_ready = salloc_arb_io_in_3_ready; // @[InputUnit.scala 295:36]
  assign route_arbiter_io_in_0_valid = states_0_g == 3'h1; // @[InputUnit.scala 212:22]
  assign route_arbiter_io_in_0_bits_flow_ingress_node = states_0_flow_ingress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_0_bits_flow_egress_node = states_0_flow_egress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_1_valid = states_1_g == 3'h1; // @[InputUnit.scala 212:22]
  assign route_arbiter_io_in_1_bits_flow_ingress_node = states_1_flow_ingress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_1_bits_flow_egress_node = states_1_flow_egress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_2_valid = states_2_g == 3'h1; // @[InputUnit.scala 212:22]
  assign route_arbiter_io_in_2_bits_flow_ingress_node = states_2_flow_ingress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_2_bits_flow_egress_node = states_2_flow_egress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_3_valid = states_3_g == 3'h1; // @[InputUnit.scala 212:22]
  assign route_arbiter_io_in_3_bits_flow_ingress_node = states_3_flow_ingress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_3_bits_flow_egress_node = states_3_flow_egress_node; // @[InputUnit.scala 213:19]
  assign salloc_arb_clock = clock;
  assign salloc_arb_reset = reset;
  assign salloc_arb_io_in_0_valid = states_0_g == 3'h3 & credit_available & input_buffer_io_deq_0_valid; // @[InputUnit.scala 288:50]
  assign salloc_arb_io_in_0_bits_vc_sel_2_0 = states_0_vc_sel_2_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_0_bits_vc_sel_1_0 = states_0_vc_sel_1_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_0_bits_vc_sel_0_0 = states_0_vc_sel_0_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_0_bits_tail = input_buffer_io_deq_0_bits_tail; // @[InputUnit.scala 291:19]
  assign salloc_arb_io_in_1_valid = states_1_g == 3'h3 & credit_available_1 & input_buffer_io_deq_1_valid; // @[InputUnit.scala 288:50]
  assign salloc_arb_io_in_1_bits_vc_sel_2_0 = states_1_vc_sel_2_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_1_bits_vc_sel_1_0 = states_1_vc_sel_1_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_1_bits_vc_sel_1_1 = 1'h0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_1_bits_vc_sel_0_0 = states_1_vc_sel_0_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_1_bits_vc_sel_0_1 = states_1_vc_sel_0_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_1_bits_tail = input_buffer_io_deq_1_bits_tail; // @[InputUnit.scala 291:19]
  assign salloc_arb_io_in_2_valid = states_2_g == 3'h3 & credit_available_2 & input_buffer_io_deq_2_valid; // @[InputUnit.scala 288:50]
  assign salloc_arb_io_in_2_bits_vc_sel_2_0 = states_2_vc_sel_2_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_1_0 = states_2_vc_sel_1_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_1_1 = states_2_vc_sel_1_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_1_2 = 1'h0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_0_0 = states_2_vc_sel_0_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_0_1 = states_2_vc_sel_0_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_0_2 = states_2_vc_sel_0_2; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_tail = input_buffer_io_deq_2_bits_tail; // @[InputUnit.scala 291:19]
  assign salloc_arb_io_in_3_valid = states_3_g == 3'h3 & credit_available_3 & input_buffer_io_deq_3_valid; // @[InputUnit.scala 288:50]
  assign salloc_arb_io_in_3_bits_vc_sel_2_0 = states_3_vc_sel_2_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_1_0 = states_3_vc_sel_1_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_1_1 = states_3_vc_sel_1_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_1_2 = states_3_vc_sel_1_2; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_1_3 = 1'h0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_0_0 = states_3_vc_sel_0_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_0_1 = states_3_vc_sel_0_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_0_2 = states_3_vc_sel_0_2; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_0_3 = states_3_vc_sel_0_3; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_tail = input_buffer_io_deq_3_bits_tail; // @[InputUnit.scala 291:19]
  assign salloc_arb_io_out_0_ready = io_salloc_req_0_ready; // @[InputUnit.scala 302:17 303:19 304:39]
  always @(posedge clock) begin
    if (reset) begin // @[InputUnit.scala 377:23]
      states_0_g <= 3'h0; // @[InputUnit.scala 378:24]
    end else if (_T_60 & input_buffer_io_deq_0_bits_tail) begin // @[InputUnit.scala 292:35]
      states_0_g <= 3'h0; // @[InputUnit.scala 293:13]
    end else if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[0]) begin // @[InputUnit.scala 270:29]
        states_0_g <= 3'h3; // @[InputUnit.scala 272:21]
      end else begin
        states_0_g <= _GEN_222;
      end
    end else begin
      states_0_g <= _GEN_222;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[0]) begin // @[InputUnit.scala 270:29]
        states_0_vc_sel_2_0 <= io_vcalloc_resp_vc_sel_2_0; // @[InputUnit.scala 271:26]
      end else begin
        states_0_vc_sel_2_0 <= _GEN_184;
      end
    end else begin
      states_0_vc_sel_2_0 <= _GEN_184;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[0]) begin // @[InputUnit.scala 270:29]
        states_0_vc_sel_1_0 <= io_vcalloc_resp_vc_sel_1_0; // @[InputUnit.scala 271:26]
      end else begin
        states_0_vc_sel_1_0 <= _GEN_185;
      end
    end else begin
      states_0_vc_sel_1_0 <= _GEN_185;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[0]) begin // @[InputUnit.scala 270:29]
        states_0_vc_sel_0_0 <= io_vcalloc_resp_vc_sel_0_0; // @[InputUnit.scala 271:26]
      end else begin
        states_0_vc_sel_0_0 <= _GEN_189;
      end
    end else begin
      states_0_vc_sel_0_0 <= _GEN_189;
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h0 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_0_flow_ingress_node <= io_in_flit_0_bits_flow_ingress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h0 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_0_flow_egress_node <= io_in_flit_0_bits_flow_egress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (reset) begin // @[InputUnit.scala 377:23]
      states_1_g <= 3'h0; // @[InputUnit.scala 378:24]
    end else if (_T_62 & input_buffer_io_deq_1_bits_tail) begin // @[InputUnit.scala 292:35]
      states_1_g <= 3'h0; // @[InputUnit.scala 293:13]
    end else if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_g <= 3'h3; // @[InputUnit.scala 272:21]
      end else begin
        states_1_g <= _GEN_223;
      end
    end else begin
      states_1_g <= _GEN_223;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_vc_sel_2_0 <= io_vcalloc_resp_vc_sel_2_0; // @[InputUnit.scala 271:26]
      end else begin
        states_1_vc_sel_2_0 <= _GEN_193;
      end
    end else begin
      states_1_vc_sel_2_0 <= _GEN_193;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_vc_sel_1_0 <= io_vcalloc_resp_vc_sel_1_0; // @[InputUnit.scala 271:26]
      end else begin
        states_1_vc_sel_1_0 <= _GEN_194;
      end
    end else begin
      states_1_vc_sel_1_0 <= _GEN_194;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_vc_sel_0_0 <= io_vcalloc_resp_vc_sel_0_0; // @[InputUnit.scala 271:26]
      end else begin
        states_1_vc_sel_0_0 <= _GEN_198;
      end
    end else begin
      states_1_vc_sel_0_0 <= _GEN_198;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_vc_sel_0_1 <= io_vcalloc_resp_vc_sel_0_1; // @[InputUnit.scala 271:26]
      end else begin
        states_1_vc_sel_0_1 <= _GEN_199;
      end
    end else begin
      states_1_vc_sel_0_1 <= _GEN_199;
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h1 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_1_flow_ingress_node <= io_in_flit_0_bits_flow_ingress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h1 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_1_flow_egress_node <= io_in_flit_0_bits_flow_egress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (reset) begin // @[InputUnit.scala 377:23]
      states_2_g <= 3'h0; // @[InputUnit.scala 378:24]
    end else if (_T_64 & input_buffer_io_deq_2_bits_tail) begin // @[InputUnit.scala 292:35]
      states_2_g <= 3'h0; // @[InputUnit.scala 293:13]
    end else if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_g <= 3'h3; // @[InputUnit.scala 272:21]
      end else begin
        states_2_g <= _GEN_224;
      end
    end else begin
      states_2_g <= _GEN_224;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_2_0 <= io_vcalloc_resp_vc_sel_2_0; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_2_0 <= _GEN_202;
      end
    end else begin
      states_2_vc_sel_2_0 <= _GEN_202;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_1_0 <= io_vcalloc_resp_vc_sel_1_0; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_1_0 <= _GEN_203;
      end
    end else begin
      states_2_vc_sel_1_0 <= _GEN_203;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_1_1 <= io_vcalloc_resp_vc_sel_1_1; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_1_1 <= _GEN_204;
      end
    end else begin
      states_2_vc_sel_1_1 <= _GEN_204;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_0_0 <= io_vcalloc_resp_vc_sel_0_0; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_0_0 <= _GEN_207;
      end
    end else begin
      states_2_vc_sel_0_0 <= _GEN_207;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_0_1 <= io_vcalloc_resp_vc_sel_0_1; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_0_1 <= _GEN_208;
      end
    end else begin
      states_2_vc_sel_0_1 <= _GEN_208;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_0_2 <= io_vcalloc_resp_vc_sel_0_2; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_0_2 <= _GEN_209;
      end
    end else begin
      states_2_vc_sel_0_2 <= _GEN_209;
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h2 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_2_flow_ingress_node <= io_in_flit_0_bits_flow_ingress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h2 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_2_flow_egress_node <= io_in_flit_0_bits_flow_egress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (reset) begin // @[InputUnit.scala 377:23]
      states_3_g <= 3'h0; // @[InputUnit.scala 378:24]
    end else if (_T_66 & input_buffer_io_deq_3_bits_tail) begin // @[InputUnit.scala 292:35]
      states_3_g <= 3'h0; // @[InputUnit.scala 293:13]
    end else if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_g <= 3'h3; // @[InputUnit.scala 272:21]
      end else begin
        states_3_g <= _GEN_225;
      end
    end else begin
      states_3_g <= _GEN_225;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_2_0 <= io_vcalloc_resp_vc_sel_2_0; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_2_0 <= _GEN_211;
      end
    end else begin
      states_3_vc_sel_2_0 <= _GEN_211;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_1_0 <= io_vcalloc_resp_vc_sel_1_0; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_1_0 <= _GEN_212;
      end
    end else begin
      states_3_vc_sel_1_0 <= _GEN_212;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_1_1 <= io_vcalloc_resp_vc_sel_1_1; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_1_1 <= _GEN_213;
      end
    end else begin
      states_3_vc_sel_1_1 <= _GEN_213;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_1_2 <= io_vcalloc_resp_vc_sel_1_2; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_1_2 <= _GEN_214;
      end
    end else begin
      states_3_vc_sel_1_2 <= _GEN_214;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_0_0 <= io_vcalloc_resp_vc_sel_0_0; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_0_0 <= _GEN_216;
      end
    end else begin
      states_3_vc_sel_0_0 <= _GEN_216;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_0_1 <= io_vcalloc_resp_vc_sel_0_1; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_0_1 <= _GEN_217;
      end
    end else begin
      states_3_vc_sel_0_1 <= _GEN_217;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_0_2 <= io_vcalloc_resp_vc_sel_0_2; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_0_2 <= _GEN_218;
      end
    end else begin
      states_3_vc_sel_0_2 <= _GEN_218;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_0_3 <= io_vcalloc_resp_vc_sel_0_3; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_0_3 <= _GEN_219;
      end
    end else begin
      states_3_vc_sel_0_3 <= _GEN_219;
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h3 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_3_flow_ingress_node <= io_in_flit_0_bits_flow_ingress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h3 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_3_flow_egress_node <= io_in_flit_0_bits_flow_egress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (reset) begin // @[InputUnit.scala 233:21]
      mask <= 4'h0; // @[InputUnit.scala 233:21]
    end else if (io_router_req_valid) begin // @[InputUnit.scala 239:31]
      mask <= _mask_T_2; // @[InputUnit.scala 240:10]
    end else if (_T_26) begin // @[InputUnit.scala 241:34]
      mask <= _mask_T_17; // @[InputUnit.scala 242:10]
    end
    salloc_outs_0_valid <= salloc_arb_io_out_0_ready & salloc_arb_io_out_0_valid; // @[Decoupled.scala 51:35]
    salloc_outs_0_out_vid <= _virt_channel_T_10 | _virt_channel_T_11; // @[Mux.scala 27:73]
    salloc_outs_0_flit_head <= salloc_arb_io_chosen_oh_0[0] & input_buffer_io_deq_0_bits_head |
      salloc_arb_io_chosen_oh_0[1] & input_buffer_io_deq_1_bits_head | salloc_arb_io_chosen_oh_0[2] &
      input_buffer_io_deq_2_bits_head | salloc_arb_io_chosen_oh_0[3] & input_buffer_io_deq_3_bits_head; // @[Mux.scala 27:73]
    salloc_outs_0_flit_tail <= salloc_arb_io_chosen_oh_0[0] & input_buffer_io_deq_0_bits_tail |
      salloc_arb_io_chosen_oh_0[1] & input_buffer_io_deq_1_bits_tail | salloc_arb_io_chosen_oh_0[2] &
      input_buffer_io_deq_2_bits_tail | salloc_arb_io_chosen_oh_0[3] & input_buffer_io_deq_3_bits_tail; // @[Mux.scala 27:73]
    salloc_outs_0_flit_payload <= _salloc_outs_0_flit_payload_T_9 | _salloc_outs_0_flit_payload_T_7; // @[Mux.scala 27:73]
    salloc_outs_0_flit_flow_ingress_node <= _salloc_outs_0_flit_flow_T_30 | _salloc_outs_0_flit_flow_T_28; // @[Mux.scala 27:73]
    salloc_outs_0_flit_flow_egress_node <= _salloc_outs_0_flit_flow_T_16 | _salloc_outs_0_flit_flow_T_14; // @[Mux.scala 27:73]
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T & _T_3 & ~(_GEN_3 == 3'h0)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:197 assert(states(id).g === g_i)\n"); // @[InputUnit.scala 197:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_router_req_valid & _T_3 & ~(_GEN_139 == 3'h1)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:224 assert(states(id).g === g_r)\n"); // @[InputUnit.scala 224:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_39 & vcalloc_sel[0] & _T_3 & ~vcalloc_vals_0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:274 assert(states(i).g === g_v)\n"); // @[InputUnit.scala 274:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_39 & vcalloc_sel[1] & _T_3 & ~vcalloc_vals_1) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:274 assert(states(i).g === g_v)\n"); // @[InputUnit.scala 274:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_39 & vcalloc_sel[2] & _T_3 & ~vcalloc_vals_2) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:274 assert(states(i).g === g_v)\n"); // @[InputUnit.scala 274:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_39 & vcalloc_sel[3] & _T_3 & ~vcalloc_vals_3) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:274 assert(states(i).g === g_v)\n"); // @[InputUnit.scala 274:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  states_0_g = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  states_0_vc_sel_2_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  states_0_vc_sel_1_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  states_0_vc_sel_0_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  states_0_flow_ingress_node = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  states_0_flow_egress_node = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  states_1_g = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  states_1_vc_sel_2_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  states_1_vc_sel_1_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  states_1_vc_sel_0_0 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  states_1_vc_sel_0_1 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  states_1_flow_ingress_node = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  states_1_flow_egress_node = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  states_2_g = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  states_2_vc_sel_2_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  states_2_vc_sel_1_0 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  states_2_vc_sel_1_1 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  states_2_vc_sel_0_0 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  states_2_vc_sel_0_1 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  states_2_vc_sel_0_2 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  states_2_flow_ingress_node = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  states_2_flow_egress_node = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  states_3_g = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  states_3_vc_sel_2_0 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  states_3_vc_sel_1_0 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  states_3_vc_sel_1_1 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  states_3_vc_sel_1_2 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  states_3_vc_sel_0_0 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  states_3_vc_sel_0_1 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  states_3_vc_sel_0_2 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  states_3_vc_sel_0_3 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  states_3_flow_ingress_node = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  states_3_flow_egress_node = _RAND_32[1:0];
  _RAND_33 = {1{`RANDOM}};
  mask = _RAND_33[3:0];
  _RAND_34 = {1{`RANDOM}};
  salloc_outs_0_valid = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  salloc_outs_0_out_vid = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  salloc_outs_0_flit_head = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  salloc_outs_0_flit_tail = _RAND_37[0:0];
  _RAND_38 = {2{`RANDOM}};
  salloc_outs_0_flit_payload = _RAND_38[63:0];
  _RAND_39 = {1{`RANDOM}};
  salloc_outs_0_flit_flow_ingress_node = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  salloc_outs_0_flit_flow_egress_node = _RAND_40[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (_T & ~reset) begin
      assert(1'h1); // @[InputUnit.scala 196:13]
    end
    //
    if (_T & _T_3) begin
      assert(_GEN_3 == 3'h0); // @[InputUnit.scala 197:13]
    end
    //
    if (io_router_req_valid & _T_3) begin
      assert(_GEN_139 == 3'h1); // @[InputUnit.scala 224:11]
    end
    //
    if (_T_39 & vcalloc_sel[0] & _T_3) begin
      assert(vcalloc_vals_0); // @[InputUnit.scala 274:17]
    end
    //
    if (_T_39 & vcalloc_sel[1] & _T_3) begin
      assert(vcalloc_vals_1); // @[InputUnit.scala 274:17]
    end
    //
    if (_T_39 & vcalloc_sel[2] & _T_3) begin
      assert(vcalloc_vals_2); // @[InputUnit.scala 274:17]
    end
    //
    if (_T_39 & vcalloc_sel[3] & _T_3) begin
      assert(vcalloc_vals_3); // @[InputUnit.scala 274:17]
    end
  end
endmodule
module Queue_8(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_head,
  input         io_enq_bits_tail,
  input  [63:0] io_enq_bits_payload,
  input  [1:0]  io_enq_bits_flow_ingress_node,
  input  [1:0]  io_enq_bits_flow_egress_node,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_head,
  output        io_deq_bits_tail,
  output [63:0] io_deq_bits_payload,
  output [1:0]  io_deq_bits_flow_ingress_node,
  output [1:0]  io_deq_bits_flow_egress_node
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg  ram_head [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_head_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_head_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_head_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_tail [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_tail_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_tail_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_tail_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_en; // @[Decoupled.scala 273:95]
  reg [63:0] ram_payload [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_payload_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_payload_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [63:0] ram_payload_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [63:0] ram_payload_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_payload_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_payload_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_payload_MPORT_en; // @[Decoupled.scala 273:95]
  reg [1:0] ram_flow_ingress_node [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_flow_ingress_node_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_flow_ingress_node_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [1:0] ram_flow_ingress_node_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_flow_ingress_node_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_flow_ingress_node_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_flow_ingress_node_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_flow_ingress_node_MPORT_en; // @[Decoupled.scala 273:95]
  reg [1:0] ram_flow_egress_node [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_flow_egress_node_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_flow_egress_node_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [1:0] ram_flow_egress_node_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_flow_egress_node_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_flow_egress_node_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_flow_egress_node_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_flow_egress_node_MPORT_en; // @[Decoupled.scala 273:95]
  reg  enq_ptr_value; // @[Counter.scala 61:40]
  reg  deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  assign ram_head_io_deq_bits_MPORT_en = 1'h1;
  assign ram_head_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_head_io_deq_bits_MPORT_data = ram_head[ram_head_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_head_MPORT_data = io_enq_bits_head;
  assign ram_head_MPORT_addr = enq_ptr_value;
  assign ram_head_MPORT_mask = 1'h1;
  assign ram_head_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tail_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tail_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_tail_io_deq_bits_MPORT_data = ram_tail[ram_tail_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_tail_MPORT_data = io_enq_bits_tail;
  assign ram_tail_MPORT_addr = enq_ptr_value;
  assign ram_tail_MPORT_mask = 1'h1;
  assign ram_tail_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_payload_io_deq_bits_MPORT_en = 1'h1;
  assign ram_payload_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_payload_io_deq_bits_MPORT_data = ram_payload[ram_payload_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_payload_MPORT_data = io_enq_bits_payload;
  assign ram_payload_MPORT_addr = enq_ptr_value;
  assign ram_payload_MPORT_mask = 1'h1;
  assign ram_payload_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_flow_ingress_node_io_deq_bits_MPORT_en = 1'h1;
  assign ram_flow_ingress_node_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_flow_ingress_node_io_deq_bits_MPORT_data =
    ram_flow_ingress_node[ram_flow_ingress_node_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_flow_ingress_node_MPORT_data = io_enq_bits_flow_ingress_node;
  assign ram_flow_ingress_node_MPORT_addr = enq_ptr_value;
  assign ram_flow_ingress_node_MPORT_mask = 1'h1;
  assign ram_flow_ingress_node_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_flow_egress_node_io_deq_bits_MPORT_en = 1'h1;
  assign ram_flow_egress_node_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_flow_egress_node_io_deq_bits_MPORT_data = ram_flow_egress_node[ram_flow_egress_node_io_deq_bits_MPORT_addr]
    ; // @[Decoupled.scala 273:95]
  assign ram_flow_egress_node_MPORT_data = io_enq_bits_flow_egress_node;
  assign ram_flow_egress_node_MPORT_addr = enq_ptr_value;
  assign ram_flow_egress_node_MPORT_mask = 1'h1;
  assign ram_flow_egress_node_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_head = ram_head_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_tail = ram_tail_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_payload = ram_payload_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_flow_ingress_node = ram_flow_ingress_node_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_flow_egress_node = ram_flow_egress_node_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  always @(posedge clock) begin
    if (ram_head_MPORT_en & ram_head_MPORT_mask) begin
      ram_head[ram_head_MPORT_addr] <= ram_head_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_tail_MPORT_en & ram_tail_MPORT_mask) begin
      ram_tail[ram_tail_MPORT_addr] <= ram_tail_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_payload_MPORT_en & ram_payload_MPORT_mask) begin
      ram_payload[ram_payload_MPORT_addr] <= ram_payload_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_flow_ingress_node_MPORT_en & ram_flow_ingress_node_MPORT_mask) begin
      ram_flow_ingress_node[ram_flow_ingress_node_MPORT_addr] <= ram_flow_ingress_node_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_flow_egress_node_MPORT_en & ram_flow_egress_node_MPORT_mask) begin
      ram_flow_egress_node[ram_flow_egress_node_MPORT_addr] <= ram_flow_egress_node_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_head[initvar] = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_tail[initvar] = _RAND_1[0:0];
  _RAND_2 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload[initvar] = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_flow_ingress_node[initvar] = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_flow_egress_node[initvar] = _RAND_4[1:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  enq_ptr_value = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  deq_ptr_value = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  maybe_full = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_9(
  input   clock,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input   io_enq_bits_vc_sel_2_0,
  input   io_enq_bits_vc_sel_1_0,
  input   io_enq_bits_vc_sel_1_1,
  input   io_enq_bits_vc_sel_1_2,
  input   io_enq_bits_vc_sel_1_3,
  input   io_enq_bits_vc_sel_0_0,
  input   io_enq_bits_vc_sel_0_1,
  input   io_enq_bits_vc_sel_0_2,
  input   io_enq_bits_vc_sel_0_3,
  input   io_deq_ready,
  output  io_deq_valid,
  output  io_deq_bits_vc_sel_2_0,
  output  io_deq_bits_vc_sel_1_0,
  output  io_deq_bits_vc_sel_1_1,
  output  io_deq_bits_vc_sel_1_2,
  output  io_deq_bits_vc_sel_1_3,
  output  io_deq_bits_vc_sel_0_0,
  output  io_deq_bits_vc_sel_0_1,
  output  io_deq_bits_vc_sel_0_2,
  output  io_deq_bits_vc_sel_0_3
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  reg  ram_vc_sel_2_0 [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_2_0_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_2_0_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_2_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_2_0_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_2_0_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_2_0_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_2_0_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_vc_sel_1_0 [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_0_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_0_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_0_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_0_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_0_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_0_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_vc_sel_1_1 [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_1_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_1_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_1_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_1_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_1_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_1_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_vc_sel_1_2 [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_2_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_2_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_2_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_2_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_2_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_2_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_vc_sel_1_3 [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_3_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_3_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_3_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_3_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_3_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_3_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_vc_sel_0_0 [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_0_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_0_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_0_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_0_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_0_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_0_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_vc_sel_0_1 [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_1_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_1_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_1_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_1_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_1_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_1_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_vc_sel_0_2 [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_2_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_2_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_2_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_2_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_2_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_2_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_vc_sel_0_3 [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_3_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_3_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_3_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_3_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_3_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_3_MPORT_en; // @[Decoupled.scala 273:95]
  reg  enq_ptr_value; // @[Counter.scala 61:40]
  reg  deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  assign ram_vc_sel_2_0_io_deq_bits_MPORT_en = 1'h1;
  assign ram_vc_sel_2_0_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_vc_sel_2_0_io_deq_bits_MPORT_data = ram_vc_sel_2_0[ram_vc_sel_2_0_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_vc_sel_2_0_MPORT_data = io_enq_bits_vc_sel_2_0;
  assign ram_vc_sel_2_0_MPORT_addr = enq_ptr_value;
  assign ram_vc_sel_2_0_MPORT_mask = 1'h1;
  assign ram_vc_sel_2_0_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_vc_sel_1_0_io_deq_bits_MPORT_en = 1'h1;
  assign ram_vc_sel_1_0_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_vc_sel_1_0_io_deq_bits_MPORT_data = ram_vc_sel_1_0[ram_vc_sel_1_0_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_vc_sel_1_0_MPORT_data = io_enq_bits_vc_sel_1_0;
  assign ram_vc_sel_1_0_MPORT_addr = enq_ptr_value;
  assign ram_vc_sel_1_0_MPORT_mask = 1'h1;
  assign ram_vc_sel_1_0_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_vc_sel_1_1_io_deq_bits_MPORT_en = 1'h1;
  assign ram_vc_sel_1_1_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_vc_sel_1_1_io_deq_bits_MPORT_data = ram_vc_sel_1_1[ram_vc_sel_1_1_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_vc_sel_1_1_MPORT_data = io_enq_bits_vc_sel_1_1;
  assign ram_vc_sel_1_1_MPORT_addr = enq_ptr_value;
  assign ram_vc_sel_1_1_MPORT_mask = 1'h1;
  assign ram_vc_sel_1_1_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_vc_sel_1_2_io_deq_bits_MPORT_en = 1'h1;
  assign ram_vc_sel_1_2_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_vc_sel_1_2_io_deq_bits_MPORT_data = ram_vc_sel_1_2[ram_vc_sel_1_2_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_vc_sel_1_2_MPORT_data = io_enq_bits_vc_sel_1_2;
  assign ram_vc_sel_1_2_MPORT_addr = enq_ptr_value;
  assign ram_vc_sel_1_2_MPORT_mask = 1'h1;
  assign ram_vc_sel_1_2_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_vc_sel_1_3_io_deq_bits_MPORT_en = 1'h1;
  assign ram_vc_sel_1_3_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_vc_sel_1_3_io_deq_bits_MPORT_data = ram_vc_sel_1_3[ram_vc_sel_1_3_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_vc_sel_1_3_MPORT_data = io_enq_bits_vc_sel_1_3;
  assign ram_vc_sel_1_3_MPORT_addr = enq_ptr_value;
  assign ram_vc_sel_1_3_MPORT_mask = 1'h1;
  assign ram_vc_sel_1_3_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_vc_sel_0_0_io_deq_bits_MPORT_en = 1'h1;
  assign ram_vc_sel_0_0_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_vc_sel_0_0_io_deq_bits_MPORT_data = ram_vc_sel_0_0[ram_vc_sel_0_0_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_vc_sel_0_0_MPORT_data = io_enq_bits_vc_sel_0_0;
  assign ram_vc_sel_0_0_MPORT_addr = enq_ptr_value;
  assign ram_vc_sel_0_0_MPORT_mask = 1'h1;
  assign ram_vc_sel_0_0_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_vc_sel_0_1_io_deq_bits_MPORT_en = 1'h1;
  assign ram_vc_sel_0_1_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_vc_sel_0_1_io_deq_bits_MPORT_data = ram_vc_sel_0_1[ram_vc_sel_0_1_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_vc_sel_0_1_MPORT_data = io_enq_bits_vc_sel_0_1;
  assign ram_vc_sel_0_1_MPORT_addr = enq_ptr_value;
  assign ram_vc_sel_0_1_MPORT_mask = 1'h1;
  assign ram_vc_sel_0_1_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_vc_sel_0_2_io_deq_bits_MPORT_en = 1'h1;
  assign ram_vc_sel_0_2_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_vc_sel_0_2_io_deq_bits_MPORT_data = ram_vc_sel_0_2[ram_vc_sel_0_2_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_vc_sel_0_2_MPORT_data = io_enq_bits_vc_sel_0_2;
  assign ram_vc_sel_0_2_MPORT_addr = enq_ptr_value;
  assign ram_vc_sel_0_2_MPORT_mask = 1'h1;
  assign ram_vc_sel_0_2_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_vc_sel_0_3_io_deq_bits_MPORT_en = 1'h1;
  assign ram_vc_sel_0_3_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_vc_sel_0_3_io_deq_bits_MPORT_data = ram_vc_sel_0_3[ram_vc_sel_0_3_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_vc_sel_0_3_MPORT_data = io_enq_bits_vc_sel_0_3;
  assign ram_vc_sel_0_3_MPORT_addr = enq_ptr_value;
  assign ram_vc_sel_0_3_MPORT_mask = 1'h1;
  assign ram_vc_sel_0_3_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_vc_sel_2_0 = ram_vc_sel_2_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_vc_sel_1_0 = ram_vc_sel_1_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_vc_sel_1_1 = ram_vc_sel_1_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_vc_sel_1_2 = ram_vc_sel_1_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_vc_sel_1_3 = ram_vc_sel_1_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_vc_sel_0_0 = ram_vc_sel_0_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_vc_sel_0_1 = ram_vc_sel_0_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_vc_sel_0_2 = ram_vc_sel_0_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_vc_sel_0_3 = ram_vc_sel_0_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  always @(posedge clock) begin
    if (ram_vc_sel_2_0_MPORT_en & ram_vc_sel_2_0_MPORT_mask) begin
      ram_vc_sel_2_0[ram_vc_sel_2_0_MPORT_addr] <= ram_vc_sel_2_0_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_vc_sel_1_0_MPORT_en & ram_vc_sel_1_0_MPORT_mask) begin
      ram_vc_sel_1_0[ram_vc_sel_1_0_MPORT_addr] <= ram_vc_sel_1_0_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_vc_sel_1_1_MPORT_en & ram_vc_sel_1_1_MPORT_mask) begin
      ram_vc_sel_1_1[ram_vc_sel_1_1_MPORT_addr] <= ram_vc_sel_1_1_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_vc_sel_1_2_MPORT_en & ram_vc_sel_1_2_MPORT_mask) begin
      ram_vc_sel_1_2[ram_vc_sel_1_2_MPORT_addr] <= ram_vc_sel_1_2_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_vc_sel_1_3_MPORT_en & ram_vc_sel_1_3_MPORT_mask) begin
      ram_vc_sel_1_3[ram_vc_sel_1_3_MPORT_addr] <= ram_vc_sel_1_3_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_vc_sel_0_0_MPORT_en & ram_vc_sel_0_0_MPORT_mask) begin
      ram_vc_sel_0_0[ram_vc_sel_0_0_MPORT_addr] <= ram_vc_sel_0_0_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_vc_sel_0_1_MPORT_en & ram_vc_sel_0_1_MPORT_mask) begin
      ram_vc_sel_0_1[ram_vc_sel_0_1_MPORT_addr] <= ram_vc_sel_0_1_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_vc_sel_0_2_MPORT_en & ram_vc_sel_0_2_MPORT_mask) begin
      ram_vc_sel_0_2[ram_vc_sel_0_2_MPORT_addr] <= ram_vc_sel_0_2_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_vc_sel_0_3_MPORT_en & ram_vc_sel_0_3_MPORT_mask) begin
      ram_vc_sel_0_3[ram_vc_sel_0_3_MPORT_addr] <= ram_vc_sel_0_3_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_vc_sel_2_0[initvar] = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_vc_sel_1_0[initvar] = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_vc_sel_1_1[initvar] = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_vc_sel_1_2[initvar] = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_vc_sel_1_3[initvar] = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_vc_sel_0_0[initvar] = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_vc_sel_0_1[initvar] = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_vc_sel_0_2[initvar] = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_vc_sel_0_3[initvar] = _RAND_8[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  enq_ptr_value = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  deq_ptr_value = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  maybe_full = _RAND_11[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_11(
  input   clock,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input   io_enq_bits_vc_sel_2_0,
  input   io_enq_bits_vc_sel_1_0,
  input   io_enq_bits_vc_sel_1_1,
  input   io_enq_bits_vc_sel_1_2,
  input   io_enq_bits_vc_sel_1_3,
  input   io_enq_bits_vc_sel_0_0,
  input   io_enq_bits_vc_sel_0_1,
  input   io_enq_bits_vc_sel_0_2,
  input   io_enq_bits_vc_sel_0_3,
  input   io_deq_ready,
  output  io_deq_valid,
  output  io_deq_bits_vc_sel_2_0,
  output  io_deq_bits_vc_sel_1_0,
  output  io_deq_bits_vc_sel_1_1,
  output  io_deq_bits_vc_sel_1_2,
  output  io_deq_bits_vc_sel_1_3,
  output  io_deq_bits_vc_sel_0_0,
  output  io_deq_bits_vc_sel_0_1,
  output  io_deq_bits_vc_sel_0_2,
  output  io_deq_bits_vc_sel_0_3
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  reg  ram_vc_sel_2_0 [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_2_0_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_2_0_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_2_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_2_0_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_2_0_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_2_0_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_2_0_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_vc_sel_1_0 [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_0_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_0_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_0_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_0_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_0_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_0_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_vc_sel_1_1 [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_1_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_1_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_1_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_1_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_1_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_1_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_vc_sel_1_2 [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_2_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_2_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_2_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_2_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_2_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_2_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_vc_sel_1_3 [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_3_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_3_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_3_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_3_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_3_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_3_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_vc_sel_0_0 [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_0_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_0_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_0_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_0_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_0_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_0_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_vc_sel_0_1 [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_1_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_1_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_1_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_1_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_1_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_1_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_vc_sel_0_2 [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_2_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_2_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_2_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_2_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_2_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_2_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_vc_sel_0_3 [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_3_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_3_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_3_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_3_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_3_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_3_MPORT_en; // @[Decoupled.scala 273:95]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 278:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  assign ram_vc_sel_2_0_io_deq_bits_MPORT_en = 1'h1;
  assign ram_vc_sel_2_0_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_vc_sel_2_0_io_deq_bits_MPORT_data = ram_vc_sel_2_0[ram_vc_sel_2_0_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_vc_sel_2_0_MPORT_data = io_enq_bits_vc_sel_2_0;
  assign ram_vc_sel_2_0_MPORT_addr = 1'h0;
  assign ram_vc_sel_2_0_MPORT_mask = 1'h1;
  assign ram_vc_sel_2_0_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_vc_sel_1_0_io_deq_bits_MPORT_en = 1'h1;
  assign ram_vc_sel_1_0_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_vc_sel_1_0_io_deq_bits_MPORT_data = ram_vc_sel_1_0[ram_vc_sel_1_0_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_vc_sel_1_0_MPORT_data = io_enq_bits_vc_sel_1_0;
  assign ram_vc_sel_1_0_MPORT_addr = 1'h0;
  assign ram_vc_sel_1_0_MPORT_mask = 1'h1;
  assign ram_vc_sel_1_0_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_vc_sel_1_1_io_deq_bits_MPORT_en = 1'h1;
  assign ram_vc_sel_1_1_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_vc_sel_1_1_io_deq_bits_MPORT_data = ram_vc_sel_1_1[ram_vc_sel_1_1_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_vc_sel_1_1_MPORT_data = io_enq_bits_vc_sel_1_1;
  assign ram_vc_sel_1_1_MPORT_addr = 1'h0;
  assign ram_vc_sel_1_1_MPORT_mask = 1'h1;
  assign ram_vc_sel_1_1_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_vc_sel_1_2_io_deq_bits_MPORT_en = 1'h1;
  assign ram_vc_sel_1_2_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_vc_sel_1_2_io_deq_bits_MPORT_data = ram_vc_sel_1_2[ram_vc_sel_1_2_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_vc_sel_1_2_MPORT_data = io_enq_bits_vc_sel_1_2;
  assign ram_vc_sel_1_2_MPORT_addr = 1'h0;
  assign ram_vc_sel_1_2_MPORT_mask = 1'h1;
  assign ram_vc_sel_1_2_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_vc_sel_1_3_io_deq_bits_MPORT_en = 1'h1;
  assign ram_vc_sel_1_3_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_vc_sel_1_3_io_deq_bits_MPORT_data = ram_vc_sel_1_3[ram_vc_sel_1_3_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_vc_sel_1_3_MPORT_data = io_enq_bits_vc_sel_1_3;
  assign ram_vc_sel_1_3_MPORT_addr = 1'h0;
  assign ram_vc_sel_1_3_MPORT_mask = 1'h1;
  assign ram_vc_sel_1_3_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_vc_sel_0_0_io_deq_bits_MPORT_en = 1'h1;
  assign ram_vc_sel_0_0_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_vc_sel_0_0_io_deq_bits_MPORT_data = ram_vc_sel_0_0[ram_vc_sel_0_0_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_vc_sel_0_0_MPORT_data = io_enq_bits_vc_sel_0_0;
  assign ram_vc_sel_0_0_MPORT_addr = 1'h0;
  assign ram_vc_sel_0_0_MPORT_mask = 1'h1;
  assign ram_vc_sel_0_0_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_vc_sel_0_1_io_deq_bits_MPORT_en = 1'h1;
  assign ram_vc_sel_0_1_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_vc_sel_0_1_io_deq_bits_MPORT_data = ram_vc_sel_0_1[ram_vc_sel_0_1_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_vc_sel_0_1_MPORT_data = io_enq_bits_vc_sel_0_1;
  assign ram_vc_sel_0_1_MPORT_addr = 1'h0;
  assign ram_vc_sel_0_1_MPORT_mask = 1'h1;
  assign ram_vc_sel_0_1_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_vc_sel_0_2_io_deq_bits_MPORT_en = 1'h1;
  assign ram_vc_sel_0_2_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_vc_sel_0_2_io_deq_bits_MPORT_data = ram_vc_sel_0_2[ram_vc_sel_0_2_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_vc_sel_0_2_MPORT_data = io_enq_bits_vc_sel_0_2;
  assign ram_vc_sel_0_2_MPORT_addr = 1'h0;
  assign ram_vc_sel_0_2_MPORT_mask = 1'h1;
  assign ram_vc_sel_0_2_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_vc_sel_0_3_io_deq_bits_MPORT_en = 1'h1;
  assign ram_vc_sel_0_3_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_vc_sel_0_3_io_deq_bits_MPORT_data = ram_vc_sel_0_3[ram_vc_sel_0_3_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_vc_sel_0_3_MPORT_data = io_enq_bits_vc_sel_0_3;
  assign ram_vc_sel_0_3_MPORT_addr = 1'h0;
  assign ram_vc_sel_0_3_MPORT_mask = 1'h1;
  assign ram_vc_sel_0_3_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = io_deq_ready | empty; // @[Decoupled.scala 303:16 323:{24,39}]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_vc_sel_2_0 = ram_vc_sel_2_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_vc_sel_1_0 = ram_vc_sel_1_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_vc_sel_1_1 = ram_vc_sel_1_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_vc_sel_1_2 = ram_vc_sel_1_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_vc_sel_1_3 = ram_vc_sel_1_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_vc_sel_0_0 = ram_vc_sel_0_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_vc_sel_0_1 = ram_vc_sel_0_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_vc_sel_0_2 = ram_vc_sel_0_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_vc_sel_0_3 = ram_vc_sel_0_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  always @(posedge clock) begin
    if (ram_vc_sel_2_0_MPORT_en & ram_vc_sel_2_0_MPORT_mask) begin
      ram_vc_sel_2_0[ram_vc_sel_2_0_MPORT_addr] <= ram_vc_sel_2_0_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_vc_sel_1_0_MPORT_en & ram_vc_sel_1_0_MPORT_mask) begin
      ram_vc_sel_1_0[ram_vc_sel_1_0_MPORT_addr] <= ram_vc_sel_1_0_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_vc_sel_1_1_MPORT_en & ram_vc_sel_1_1_MPORT_mask) begin
      ram_vc_sel_1_1[ram_vc_sel_1_1_MPORT_addr] <= ram_vc_sel_1_1_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_vc_sel_1_2_MPORT_en & ram_vc_sel_1_2_MPORT_mask) begin
      ram_vc_sel_1_2[ram_vc_sel_1_2_MPORT_addr] <= ram_vc_sel_1_2_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_vc_sel_1_3_MPORT_en & ram_vc_sel_1_3_MPORT_mask) begin
      ram_vc_sel_1_3[ram_vc_sel_1_3_MPORT_addr] <= ram_vc_sel_1_3_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_vc_sel_0_0_MPORT_en & ram_vc_sel_0_0_MPORT_mask) begin
      ram_vc_sel_0_0[ram_vc_sel_0_0_MPORT_addr] <= ram_vc_sel_0_0_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_vc_sel_0_1_MPORT_en & ram_vc_sel_0_1_MPORT_mask) begin
      ram_vc_sel_0_1[ram_vc_sel_0_1_MPORT_addr] <= ram_vc_sel_0_1_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_vc_sel_0_2_MPORT_en & ram_vc_sel_0_2_MPORT_mask) begin
      ram_vc_sel_0_2[ram_vc_sel_0_2_MPORT_addr] <= ram_vc_sel_0_2_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_vc_sel_0_3_MPORT_en & ram_vc_sel_0_3_MPORT_mask) begin
      ram_vc_sel_0_3[ram_vc_sel_0_3_MPORT_addr] <= ram_vc_sel_0_3_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_vc_sel_2_0[initvar] = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_vc_sel_1_0[initvar] = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_vc_sel_1_1[initvar] = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_vc_sel_1_2[initvar] = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_vc_sel_1_3[initvar] = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_vc_sel_0_0[initvar] = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_vc_sel_0_1[initvar] = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_vc_sel_0_2[initvar] = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_vc_sel_0_3[initvar] = _RAND_8[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  maybe_full = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IngressUnit(
  input         clock,
  input         reset,
  output        io_router_req_valid,
  output [1:0]  io_router_req_bits_flow_ingress_node,
  output [1:0]  io_router_req_bits_flow_egress_node,
  input         io_router_resp_vc_sel_1_0,
  input         io_router_resp_vc_sel_1_1,
  input         io_router_resp_vc_sel_1_2,
  input         io_router_resp_vc_sel_1_3,
  input         io_router_resp_vc_sel_0_0,
  input         io_router_resp_vc_sel_0_1,
  input         io_router_resp_vc_sel_0_2,
  input         io_router_resp_vc_sel_0_3,
  input         io_vcalloc_req_ready,
  output        io_vcalloc_req_valid,
  output        io_vcalloc_req_bits_vc_sel_2_0,
  output        io_vcalloc_req_bits_vc_sel_1_0,
  output        io_vcalloc_req_bits_vc_sel_1_1,
  output        io_vcalloc_req_bits_vc_sel_1_2,
  output        io_vcalloc_req_bits_vc_sel_1_3,
  output        io_vcalloc_req_bits_vc_sel_0_0,
  output        io_vcalloc_req_bits_vc_sel_0_1,
  output        io_vcalloc_req_bits_vc_sel_0_2,
  output        io_vcalloc_req_bits_vc_sel_0_3,
  input         io_vcalloc_resp_vc_sel_2_0,
  input         io_vcalloc_resp_vc_sel_1_0,
  input         io_vcalloc_resp_vc_sel_1_1,
  input         io_vcalloc_resp_vc_sel_1_2,
  input         io_vcalloc_resp_vc_sel_1_3,
  input         io_vcalloc_resp_vc_sel_0_0,
  input         io_vcalloc_resp_vc_sel_0_1,
  input         io_vcalloc_resp_vc_sel_0_2,
  input         io_vcalloc_resp_vc_sel_0_3,
  input         io_out_credit_available_2_0,
  input         io_out_credit_available_1_0,
  input         io_out_credit_available_1_1,
  input         io_out_credit_available_1_2,
  input         io_out_credit_available_1_3,
  input         io_out_credit_available_0_0,
  input         io_out_credit_available_0_1,
  input         io_out_credit_available_0_2,
  input         io_out_credit_available_0_3,
  input         io_salloc_req_0_ready,
  output        io_salloc_req_0_valid,
  output        io_salloc_req_0_bits_vc_sel_2_0,
  output        io_salloc_req_0_bits_vc_sel_1_0,
  output        io_salloc_req_0_bits_vc_sel_1_1,
  output        io_salloc_req_0_bits_vc_sel_1_2,
  output        io_salloc_req_0_bits_vc_sel_1_3,
  output        io_salloc_req_0_bits_vc_sel_0_0,
  output        io_salloc_req_0_bits_vc_sel_0_1,
  output        io_salloc_req_0_bits_vc_sel_0_2,
  output        io_salloc_req_0_bits_vc_sel_0_3,
  output        io_salloc_req_0_bits_tail,
  output        io_out_0_valid,
  output        io_out_0_bits_flit_head,
  output        io_out_0_bits_flit_tail,
  output [63:0] io_out_0_bits_flit_payload,
  output [1:0]  io_out_0_bits_flit_flow_ingress_node,
  output [1:0]  io_out_0_bits_flit_flow_egress_node,
  output [1:0]  io_out_0_bits_out_virt_channel,
  output        io_in_ready,
  input         io_in_valid,
  input         io_in_bits_head,
  input         io_in_bits_tail,
  input  [63:0] io_in_bits_payload,
  input  [1:0]  io_in_bits_egress_id
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  route_buffer_clock; // @[IngressUnit.scala 26:28]
  wire  route_buffer_reset; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_enq_ready; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_enq_valid; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_enq_bits_head; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_enq_bits_tail; // @[IngressUnit.scala 26:28]
  wire [63:0] route_buffer_io_enq_bits_payload; // @[IngressUnit.scala 26:28]
  wire [1:0] route_buffer_io_enq_bits_flow_ingress_node; // @[IngressUnit.scala 26:28]
  wire [1:0] route_buffer_io_enq_bits_flow_egress_node; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_deq_ready; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_deq_valid; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_deq_bits_head; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_deq_bits_tail; // @[IngressUnit.scala 26:28]
  wire [63:0] route_buffer_io_deq_bits_payload; // @[IngressUnit.scala 26:28]
  wire [1:0] route_buffer_io_deq_bits_flow_ingress_node; // @[IngressUnit.scala 26:28]
  wire [1:0] route_buffer_io_deq_bits_flow_egress_node; // @[IngressUnit.scala 26:28]
  wire  route_q_clock; // @[IngressUnit.scala 27:23]
  wire  route_q_reset; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_ready; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_valid; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_2_0; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_1_0; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_1_1; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_1_2; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_1_3; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_0_0; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_0_1; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_0_2; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_0_3; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_ready; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_valid; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_2_0; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_1_0; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_1_1; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_1_2; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_1_3; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_0_0; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_0_1; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_0_2; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_0_3; // @[IngressUnit.scala 27:23]
  wire  vcalloc_buffer_clock; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_reset; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_enq_ready; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_enq_valid; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_enq_bits_head; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_enq_bits_tail; // @[IngressUnit.scala 75:30]
  wire [63:0] vcalloc_buffer_io_enq_bits_payload; // @[IngressUnit.scala 75:30]
  wire [1:0] vcalloc_buffer_io_enq_bits_flow_ingress_node; // @[IngressUnit.scala 75:30]
  wire [1:0] vcalloc_buffer_io_enq_bits_flow_egress_node; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_deq_ready; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_deq_valid; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_deq_bits_head; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_deq_bits_tail; // @[IngressUnit.scala 75:30]
  wire [63:0] vcalloc_buffer_io_deq_bits_payload; // @[IngressUnit.scala 75:30]
  wire [1:0] vcalloc_buffer_io_deq_bits_flow_ingress_node; // @[IngressUnit.scala 75:30]
  wire [1:0] vcalloc_buffer_io_deq_bits_flow_egress_node; // @[IngressUnit.scala 75:30]
  wire  vcalloc_q_clock; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_reset; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_ready; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_valid; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_2_0; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_1_0; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_1_1; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_1_2; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_1_3; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_0_0; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_0_1; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_0_2; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_0_3; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_ready; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_valid; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_2_0; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_1_0; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_1_1; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_1_2; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_1_3; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_0_0; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_0_1; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_0_2; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_0_3; // @[IngressUnit.scala 76:25]
  wire  _T = 2'h0 == io_in_bits_egress_id; // @[IngressUnit.scala 30:72]
  wire  _T_1 = 2'h1 == io_in_bits_egress_id; // @[IngressUnit.scala 30:72]
  wire  _T_2 = 2'h2 == io_in_bits_egress_id; // @[IngressUnit.scala 30:72]
  wire  _T_3 = 2'h3 == io_in_bits_egress_id; // @[IngressUnit.scala 30:72]
  wire  _T_6 = _T | _T_1 | _T_2 | _T_3; // @[package.scala 73:59]
  wire  _T_11 = ~reset; // @[IngressUnit.scala 30:9]
  wire [1:0] _route_buffer_io_enq_bits_flow_egress_node_T_6 = _T_2 ? 2'h2 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _route_buffer_io_enq_bits_flow_egress_node_T_7 = _T_3 ? 2'h3 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _GEN_11 = {{1'd0}, _T_1}; // @[Mux.scala 27:73]
  wire [1:0] _route_buffer_io_enq_bits_flow_egress_node_T_9 = _GEN_11 | _route_buffer_io_enq_bits_flow_egress_node_T_6; // @[Mux.scala 27:73]
  wire  at_dest = route_buffer_io_enq_bits_flow_egress_node == 2'h0; // @[IngressUnit.scala 55:59]
  wire  _T_13 = io_in_ready & io_in_valid; // @[Decoupled.scala 51:35]
  wire  _vcalloc_buffer_io_enq_valid_T = ~route_buffer_io_deq_bits_head; // @[IngressUnit.scala 88:30]
  wire  _vcalloc_buffer_io_enq_valid_T_1 = route_q_io_deq_valid | ~route_buffer_io_deq_bits_head; // @[IngressUnit.scala 88:27]
  wire  _vcalloc_buffer_io_enq_valid_T_2 = route_buffer_io_deq_valid & _vcalloc_buffer_io_enq_valid_T_1; // @[IngressUnit.scala 87:61]
  wire  _vcalloc_buffer_io_enq_valid_T_4 = io_vcalloc_req_ready | _vcalloc_buffer_io_enq_valid_T; // @[IngressUnit.scala 89:27]
  wire  _io_vcalloc_req_valid_T_1 = route_buffer_io_deq_valid & route_q_io_deq_valid & route_buffer_io_deq_bits_head; // @[IngressUnit.scala 91:78]
  wire  _route_buffer_io_deq_ready_T_2 = vcalloc_buffer_io_enq_ready & _vcalloc_buffer_io_enq_valid_T_1; // @[IngressUnit.scala 93:61]
  wire  _route_buffer_io_deq_ready_T_5 = _route_buffer_io_deq_ready_T_2 & _vcalloc_buffer_io_enq_valid_T_4; // @[IngressUnit.scala 94:37]
  wire  _route_buffer_io_deq_ready_T_7 = vcalloc_q_io_enq_ready | _vcalloc_buffer_io_enq_valid_T; // @[IngressUnit.scala 96:29]
  wire  _route_q_io_deq_ready_T = route_buffer_io_deq_ready & route_buffer_io_deq_valid; // @[Decoupled.scala 51:35]
  wire [3:0] c_lo = {vcalloc_q_io_deq_bits_vc_sel_0_3,vcalloc_q_io_deq_bits_vc_sel_0_2,vcalloc_q_io_deq_bits_vc_sel_0_1,
    vcalloc_q_io_deq_bits_vc_sel_0_0}; // @[IngressUnit.scala 107:41]
  wire [8:0] _c_T = {vcalloc_q_io_deq_bits_vc_sel_2_0,vcalloc_q_io_deq_bits_vc_sel_1_3,vcalloc_q_io_deq_bits_vc_sel_1_2,
    vcalloc_q_io_deq_bits_vc_sel_1_1,vcalloc_q_io_deq_bits_vc_sel_1_0,vcalloc_q_io_deq_bits_vc_sel_0_3,
    vcalloc_q_io_deq_bits_vc_sel_0_2,vcalloc_q_io_deq_bits_vc_sel_0_1,vcalloc_q_io_deq_bits_vc_sel_0_0}; // @[IngressUnit.scala 107:41]
  wire [8:0] _c_T_1 = {io_out_credit_available_2_0,io_out_credit_available_1_3,io_out_credit_available_1_2,
    io_out_credit_available_1_1,io_out_credit_available_1_0,io_out_credit_available_0_3,io_out_credit_available_0_2,
    io_out_credit_available_0_1,io_out_credit_available_0_0}; // @[IngressUnit.scala 107:74]
  wire [8:0] _c_T_2 = _c_T & _c_T_1; // @[IngressUnit.scala 107:48]
  wire  c = _c_T_2 != 9'h0; // @[IngressUnit.scala 107:82]
  wire  _vcalloc_q_io_deq_ready_T = vcalloc_buffer_io_deq_ready & vcalloc_buffer_io_deq_valid; // @[Decoupled.scala 51:35]
  reg  out_bundle_valid; // @[IngressUnit.scala 116:8]
  reg  out_bundle_bits_flit_head; // @[IngressUnit.scala 116:8]
  reg  out_bundle_bits_flit_tail; // @[IngressUnit.scala 116:8]
  reg [63:0] out_bundle_bits_flit_payload; // @[IngressUnit.scala 116:8]
  reg [1:0] out_bundle_bits_flit_flow_ingress_node; // @[IngressUnit.scala 116:8]
  reg [1:0] out_bundle_bits_flit_flow_egress_node; // @[IngressUnit.scala 116:8]
  reg [1:0] out_bundle_bits_out_virt_channel; // @[IngressUnit.scala 116:8]
  wire  out_channel_oh_0 = vcalloc_q_io_deq_bits_vc_sel_0_0 | vcalloc_q_io_deq_bits_vc_sel_0_1 |
    vcalloc_q_io_deq_bits_vc_sel_0_2 | vcalloc_q_io_deq_bits_vc_sel_0_3; // @[IngressUnit.scala 123:67]
  wire  out_channel_oh_1 = vcalloc_q_io_deq_bits_vc_sel_1_0 | vcalloc_q_io_deq_bits_vc_sel_1_1 |
    vcalloc_q_io_deq_bits_vc_sel_1_2 | vcalloc_q_io_deq_bits_vc_sel_1_3; // @[IngressUnit.scala 123:67]
  wire [1:0] out_bundle_bits_out_virt_channel_hi_1 = c_lo[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] out_bundle_bits_out_virt_channel_lo_1 = c_lo[1:0]; // @[OneHot.scala 31:18]
  wire  _out_bundle_bits_out_virt_channel_T_1 = |out_bundle_bits_out_virt_channel_hi_1; // @[OneHot.scala 32:14]
  wire [1:0] _out_bundle_bits_out_virt_channel_T_2 = out_bundle_bits_out_virt_channel_hi_1 |
    out_bundle_bits_out_virt_channel_lo_1; // @[OneHot.scala 32:28]
  wire [1:0] _out_bundle_bits_out_virt_channel_T_4 = {_out_bundle_bits_out_virt_channel_T_1,
    _out_bundle_bits_out_virt_channel_T_2[1]}; // @[Cat.scala 33:92]
  wire [3:0] _out_bundle_bits_out_virt_channel_T_5 = {vcalloc_q_io_deq_bits_vc_sel_1_3,vcalloc_q_io_deq_bits_vc_sel_1_2,
    vcalloc_q_io_deq_bits_vc_sel_1_1,vcalloc_q_io_deq_bits_vc_sel_1_0}; // @[OneHot.scala 22:45]
  wire [1:0] out_bundle_bits_out_virt_channel_hi_3 = _out_bundle_bits_out_virt_channel_T_5[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] out_bundle_bits_out_virt_channel_lo_3 = _out_bundle_bits_out_virt_channel_T_5[1:0]; // @[OneHot.scala 31:18]
  wire  _out_bundle_bits_out_virt_channel_T_6 = |out_bundle_bits_out_virt_channel_hi_3; // @[OneHot.scala 32:14]
  wire [1:0] _out_bundle_bits_out_virt_channel_T_7 = out_bundle_bits_out_virt_channel_hi_3 |
    out_bundle_bits_out_virt_channel_lo_3; // @[OneHot.scala 32:28]
  wire [1:0] _out_bundle_bits_out_virt_channel_T_9 = {_out_bundle_bits_out_virt_channel_T_6,
    _out_bundle_bits_out_virt_channel_T_7[1]}; // @[Cat.scala 33:92]
  wire [1:0] _out_bundle_bits_out_virt_channel_T_10 = out_channel_oh_0 ? _out_bundle_bits_out_virt_channel_T_4 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _out_bundle_bits_out_virt_channel_T_11 = out_channel_oh_1 ? _out_bundle_bits_out_virt_channel_T_9 : 2'h0; // @[Mux.scala 27:73]
  Queue_8 route_buffer ( // @[IngressUnit.scala 26:28]
    .clock(route_buffer_clock),
    .reset(route_buffer_reset),
    .io_enq_ready(route_buffer_io_enq_ready),
    .io_enq_valid(route_buffer_io_enq_valid),
    .io_enq_bits_head(route_buffer_io_enq_bits_head),
    .io_enq_bits_tail(route_buffer_io_enq_bits_tail),
    .io_enq_bits_payload(route_buffer_io_enq_bits_payload),
    .io_enq_bits_flow_ingress_node(route_buffer_io_enq_bits_flow_ingress_node),
    .io_enq_bits_flow_egress_node(route_buffer_io_enq_bits_flow_egress_node),
    .io_deq_ready(route_buffer_io_deq_ready),
    .io_deq_valid(route_buffer_io_deq_valid),
    .io_deq_bits_head(route_buffer_io_deq_bits_head),
    .io_deq_bits_tail(route_buffer_io_deq_bits_tail),
    .io_deq_bits_payload(route_buffer_io_deq_bits_payload),
    .io_deq_bits_flow_ingress_node(route_buffer_io_deq_bits_flow_ingress_node),
    .io_deq_bits_flow_egress_node(route_buffer_io_deq_bits_flow_egress_node)
  );
  Queue_9 route_q ( // @[IngressUnit.scala 27:23]
    .clock(route_q_clock),
    .reset(route_q_reset),
    .io_enq_ready(route_q_io_enq_ready),
    .io_enq_valid(route_q_io_enq_valid),
    .io_enq_bits_vc_sel_2_0(route_q_io_enq_bits_vc_sel_2_0),
    .io_enq_bits_vc_sel_1_0(route_q_io_enq_bits_vc_sel_1_0),
    .io_enq_bits_vc_sel_1_1(route_q_io_enq_bits_vc_sel_1_1),
    .io_enq_bits_vc_sel_1_2(route_q_io_enq_bits_vc_sel_1_2),
    .io_enq_bits_vc_sel_1_3(route_q_io_enq_bits_vc_sel_1_3),
    .io_enq_bits_vc_sel_0_0(route_q_io_enq_bits_vc_sel_0_0),
    .io_enq_bits_vc_sel_0_1(route_q_io_enq_bits_vc_sel_0_1),
    .io_enq_bits_vc_sel_0_2(route_q_io_enq_bits_vc_sel_0_2),
    .io_enq_bits_vc_sel_0_3(route_q_io_enq_bits_vc_sel_0_3),
    .io_deq_ready(route_q_io_deq_ready),
    .io_deq_valid(route_q_io_deq_valid),
    .io_deq_bits_vc_sel_2_0(route_q_io_deq_bits_vc_sel_2_0),
    .io_deq_bits_vc_sel_1_0(route_q_io_deq_bits_vc_sel_1_0),
    .io_deq_bits_vc_sel_1_1(route_q_io_deq_bits_vc_sel_1_1),
    .io_deq_bits_vc_sel_1_2(route_q_io_deq_bits_vc_sel_1_2),
    .io_deq_bits_vc_sel_1_3(route_q_io_deq_bits_vc_sel_1_3),
    .io_deq_bits_vc_sel_0_0(route_q_io_deq_bits_vc_sel_0_0),
    .io_deq_bits_vc_sel_0_1(route_q_io_deq_bits_vc_sel_0_1),
    .io_deq_bits_vc_sel_0_2(route_q_io_deq_bits_vc_sel_0_2),
    .io_deq_bits_vc_sel_0_3(route_q_io_deq_bits_vc_sel_0_3)
  );
  Queue_8 vcalloc_buffer ( // @[IngressUnit.scala 75:30]
    .clock(vcalloc_buffer_clock),
    .reset(vcalloc_buffer_reset),
    .io_enq_ready(vcalloc_buffer_io_enq_ready),
    .io_enq_valid(vcalloc_buffer_io_enq_valid),
    .io_enq_bits_head(vcalloc_buffer_io_enq_bits_head),
    .io_enq_bits_tail(vcalloc_buffer_io_enq_bits_tail),
    .io_enq_bits_payload(vcalloc_buffer_io_enq_bits_payload),
    .io_enq_bits_flow_ingress_node(vcalloc_buffer_io_enq_bits_flow_ingress_node),
    .io_enq_bits_flow_egress_node(vcalloc_buffer_io_enq_bits_flow_egress_node),
    .io_deq_ready(vcalloc_buffer_io_deq_ready),
    .io_deq_valid(vcalloc_buffer_io_deq_valid),
    .io_deq_bits_head(vcalloc_buffer_io_deq_bits_head),
    .io_deq_bits_tail(vcalloc_buffer_io_deq_bits_tail),
    .io_deq_bits_payload(vcalloc_buffer_io_deq_bits_payload),
    .io_deq_bits_flow_ingress_node(vcalloc_buffer_io_deq_bits_flow_ingress_node),
    .io_deq_bits_flow_egress_node(vcalloc_buffer_io_deq_bits_flow_egress_node)
  );
  Queue_11 vcalloc_q ( // @[IngressUnit.scala 76:25]
    .clock(vcalloc_q_clock),
    .reset(vcalloc_q_reset),
    .io_enq_ready(vcalloc_q_io_enq_ready),
    .io_enq_valid(vcalloc_q_io_enq_valid),
    .io_enq_bits_vc_sel_2_0(vcalloc_q_io_enq_bits_vc_sel_2_0),
    .io_enq_bits_vc_sel_1_0(vcalloc_q_io_enq_bits_vc_sel_1_0),
    .io_enq_bits_vc_sel_1_1(vcalloc_q_io_enq_bits_vc_sel_1_1),
    .io_enq_bits_vc_sel_1_2(vcalloc_q_io_enq_bits_vc_sel_1_2),
    .io_enq_bits_vc_sel_1_3(vcalloc_q_io_enq_bits_vc_sel_1_3),
    .io_enq_bits_vc_sel_0_0(vcalloc_q_io_enq_bits_vc_sel_0_0),
    .io_enq_bits_vc_sel_0_1(vcalloc_q_io_enq_bits_vc_sel_0_1),
    .io_enq_bits_vc_sel_0_2(vcalloc_q_io_enq_bits_vc_sel_0_2),
    .io_enq_bits_vc_sel_0_3(vcalloc_q_io_enq_bits_vc_sel_0_3),
    .io_deq_ready(vcalloc_q_io_deq_ready),
    .io_deq_valid(vcalloc_q_io_deq_valid),
    .io_deq_bits_vc_sel_2_0(vcalloc_q_io_deq_bits_vc_sel_2_0),
    .io_deq_bits_vc_sel_1_0(vcalloc_q_io_deq_bits_vc_sel_1_0),
    .io_deq_bits_vc_sel_1_1(vcalloc_q_io_deq_bits_vc_sel_1_1),
    .io_deq_bits_vc_sel_1_2(vcalloc_q_io_deq_bits_vc_sel_1_2),
    .io_deq_bits_vc_sel_1_3(vcalloc_q_io_deq_bits_vc_sel_1_3),
    .io_deq_bits_vc_sel_0_0(vcalloc_q_io_deq_bits_vc_sel_0_0),
    .io_deq_bits_vc_sel_0_1(vcalloc_q_io_deq_bits_vc_sel_0_1),
    .io_deq_bits_vc_sel_0_2(vcalloc_q_io_deq_bits_vc_sel_0_2),
    .io_deq_bits_vc_sel_0_3(vcalloc_q_io_deq_bits_vc_sel_0_3)
  );
  assign io_router_req_valid = io_in_valid & route_buffer_io_enq_ready & io_in_bits_head & ~at_dest; // @[IngressUnit.scala 58:86]
  assign io_router_req_bits_flow_ingress_node = route_buffer_io_enq_bits_flow_ingress_node; // @[IngressUnit.scala 53:27]
  assign io_router_req_bits_flow_egress_node = route_buffer_io_enq_bits_flow_egress_node; // @[IngressUnit.scala 53:27]
  assign io_vcalloc_req_valid = _io_vcalloc_req_valid_T_1 & vcalloc_buffer_io_enq_ready & vcalloc_q_io_enq_ready; // @[IngressUnit.scala 92:41]
  assign io_vcalloc_req_bits_vc_sel_2_0 = route_q_io_deq_bits_vc_sel_2_0; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_1_0 = route_q_io_deq_bits_vc_sel_1_0; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_1_1 = route_q_io_deq_bits_vc_sel_1_1; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_1_2 = route_q_io_deq_bits_vc_sel_1_2; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_1_3 = route_q_io_deq_bits_vc_sel_1_3; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_0_0 = route_q_io_deq_bits_vc_sel_0_0; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_0_1 = route_q_io_deq_bits_vc_sel_0_1; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_0_2 = route_q_io_deq_bits_vc_sel_0_2; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_0_3 = route_q_io_deq_bits_vc_sel_0_3; // @[IngressUnit.scala 81:30]
  assign io_salloc_req_0_valid = vcalloc_buffer_io_deq_valid & vcalloc_q_io_deq_valid & c; // @[IngressUnit.scala 109:83]
  assign io_salloc_req_0_bits_vc_sel_2_0 = vcalloc_q_io_deq_bits_vc_sel_2_0; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_1_0 = vcalloc_q_io_deq_bits_vc_sel_1_0; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_1_1 = vcalloc_q_io_deq_bits_vc_sel_1_1; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_1_2 = vcalloc_q_io_deq_bits_vc_sel_1_2; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_1_3 = vcalloc_q_io_deq_bits_vc_sel_1_3; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_0_0 = vcalloc_q_io_deq_bits_vc_sel_0_0; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_0_1 = vcalloc_q_io_deq_bits_vc_sel_0_1; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_0_2 = vcalloc_q_io_deq_bits_vc_sel_0_2; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_0_3 = vcalloc_q_io_deq_bits_vc_sel_0_3; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_tail = vcalloc_buffer_io_deq_bits_tail; // @[IngressUnit.scala 105:30]
  assign io_out_0_valid = out_bundle_valid; // @[IngressUnit.scala 118:13]
  assign io_out_0_bits_flit_head = out_bundle_bits_flit_head; // @[IngressUnit.scala 118:13]
  assign io_out_0_bits_flit_tail = out_bundle_bits_flit_tail; // @[IngressUnit.scala 118:13]
  assign io_out_0_bits_flit_payload = out_bundle_bits_flit_payload; // @[IngressUnit.scala 118:13]
  assign io_out_0_bits_flit_flow_ingress_node = out_bundle_bits_flit_flow_ingress_node; // @[IngressUnit.scala 118:13]
  assign io_out_0_bits_flit_flow_egress_node = out_bundle_bits_flit_flow_egress_node; // @[IngressUnit.scala 118:13]
  assign io_out_0_bits_out_virt_channel = out_bundle_bits_out_virt_channel; // @[IngressUnit.scala 118:13]
  assign io_in_ready = route_buffer_io_enq_ready; // @[IngressUnit.scala 59:44]
  assign route_buffer_clock = clock;
  assign route_buffer_reset = reset;
  assign route_buffer_io_enq_valid = io_in_valid; // @[IngressUnit.scala 56:44]
  assign route_buffer_io_enq_bits_head = io_in_bits_head; // @[IngressUnit.scala 32:33]
  assign route_buffer_io_enq_bits_tail = io_in_bits_tail; // @[IngressUnit.scala 33:33]
  assign route_buffer_io_enq_bits_payload = io_in_bits_payload; // @[IngressUnit.scala 50:36]
  assign route_buffer_io_enq_bits_flow_ingress_node = 2'h0; // @[IngressUnit.scala 38:51]
  assign route_buffer_io_enq_bits_flow_egress_node = _route_buffer_io_enq_bits_flow_egress_node_T_9 |
    _route_buffer_io_enq_bits_flow_egress_node_T_7; // @[Mux.scala 27:73]
  assign route_buffer_io_deq_ready = _route_buffer_io_deq_ready_T_5 & _route_buffer_io_deq_ready_T_7; // @[IngressUnit.scala 95:37]
  assign route_q_clock = clock;
  assign route_q_reset = reset;
  assign route_q_io_enq_valid = _T_13 & io_in_bits_head & at_dest | io_router_req_valid; // @[IngressUnit.scala 62:24 64:53 65:26]
  assign route_q_io_enq_bits_vc_sel_2_0 = _T_13 & io_in_bits_head & at_dest & _T; // @[IngressUnit.scala 63:23 64:53]
  assign route_q_io_enq_bits_vc_sel_1_0 = _T_13 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_1_0; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_1_1 = _T_13 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_1_1; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_1_2 = _T_13 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_1_2; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_1_3 = _T_13 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_1_3; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_0_0 = _T_13 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_0_0; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_0_1 = _T_13 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_0_1; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_0_2 = _T_13 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_0_2; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_0_3 = _T_13 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_0_3; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_deq_ready = _route_q_io_deq_ready_T & route_buffer_io_deq_bits_tail; // @[IngressUnit.scala 97:55]
  assign vcalloc_buffer_clock = clock;
  assign vcalloc_buffer_reset = reset;
  assign vcalloc_buffer_io_enq_valid = _vcalloc_buffer_io_enq_valid_T_2 & _vcalloc_buffer_io_enq_valid_T_4; // @[IngressUnit.scala 88:37]
  assign vcalloc_buffer_io_enq_bits_head = route_buffer_io_deq_bits_head; // @[IngressUnit.scala 79:30]
  assign vcalloc_buffer_io_enq_bits_tail = route_buffer_io_deq_bits_tail; // @[IngressUnit.scala 79:30]
  assign vcalloc_buffer_io_enq_bits_payload = route_buffer_io_deq_bits_payload; // @[IngressUnit.scala 79:30]
  assign vcalloc_buffer_io_enq_bits_flow_ingress_node = route_buffer_io_deq_bits_flow_ingress_node; // @[IngressUnit.scala 79:30]
  assign vcalloc_buffer_io_enq_bits_flow_egress_node = route_buffer_io_deq_bits_flow_egress_node; // @[IngressUnit.scala 79:30]
  assign vcalloc_buffer_io_deq_ready = io_salloc_req_0_ready & vcalloc_q_io_deq_valid & c; // @[IngressUnit.scala 110:83]
  assign vcalloc_q_clock = clock;
  assign vcalloc_q_reset = reset;
  assign vcalloc_q_io_enq_valid = io_vcalloc_req_ready & io_vcalloc_req_valid; // @[Decoupled.scala 51:35]
  assign vcalloc_q_io_enq_bits_vc_sel_2_0 = io_vcalloc_resp_vc_sel_2_0; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_1_0 = io_vcalloc_resp_vc_sel_1_0; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_1_1 = io_vcalloc_resp_vc_sel_1_1; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_1_2 = io_vcalloc_resp_vc_sel_1_2; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_1_3 = io_vcalloc_resp_vc_sel_1_3; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_0_0 = io_vcalloc_resp_vc_sel_0_0; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_0_1 = io_vcalloc_resp_vc_sel_0_1; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_0_2 = io_vcalloc_resp_vc_sel_0_2; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_0_3 = io_vcalloc_resp_vc_sel_0_3; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_deq_ready = vcalloc_buffer_io_deq_bits_tail & _vcalloc_q_io_deq_ready_T; // @[IngressUnit.scala 111:42]
  always @(posedge clock) begin
    out_bundle_valid <= vcalloc_buffer_io_deq_ready & vcalloc_buffer_io_deq_valid; // @[Decoupled.scala 51:35]
    out_bundle_bits_flit_head <= vcalloc_buffer_io_deq_bits_head; // @[IngressUnit.scala 121:24]
    out_bundle_bits_flit_tail <= vcalloc_buffer_io_deq_bits_tail; // @[IngressUnit.scala 121:24]
    out_bundle_bits_flit_payload <= vcalloc_buffer_io_deq_bits_payload; // @[IngressUnit.scala 121:24]
    out_bundle_bits_flit_flow_ingress_node <= vcalloc_buffer_io_deq_bits_flow_ingress_node; // @[IngressUnit.scala 121:24]
    out_bundle_bits_flit_flow_egress_node <= vcalloc_buffer_io_deq_bits_flow_egress_node; // @[IngressUnit.scala 121:24]
    out_bundle_bits_out_virt_channel <= _out_bundle_bits_out_virt_channel_T_10 | _out_bundle_bits_out_virt_channel_T_11; // @[Mux.scala 27:73]
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~(io_in_valid & ~_T_6))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at IngressUnit.scala:30 assert(!(io.in.valid && !cParam.possibleFlows.toSeq.map(_.egressId.U === io.in.bits.egress_id).orR))\n"
            ); // @[IngressUnit.scala 30:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_11 & ~(~(route_q_io_enq_valid & ~route_q_io_enq_ready))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at IngressUnit.scala:73 assert(!(route_q.io.enq.valid && !route_q.io.enq.ready))\n"); // @[IngressUnit.scala 73:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_11 & ~(~(vcalloc_q_io_enq_valid & ~vcalloc_q_io_enq_ready))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at IngressUnit.scala:102 assert(!(vcalloc_q.io.enq.valid && !vcalloc_q.io.enq.ready))\n"
            ); // @[IngressUnit.scala 102:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  out_bundle_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  out_bundle_bits_flit_head = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  out_bundle_bits_flit_tail = _RAND_2[0:0];
  _RAND_3 = {2{`RANDOM}};
  out_bundle_bits_flit_payload = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  out_bundle_bits_flit_flow_ingress_node = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  out_bundle_bits_flit_flow_egress_node = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  out_bundle_bits_out_virt_channel = _RAND_6[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(~(io_in_valid & ~_T_6)); // @[IngressUnit.scala 30:9]
    end
    //
    if (_T_11) begin
      assert(~(route_q_io_enq_valid & ~route_q_io_enq_ready)); // @[IngressUnit.scala 73:9]
    end
    //
    if (_T_11) begin
      assert(~(vcalloc_q_io_enq_valid & ~vcalloc_q_io_enq_ready)); // @[IngressUnit.scala 102:9]
    end
  end
endmodule
module OutputUnit(
  input         clock,
  input         reset,
  input         io_in_0_valid,
  input         io_in_0_bits_head,
  input         io_in_0_bits_tail,
  input  [63:0] io_in_0_bits_payload,
  input  [1:0]  io_in_0_bits_flow_ingress_node,
  input  [1:0]  io_in_0_bits_flow_egress_node,
  input  [1:0]  io_in_0_bits_virt_channel_id,
  output        io_credit_available_0,
  output        io_credit_available_1,
  output        io_credit_available_2,
  output        io_credit_available_3,
  output        io_channel_status_0_occupied,
  output        io_channel_status_1_occupied,
  output        io_channel_status_2_occupied,
  output        io_channel_status_3_occupied,
  input         io_allocs_0_alloc,
  input         io_allocs_1_alloc,
  input         io_allocs_2_alloc,
  input         io_allocs_3_alloc,
  input         io_credit_alloc_0_alloc,
  input         io_credit_alloc_1_alloc,
  input         io_credit_alloc_2_alloc,
  input         io_credit_alloc_3_alloc,
  output        io_out_flit_0_valid,
  output        io_out_flit_0_bits_head,
  output        io_out_flit_0_bits_tail,
  output [63:0] io_out_flit_0_bits_payload,
  output [1:0]  io_out_flit_0_bits_flow_ingress_node,
  output [1:0]  io_out_flit_0_bits_flow_egress_node,
  output [1:0]  io_out_flit_0_bits_virt_channel_id,
  input  [3:0]  io_out_credit_return,
  input  [3:0]  io_out_vc_free
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg  states_3_occupied; // @[OutputUnit.scala 66:19]
  reg [2:0] states_3_c; // @[OutputUnit.scala 66:19]
  reg  states_2_occupied; // @[OutputUnit.scala 66:19]
  reg [2:0] states_2_c; // @[OutputUnit.scala 66:19]
  reg  states_1_occupied; // @[OutputUnit.scala 66:19]
  reg [2:0] states_1_c; // @[OutputUnit.scala 66:19]
  reg  states_0_occupied; // @[OutputUnit.scala 66:19]
  reg [2:0] states_0_c; // @[OutputUnit.scala 66:19]
  wire  _GEN_0 = io_out_vc_free[0] ? 1'h0 : states_0_occupied; // @[OutputUnit.scala 74:30 76:18 66:19]
  wire  _GEN_1 = io_out_vc_free[1] ? 1'h0 : states_1_occupied; // @[OutputUnit.scala 74:30 76:18 66:19]
  wire  _GEN_2 = io_out_vc_free[2] ? 1'h0 : states_2_occupied; // @[OutputUnit.scala 74:30 76:18 66:19]
  wire  _GEN_3 = io_out_vc_free[3] ? 1'h0 : states_3_occupied; // @[OutputUnit.scala 74:30 76:18 66:19]
  wire  _GEN_4 = io_allocs_0_alloc | _GEN_0; // @[OutputUnit.scala 83:20 84:18]
  wire  _GEN_10 = io_allocs_1_alloc | _GEN_1; // @[OutputUnit.scala 83:20 84:18]
  wire  _GEN_16 = io_allocs_2_alloc | _GEN_2; // @[OutputUnit.scala 83:20 84:18]
  wire  _GEN_22 = io_allocs_3_alloc | _GEN_3; // @[OutputUnit.scala 83:20 84:18]
  wire  free = io_out_credit_return[0]; // @[OutputUnit.scala 94:36]
  wire [2:0] _GEN_5 = {{2'd0}, free}; // @[OutputUnit.scala 97:18]
  wire [3:0] _states_0_c_T = states_0_c + _GEN_5; // @[OutputUnit.scala 97:18]
  wire [3:0] _GEN_7 = {{3'd0}, io_credit_alloc_0_alloc}; // @[OutputUnit.scala 97:26]
  wire [3:0] _states_0_c_T_2 = _states_0_c_T - _GEN_7; // @[OutputUnit.scala 97:26]
  wire  free_1 = io_out_credit_return[1]; // @[OutputUnit.scala 94:36]
  wire [2:0] _GEN_9 = {{2'd0}, free_1}; // @[OutputUnit.scala 97:18]
  wire [3:0] _states_1_c_T = states_1_c + _GEN_9; // @[OutputUnit.scala 97:18]
  wire [3:0] _GEN_11 = {{3'd0}, io_credit_alloc_1_alloc}; // @[OutputUnit.scala 97:26]
  wire [3:0] _states_1_c_T_2 = _states_1_c_T - _GEN_11; // @[OutputUnit.scala 97:26]
  wire  free_2 = io_out_credit_return[2]; // @[OutputUnit.scala 94:36]
  wire [2:0] _GEN_13 = {{2'd0}, free_2}; // @[OutputUnit.scala 97:18]
  wire [3:0] _states_2_c_T = states_2_c + _GEN_13; // @[OutputUnit.scala 97:18]
  wire [3:0] _GEN_15 = {{3'd0}, io_credit_alloc_2_alloc}; // @[OutputUnit.scala 97:26]
  wire [3:0] _states_2_c_T_2 = _states_2_c_T - _GEN_15; // @[OutputUnit.scala 97:26]
  wire  free_3 = io_out_credit_return[3]; // @[OutputUnit.scala 94:36]
  wire [2:0] _GEN_17 = {{2'd0}, free_3}; // @[OutputUnit.scala 97:18]
  wire [3:0] _states_3_c_T = states_3_c + _GEN_17; // @[OutputUnit.scala 97:18]
  wire [3:0] _GEN_19 = {{3'd0}, io_credit_alloc_3_alloc}; // @[OutputUnit.scala 97:26]
  wire [3:0] _states_3_c_T_2 = _states_3_c_T - _GEN_19; // @[OutputUnit.scala 97:26]
  wire [3:0] _GEN_32 = reset ? 4'h5 : _states_0_c_T_2; // @[OutputUnit.scala 103:23 105:29 97:11]
  wire [3:0] _GEN_33 = reset ? 4'h5 : _states_1_c_T_2; // @[OutputUnit.scala 103:23 105:29 97:11]
  wire [3:0] _GEN_34 = reset ? 4'h5 : _states_2_c_T_2; // @[OutputUnit.scala 103:23 105:29 97:11]
  wire [3:0] _GEN_35 = reset ? 4'h5 : _states_3_c_T_2; // @[OutputUnit.scala 103:23 105:29 97:11]
  assign io_credit_available_0 = states_0_c != 3'h0; // @[OutputUnit.scala 90:14]
  assign io_credit_available_1 = states_1_c != 3'h0; // @[OutputUnit.scala 90:14]
  assign io_credit_available_2 = states_2_c != 3'h0; // @[OutputUnit.scala 90:14]
  assign io_credit_available_3 = states_3_c != 3'h0; // @[OutputUnit.scala 90:14]
  assign io_channel_status_0_occupied = io_out_vc_free[0] ? 1'h0 : states_0_occupied; // @[OutputUnit.scala 74:30 76:18 66:19]
  assign io_channel_status_1_occupied = io_out_vc_free[1] ? 1'h0 : states_1_occupied; // @[OutputUnit.scala 74:30 76:18 66:19]
  assign io_channel_status_2_occupied = io_out_vc_free[2] ? 1'h0 : states_2_occupied; // @[OutputUnit.scala 74:30 76:18 66:19]
  assign io_channel_status_3_occupied = io_out_vc_free[3] ? 1'h0 : states_3_occupied; // @[OutputUnit.scala 74:30 76:18 66:19]
  assign io_out_flit_0_valid = io_in_0_valid; // @[OutputUnit.scala 71:15]
  assign io_out_flit_0_bits_head = io_in_0_bits_head; // @[OutputUnit.scala 71:15]
  assign io_out_flit_0_bits_tail = io_in_0_bits_tail; // @[OutputUnit.scala 71:15]
  assign io_out_flit_0_bits_payload = io_in_0_bits_payload; // @[OutputUnit.scala 71:15]
  assign io_out_flit_0_bits_flow_ingress_node = io_in_0_bits_flow_ingress_node; // @[OutputUnit.scala 71:15]
  assign io_out_flit_0_bits_flow_egress_node = io_in_0_bits_flow_egress_node; // @[OutputUnit.scala 71:15]
  assign io_out_flit_0_bits_virt_channel_id = io_in_0_bits_virt_channel_id; // @[OutputUnit.scala 71:15]
  always @(posedge clock) begin
    if (reset) begin // @[OutputUnit.scala 103:23]
      states_3_occupied <= 1'h0; // @[OutputUnit.scala 104:31]
    end else begin
      states_3_occupied <= _GEN_22;
    end
    states_3_c <= _GEN_35[2:0];
    if (reset) begin // @[OutputUnit.scala 103:23]
      states_2_occupied <= 1'h0; // @[OutputUnit.scala 104:31]
    end else begin
      states_2_occupied <= _GEN_16;
    end
    states_2_c <= _GEN_34[2:0];
    if (reset) begin // @[OutputUnit.scala 103:23]
      states_1_occupied <= 1'h0; // @[OutputUnit.scala 104:31]
    end else begin
      states_1_occupied <= _GEN_10;
    end
    states_1_c <= _GEN_33[2:0];
    if (reset) begin // @[OutputUnit.scala 103:23]
      states_0_occupied <= 1'h0; // @[OutputUnit.scala 104:31]
    end else begin
      states_0_occupied <= _GEN_4;
    end
    states_0_c <= _GEN_32[2:0];
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_out_vc_free[0] & ~reset & ~states_0_occupied) begin
          $fwrite(32'h80000002,"Assertion failed\n    at OutputUnit.scala:75 assert(s.occupied)\n"); // @[OutputUnit.scala 75:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_out_vc_free[1] & ~reset & ~states_1_occupied) begin
          $fwrite(32'h80000002,"Assertion failed\n    at OutputUnit.scala:75 assert(s.occupied)\n"); // @[OutputUnit.scala 75:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_out_vc_free[2] & ~reset & ~states_2_occupied) begin
          $fwrite(32'h80000002,"Assertion failed\n    at OutputUnit.scala:75 assert(s.occupied)\n"); // @[OutputUnit.scala 75:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_out_vc_free[3] & ~reset & ~states_3_occupied) begin
          $fwrite(32'h80000002,"Assertion failed\n    at OutputUnit.scala:75 assert(s.occupied)\n"); // @[OutputUnit.scala 75:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  states_3_occupied = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  states_3_c = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  states_2_occupied = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  states_2_c = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  states_1_occupied = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  states_1_c = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  states_0_occupied = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  states_0_c = _RAND_7[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (io_out_vc_free[0] & ~reset) begin
      assert(states_0_occupied); // @[OutputUnit.scala 75:13]
    end
    //
    if (io_out_vc_free[1] & ~reset) begin
      assert(states_1_occupied); // @[OutputUnit.scala 75:13]
    end
    //
    if (io_out_vc_free[2] & ~reset) begin
      assert(states_2_occupied); // @[OutputUnit.scala 75:13]
    end
    //
    if (io_out_vc_free[3] & ~reset) begin
      assert(states_3_occupied); // @[OutputUnit.scala 75:13]
    end
  end
endmodule
module Queue_12(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_head,
  input         io_enq_bits_tail,
  input  [63:0] io_enq_bits_payload,
  input  [1:0]  io_enq_bits_ingress_id,
  output        io_deq_valid,
  output        io_deq_bits_head,
  output        io_deq_bits_tail,
  output [63:0] io_deq_bits_payload,
  output [1:0]  io_deq_bits_ingress_id,
  output [1:0]  io_count
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg  ram_head [0:2]; // @[Decoupled.scala 273:95]
  wire  ram_head_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [1:0] ram_head_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_head_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_head_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_tail [0:2]; // @[Decoupled.scala 273:95]
  wire  ram_tail_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [1:0] ram_tail_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_tail_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_tail_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_en; // @[Decoupled.scala 273:95]
  reg [63:0] ram_payload [0:2]; // @[Decoupled.scala 273:95]
  wire  ram_payload_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [1:0] ram_payload_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [63:0] ram_payload_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [63:0] ram_payload_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_payload_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_payload_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_payload_MPORT_en; // @[Decoupled.scala 273:95]
  reg [1:0] ram_ingress_id [0:2]; // @[Decoupled.scala 273:95]
  wire  ram_ingress_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [1:0] ram_ingress_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [1:0] ram_ingress_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_ingress_id_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_ingress_id_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_ingress_id_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_ingress_id_MPORT_en; // @[Decoupled.scala 273:95]
  reg [1:0] enq_ptr_value; // @[Counter.scala 61:40]
  reg [1:0] deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  wrap = enq_ptr_value == 2'h2; // @[Counter.scala 73:24]
  wire [1:0] _value_T_1 = enq_ptr_value + 2'h1; // @[Counter.scala 77:24]
  wire  do_enq = empty ? 1'h0 : _do_enq_T; // @[Decoupled.scala 315:17 280:27]
  wire  wrap_1 = deq_ptr_value == 2'h2; // @[Counter.scala 73:24]
  wire [1:0] _value_T_3 = deq_ptr_value + 2'h1; // @[Counter.scala 77:24]
  wire  do_deq = empty ? 1'h0 : io_deq_valid; // @[Decoupled.scala 315:17 317:14 281:27]
  wire [1:0] ptr_diff = enq_ptr_value - deq_ptr_value; // @[Decoupled.scala 326:32]
  wire [1:0] _io_count_T = maybe_full ? 2'h3 : 2'h0; // @[Decoupled.scala 333:10]
  wire [1:0] _io_count_T_3 = 2'h3 + ptr_diff; // @[Decoupled.scala 334:57]
  wire [1:0] _io_count_T_4 = deq_ptr_value > enq_ptr_value ? _io_count_T_3 : ptr_diff; // @[Decoupled.scala 334:10]
  assign ram_head_io_deq_bits_MPORT_en = 1'h1;
  assign ram_head_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_head_io_deq_bits_MPORT_data = ram_head[ram_head_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  `else
  assign ram_head_io_deq_bits_MPORT_data = ram_head_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_1[0:0] :
    ram_head[ram_head_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_head_MPORT_data = io_enq_bits_head;
  assign ram_head_MPORT_addr = enq_ptr_value;
  assign ram_head_MPORT_mask = 1'h1;
  assign ram_head_MPORT_en = empty ? 1'h0 : _do_enq_T;
  assign ram_tail_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tail_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_tail_io_deq_bits_MPORT_data = ram_tail[ram_tail_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  `else
  assign ram_tail_io_deq_bits_MPORT_data = ram_tail_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_3[0:0] :
    ram_tail[ram_tail_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_tail_MPORT_data = io_enq_bits_tail;
  assign ram_tail_MPORT_addr = enq_ptr_value;
  assign ram_tail_MPORT_mask = 1'h1;
  assign ram_tail_MPORT_en = empty ? 1'h0 : _do_enq_T;
  assign ram_payload_io_deq_bits_MPORT_en = 1'h1;
  assign ram_payload_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_payload_io_deq_bits_MPORT_data = ram_payload[ram_payload_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  `else
  assign ram_payload_io_deq_bits_MPORT_data = ram_payload_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_5[63:0] :
    ram_payload[ram_payload_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_payload_MPORT_data = io_enq_bits_payload;
  assign ram_payload_MPORT_addr = enq_ptr_value;
  assign ram_payload_MPORT_mask = 1'h1;
  assign ram_payload_MPORT_en = empty ? 1'h0 : _do_enq_T;
  assign ram_ingress_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_ingress_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_ingress_id_io_deq_bits_MPORT_data = ram_ingress_id[ram_ingress_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  `else
  assign ram_ingress_id_io_deq_bits_MPORT_data = ram_ingress_id_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_7[1:0] :
    ram_ingress_id[ram_ingress_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_ingress_id_MPORT_data = io_enq_bits_ingress_id;
  assign ram_ingress_id_MPORT_addr = enq_ptr_value;
  assign ram_ingress_id_MPORT_mask = 1'h1;
  assign ram_ingress_id_MPORT_en = empty ? 1'h0 : _do_enq_T;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 302:16 314:{24,39}]
  assign io_deq_bits_head = empty ? io_enq_bits_head : ram_head_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_tail = empty ? io_enq_bits_tail : ram_tail_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_payload = empty ? io_enq_bits_payload : ram_payload_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_ingress_id = empty ? io_enq_bits_ingress_id : ram_ingress_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_count = ptr_match ? _io_count_T : _io_count_T_4; // @[Decoupled.scala 331:20]
  always @(posedge clock) begin
    if (ram_head_MPORT_en & ram_head_MPORT_mask) begin
      ram_head[ram_head_MPORT_addr] <= ram_head_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_tail_MPORT_en & ram_tail_MPORT_mask) begin
      ram_tail[ram_tail_MPORT_addr] <= ram_tail_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_payload_MPORT_en & ram_payload_MPORT_mask) begin
      ram_payload[ram_payload_MPORT_addr] <= ram_payload_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_ingress_id_MPORT_en & ram_ingress_id_MPORT_mask) begin
      ram_ingress_id[ram_ingress_id_MPORT_addr] <= ram_ingress_id_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 2'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      if (wrap) begin // @[Counter.scala 87:20]
        enq_ptr_value <= 2'h0; // @[Counter.scala 87:28]
      end else begin
        enq_ptr_value <= _value_T_1; // @[Counter.scala 77:15]
      end
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 2'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      if (wrap_1) begin // @[Counter.scala 87:20]
        deq_ptr_value <= 2'h0; // @[Counter.scala 87:28]
      end else begin
        deq_ptr_value <= _value_T_3; // @[Counter.scala 77:15]
      end
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      if (empty) begin // @[Decoupled.scala 315:17]
        maybe_full <= 1'h0;
      end else begin
        maybe_full <= _do_enq_T; // @[Decoupled.scala 280:27]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {1{`RANDOM}};
  _RAND_3 = {1{`RANDOM}};
  _RAND_5 = {2{`RANDOM}};
  _RAND_7 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_head[initvar] = _RAND_0[0:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_tail[initvar] = _RAND_2[0:0];
  _RAND_4 = {2{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_payload[initvar] = _RAND_4[63:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_ingress_id[initvar] = _RAND_6[1:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  enq_ptr_value = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  deq_ptr_value = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  maybe_full = _RAND_10[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module EgressUnit(
  input         clock,
  input         reset,
  input         io_in_0_valid,
  input         io_in_0_bits_head,
  input         io_in_0_bits_tail,
  input  [63:0] io_in_0_bits_payload,
  input  [1:0]  io_in_0_bits_flow_ingress_node,
  output        io_credit_available_0,
  output        io_channel_status_0_occupied,
  input         io_allocs_0_alloc,
  input         io_credit_alloc_0_alloc,
  input         io_credit_alloc_0_tail,
  output        io_out_valid,
  output        io_out_bits_head,
  output        io_out_bits_tail,
  output [63:0] io_out_bits_payload,
  output [1:0]  io_out_bits_ingress_id
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  q_clock; // @[EgressUnit.scala 22:17]
  wire  q_reset; // @[EgressUnit.scala 22:17]
  wire  q_io_enq_ready; // @[EgressUnit.scala 22:17]
  wire  q_io_enq_valid; // @[EgressUnit.scala 22:17]
  wire  q_io_enq_bits_head; // @[EgressUnit.scala 22:17]
  wire  q_io_enq_bits_tail; // @[EgressUnit.scala 22:17]
  wire [63:0] q_io_enq_bits_payload; // @[EgressUnit.scala 22:17]
  wire [1:0] q_io_enq_bits_ingress_id; // @[EgressUnit.scala 22:17]
  wire  q_io_deq_valid; // @[EgressUnit.scala 22:17]
  wire  q_io_deq_bits_head; // @[EgressUnit.scala 22:17]
  wire  q_io_deq_bits_tail; // @[EgressUnit.scala 22:17]
  wire [63:0] q_io_deq_bits_payload; // @[EgressUnit.scala 22:17]
  wire [1:0] q_io_deq_bits_ingress_id; // @[EgressUnit.scala 22:17]
  wire [1:0] q_io_count; // @[EgressUnit.scala 22:17]
  reg  channel_empty; // @[EgressUnit.scala 20:30]
  wire  _q_io_enq_bits_ingress_id_T_3 = 2'h1 == io_in_0_bits_flow_ingress_node; // @[EgressUnit.scala 31:39]
  wire  _q_io_enq_bits_ingress_id_T_6 = 2'h2 == io_in_0_bits_flow_ingress_node; // @[EgressUnit.scala 31:39]
  wire  _q_io_enq_bits_ingress_id_T_9 = 2'h3 == io_in_0_bits_flow_ingress_node; // @[EgressUnit.scala 31:39]
  wire [1:0] _q_io_enq_bits_ingress_id_T_13 = _q_io_enq_bits_ingress_id_T_3 ? 2'h1 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _q_io_enq_bits_ingress_id_T_14 = _q_io_enq_bits_ingress_id_T_6 ? 2'h2 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _q_io_enq_bits_ingress_id_T_15 = _q_io_enq_bits_ingress_id_T_9 ? 2'h3 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _q_io_enq_bits_ingress_id_T_17 = _q_io_enq_bits_ingress_id_T_13 | _q_io_enq_bits_ingress_id_T_14; // @[Mux.scala 27:73]
  wire  _GEN_0 = io_credit_alloc_0_alloc & io_credit_alloc_0_tail | channel_empty; // @[EgressUnit.scala 44:62 45:19 20:30]
  wire  _GEN_1 = io_allocs_0_alloc ? 1'h0 : _GEN_0; // @[EgressUnit.scala 49:29 50:19]
  Queue_12 q ( // @[EgressUnit.scala 22:17]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_head(q_io_enq_bits_head),
    .io_enq_bits_tail(q_io_enq_bits_tail),
    .io_enq_bits_payload(q_io_enq_bits_payload),
    .io_enq_bits_ingress_id(q_io_enq_bits_ingress_id),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_head(q_io_deq_bits_head),
    .io_deq_bits_tail(q_io_deq_bits_tail),
    .io_deq_bits_payload(q_io_deq_bits_payload),
    .io_deq_bits_ingress_id(q_io_deq_bits_ingress_id),
    .io_count(q_io_count)
  );
  assign io_credit_available_0 = q_io_count == 2'h0; // @[EgressUnit.scala 40:40]
  assign io_channel_status_0_occupied = ~channel_empty; // @[EgressUnit.scala 41:36]
  assign io_out_valid = q_io_deq_valid; // @[EgressUnit.scala 37:10]
  assign io_out_bits_head = q_io_deq_bits_head; // @[EgressUnit.scala 37:10]
  assign io_out_bits_tail = q_io_deq_bits_tail; // @[EgressUnit.scala 37:10]
  assign io_out_bits_payload = q_io_deq_bits_payload; // @[EgressUnit.scala 37:10]
  assign io_out_bits_ingress_id = q_io_deq_bits_ingress_id; // @[EgressUnit.scala 37:10]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_in_0_valid; // @[EgressUnit.scala 23:18]
  assign q_io_enq_bits_head = io_in_0_bits_head; // @[EgressUnit.scala 24:22]
  assign q_io_enq_bits_tail = io_in_0_bits_tail; // @[EgressUnit.scala 25:22]
  assign q_io_enq_bits_payload = io_in_0_bits_payload; // @[EgressUnit.scala 36:25]
  assign q_io_enq_bits_ingress_id = _q_io_enq_bits_ingress_id_T_17 | _q_io_enq_bits_ingress_id_T_15; // @[Mux.scala 27:73]
  always @(posedge clock) begin
    channel_empty <= reset | _GEN_1; // @[EgressUnit.scala 20:{30,30}]
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~(q_io_enq_valid & ~q_io_enq_ready))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at EgressUnit.scala:38 assert(!(q.io.enq.valid && !q.io.enq.ready))\n"); // @[EgressUnit.scala 38:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  channel_empty = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(~(q_io_enq_valid & ~q_io_enq_ready)); // @[EgressUnit.scala 38:9]
    end
  end
endmodule
module Switch(
  input         clock,
  input         reset,
  input         io_in_2_0_valid,
  input         io_in_2_0_bits_flit_head,
  input         io_in_2_0_bits_flit_tail,
  input  [63:0] io_in_2_0_bits_flit_payload,
  input  [1:0]  io_in_2_0_bits_flit_flow_ingress_node,
  input  [1:0]  io_in_2_0_bits_flit_flow_egress_node,
  input  [1:0]  io_in_2_0_bits_out_virt_channel,
  input         io_in_1_0_valid,
  input         io_in_1_0_bits_flit_head,
  input         io_in_1_0_bits_flit_tail,
  input  [63:0] io_in_1_0_bits_flit_payload,
  input  [1:0]  io_in_1_0_bits_flit_flow_ingress_node,
  input  [1:0]  io_in_1_0_bits_flit_flow_egress_node,
  input  [1:0]  io_in_1_0_bits_out_virt_channel,
  input         io_in_0_0_valid,
  input         io_in_0_0_bits_flit_head,
  input         io_in_0_0_bits_flit_tail,
  input  [63:0] io_in_0_0_bits_flit_payload,
  input  [1:0]  io_in_0_0_bits_flit_flow_ingress_node,
  input  [1:0]  io_in_0_0_bits_flit_flow_egress_node,
  input  [1:0]  io_in_0_0_bits_out_virt_channel,
  output        io_out_2_0_valid,
  output        io_out_2_0_bits_head,
  output        io_out_2_0_bits_tail,
  output [63:0] io_out_2_0_bits_payload,
  output [1:0]  io_out_2_0_bits_flow_ingress_node,
  output        io_out_1_0_valid,
  output        io_out_1_0_bits_head,
  output        io_out_1_0_bits_tail,
  output [63:0] io_out_1_0_bits_payload,
  output [1:0]  io_out_1_0_bits_flow_ingress_node,
  output [1:0]  io_out_1_0_bits_flow_egress_node,
  output [1:0]  io_out_1_0_bits_virt_channel_id,
  output        io_out_0_0_valid,
  output        io_out_0_0_bits_head,
  output        io_out_0_0_bits_tail,
  output [63:0] io_out_0_0_bits_payload,
  output [1:0]  io_out_0_0_bits_flow_ingress_node,
  output [1:0]  io_out_0_0_bits_flow_egress_node,
  output [1:0]  io_out_0_0_bits_virt_channel_id,
  input         io_sel_2_0_2_0,
  input         io_sel_2_0_1_0,
  input         io_sel_2_0_0_0,
  input         io_sel_1_0_2_0,
  input         io_sel_1_0_1_0,
  input         io_sel_1_0_0_0,
  input         io_sel_0_0_2_0,
  input         io_sel_0_0_1_0,
  input         io_sel_0_0_0_0
);
  wire [2:0] sel_flat = {io_sel_0_0_2_0,io_sel_0_0_1_0,io_sel_0_0_0_0}; // @[Switch.scala 46:35]
  wire [1:0] _T_3 = sel_flat[1] + sel_flat[2]; // @[Bitwise.scala 51:90]
  wire [1:0] _GEN_0 = {{1'd0}, sel_flat[0]}; // @[Bitwise.scala 51:90]
  wire [2:0] _T_5 = _GEN_0 + _T_3; // @[Bitwise.scala 51:90]
  wire  _io_out_0_0_valid_T_7 = sel_flat[0] & io_in_0_0_valid | sel_flat[1] & io_in_1_0_valid | sel_flat[2] &
    io_in_2_0_valid; // @[Mux.scala 27:73]
  wire [1:0] _io_out_0_0_bits_T_13 = sel_flat[0] ? io_in_0_0_bits_flit_flow_egress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_0_0_bits_T_14 = sel_flat[1] ? io_in_1_0_bits_flit_flow_egress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_0_0_bits_T_15 = sel_flat[2] ? io_in_2_0_bits_flit_flow_egress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_0_0_bits_T_16 = _io_out_0_0_bits_T_13 | _io_out_0_0_bits_T_14; // @[Mux.scala 27:73]
  wire [1:0] _io_out_0_0_bits_T_23 = sel_flat[0] ? io_in_0_0_bits_flit_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_0_0_bits_T_24 = sel_flat[1] ? io_in_1_0_bits_flit_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_0_0_bits_T_25 = sel_flat[2] ? io_in_2_0_bits_flit_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_0_0_bits_T_26 = _io_out_0_0_bits_T_23 | _io_out_0_0_bits_T_24; // @[Mux.scala 27:73]
  wire [63:0] _io_out_0_0_bits_T_33 = sel_flat[0] ? io_in_0_0_bits_flit_payload : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_out_0_0_bits_T_34 = sel_flat[1] ? io_in_1_0_bits_flit_payload : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_out_0_0_bits_T_35 = sel_flat[2] ? io_in_2_0_bits_flit_payload : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_out_0_0_bits_T_36 = _io_out_0_0_bits_T_33 | _io_out_0_0_bits_T_34; // @[Mux.scala 27:73]
  wire [1:0] _io_out_0_0_bits_virt_channel_id_T_3 = sel_flat[0] ? io_in_0_0_bits_out_virt_channel : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_0_0_bits_virt_channel_id_T_4 = sel_flat[1] ? io_in_1_0_bits_out_virt_channel : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_0_0_bits_virt_channel_id_T_5 = sel_flat[2] ? io_in_2_0_bits_out_virt_channel : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_0_0_bits_virt_channel_id_T_6 = _io_out_0_0_bits_virt_channel_id_T_3 |
    _io_out_0_0_bits_virt_channel_id_T_4; // @[Mux.scala 27:73]
  wire [2:0] sel_flat_1 = {io_sel_1_0_2_0,io_sel_1_0_1_0,io_sel_1_0_0_0}; // @[Switch.scala 46:35]
  wire [1:0] _T_14 = sel_flat_1[1] + sel_flat_1[2]; // @[Bitwise.scala 51:90]
  wire [1:0] _GEN_1 = {{1'd0}, sel_flat_1[0]}; // @[Bitwise.scala 51:90]
  wire [2:0] _T_16 = _GEN_1 + _T_14; // @[Bitwise.scala 51:90]
  wire  _io_out_1_0_valid_T_7 = sel_flat_1[0] & io_in_0_0_valid | sel_flat_1[1] & io_in_1_0_valid | sel_flat_1[2] &
    io_in_2_0_valid; // @[Mux.scala 27:73]
  wire [1:0] _io_out_1_0_bits_T_13 = sel_flat_1[0] ? io_in_0_0_bits_flit_flow_egress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_1_0_bits_T_14 = sel_flat_1[1] ? io_in_1_0_bits_flit_flow_egress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_1_0_bits_T_15 = sel_flat_1[2] ? io_in_2_0_bits_flit_flow_egress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_1_0_bits_T_16 = _io_out_1_0_bits_T_13 | _io_out_1_0_bits_T_14; // @[Mux.scala 27:73]
  wire [1:0] _io_out_1_0_bits_T_23 = sel_flat_1[0] ? io_in_0_0_bits_flit_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_1_0_bits_T_24 = sel_flat_1[1] ? io_in_1_0_bits_flit_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_1_0_bits_T_25 = sel_flat_1[2] ? io_in_2_0_bits_flit_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_1_0_bits_T_26 = _io_out_1_0_bits_T_23 | _io_out_1_0_bits_T_24; // @[Mux.scala 27:73]
  wire [63:0] _io_out_1_0_bits_T_33 = sel_flat_1[0] ? io_in_0_0_bits_flit_payload : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_out_1_0_bits_T_34 = sel_flat_1[1] ? io_in_1_0_bits_flit_payload : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_out_1_0_bits_T_35 = sel_flat_1[2] ? io_in_2_0_bits_flit_payload : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_out_1_0_bits_T_36 = _io_out_1_0_bits_T_33 | _io_out_1_0_bits_T_34; // @[Mux.scala 27:73]
  wire [1:0] _io_out_1_0_bits_virt_channel_id_T_3 = sel_flat_1[0] ? io_in_0_0_bits_out_virt_channel : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_1_0_bits_virt_channel_id_T_4 = sel_flat_1[1] ? io_in_1_0_bits_out_virt_channel : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_1_0_bits_virt_channel_id_T_5 = sel_flat_1[2] ? io_in_2_0_bits_out_virt_channel : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_1_0_bits_virt_channel_id_T_6 = _io_out_1_0_bits_virt_channel_id_T_3 |
    _io_out_1_0_bits_virt_channel_id_T_4; // @[Mux.scala 27:73]
  wire [2:0] sel_flat_2 = {io_sel_2_0_2_0,io_sel_2_0_1_0,io_sel_2_0_0_0}; // @[Switch.scala 46:35]
  wire [1:0] _T_25 = sel_flat_2[1] + sel_flat_2[2]; // @[Bitwise.scala 51:90]
  wire [1:0] _GEN_2 = {{1'd0}, sel_flat_2[0]}; // @[Bitwise.scala 51:90]
  wire [2:0] _T_27 = _GEN_2 + _T_25; // @[Bitwise.scala 51:90]
  wire  _io_out_2_0_valid_T_7 = sel_flat_2[0] & io_in_0_0_valid | sel_flat_2[1] & io_in_1_0_valid | sel_flat_2[2] &
    io_in_2_0_valid; // @[Mux.scala 27:73]
  wire [1:0] _io_out_2_0_bits_T_23 = sel_flat_2[0] ? io_in_0_0_bits_flit_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_2_0_bits_T_24 = sel_flat_2[1] ? io_in_1_0_bits_flit_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_2_0_bits_T_25 = sel_flat_2[2] ? io_in_2_0_bits_flit_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_2_0_bits_T_26 = _io_out_2_0_bits_T_23 | _io_out_2_0_bits_T_24; // @[Mux.scala 27:73]
  wire [63:0] _io_out_2_0_bits_T_33 = sel_flat_2[0] ? io_in_0_0_bits_flit_payload : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_out_2_0_bits_T_34 = sel_flat_2[1] ? io_in_1_0_bits_flit_payload : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_out_2_0_bits_T_35 = sel_flat_2[2] ? io_in_2_0_bits_flit_payload : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_out_2_0_bits_T_36 = _io_out_2_0_bits_T_33 | _io_out_2_0_bits_T_34; // @[Mux.scala 27:73]
  assign io_out_2_0_valid = _io_out_2_0_valid_T_7 & sel_flat_2 != 3'h0; // @[Switch.scala 48:67]
  assign io_out_2_0_bits_head = sel_flat_2[0] & io_in_0_0_bits_flit_head | sel_flat_2[1] & io_in_1_0_bits_flit_head |
    sel_flat_2[2] & io_in_2_0_bits_flit_head; // @[Mux.scala 27:73]
  assign io_out_2_0_bits_tail = sel_flat_2[0] & io_in_0_0_bits_flit_tail | sel_flat_2[1] & io_in_1_0_bits_flit_tail |
    sel_flat_2[2] & io_in_2_0_bits_flit_tail; // @[Mux.scala 27:73]
  assign io_out_2_0_bits_payload = _io_out_2_0_bits_T_36 | _io_out_2_0_bits_T_35; // @[Mux.scala 27:73]
  assign io_out_2_0_bits_flow_ingress_node = _io_out_2_0_bits_T_26 | _io_out_2_0_bits_T_25; // @[Mux.scala 27:73]
  assign io_out_1_0_valid = _io_out_1_0_valid_T_7 & sel_flat_1 != 3'h0; // @[Switch.scala 48:67]
  assign io_out_1_0_bits_head = sel_flat_1[0] & io_in_0_0_bits_flit_head | sel_flat_1[1] & io_in_1_0_bits_flit_head |
    sel_flat_1[2] & io_in_2_0_bits_flit_head; // @[Mux.scala 27:73]
  assign io_out_1_0_bits_tail = sel_flat_1[0] & io_in_0_0_bits_flit_tail | sel_flat_1[1] & io_in_1_0_bits_flit_tail |
    sel_flat_1[2] & io_in_2_0_bits_flit_tail; // @[Mux.scala 27:73]
  assign io_out_1_0_bits_payload = _io_out_1_0_bits_T_36 | _io_out_1_0_bits_T_35; // @[Mux.scala 27:73]
  assign io_out_1_0_bits_flow_ingress_node = _io_out_1_0_bits_T_26 | _io_out_1_0_bits_T_25; // @[Mux.scala 27:73]
  assign io_out_1_0_bits_flow_egress_node = _io_out_1_0_bits_T_16 | _io_out_1_0_bits_T_15; // @[Mux.scala 27:73]
  assign io_out_1_0_bits_virt_channel_id = _io_out_1_0_bits_virt_channel_id_T_6 | _io_out_1_0_bits_virt_channel_id_T_5; // @[Mux.scala 27:73]
  assign io_out_0_0_valid = _io_out_0_0_valid_T_7 & sel_flat != 3'h0; // @[Switch.scala 48:67]
  assign io_out_0_0_bits_head = sel_flat[0] & io_in_0_0_bits_flit_head | sel_flat[1] & io_in_1_0_bits_flit_head |
    sel_flat[2] & io_in_2_0_bits_flit_head; // @[Mux.scala 27:73]
  assign io_out_0_0_bits_tail = sel_flat[0] & io_in_0_0_bits_flit_tail | sel_flat[1] & io_in_1_0_bits_flit_tail |
    sel_flat[2] & io_in_2_0_bits_flit_tail; // @[Mux.scala 27:73]
  assign io_out_0_0_bits_payload = _io_out_0_0_bits_T_36 | _io_out_0_0_bits_T_35; // @[Mux.scala 27:73]
  assign io_out_0_0_bits_flow_ingress_node = _io_out_0_0_bits_T_26 | _io_out_0_0_bits_T_25; // @[Mux.scala 27:73]
  assign io_out_0_0_bits_flow_egress_node = _io_out_0_0_bits_T_16 | _io_out_0_0_bits_T_15; // @[Mux.scala 27:73]
  assign io_out_0_0_bits_virt_channel_id = _io_out_0_0_bits_virt_channel_id_T_6 | _io_out_0_0_bits_virt_channel_id_T_5; // @[Mux.scala 27:73]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(_T_5[1:0] <= 2'h1)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Switch.scala:47 assert(PopCount(sel_flat) <= 1.U)\n"); // @[Switch.scala 47:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(_T_16[1:0] <= 2'h1)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Switch.scala:47 assert(PopCount(sel_flat) <= 1.U)\n"); // @[Switch.scala 47:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(_T_27[1:0] <= 2'h1)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Switch.scala:47 assert(PopCount(sel_flat) <= 1.U)\n"); // @[Switch.scala 47:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(_T_5[1:0] <= 2'h1); // @[Switch.scala 47:13]
    end
    //
    if (~reset) begin
      assert(_T_16[1:0] <= 2'h1); // @[Switch.scala 47:13]
    end
    //
    if (~reset) begin
      assert(_T_27[1:0] <= 2'h1); // @[Switch.scala 47:13]
    end
  end
endmodule
module SwitchArbiter_2(
  input        clock,
  input        reset,
  output       io_in_0_ready,
  input        io_in_0_valid,
  input        io_in_0_bits_vc_sel_2_0,
  input        io_in_0_bits_vc_sel_1_0,
  input        io_in_0_bits_vc_sel_1_1,
  input        io_in_0_bits_vc_sel_1_2,
  input        io_in_0_bits_vc_sel_1_3,
  input        io_in_0_bits_vc_sel_0_0,
  input        io_in_0_bits_vc_sel_0_1,
  input        io_in_0_bits_vc_sel_0_2,
  input        io_in_0_bits_vc_sel_0_3,
  input        io_in_0_bits_tail,
  output       io_in_1_ready,
  input        io_in_1_valid,
  input        io_in_1_bits_vc_sel_2_0,
  input        io_in_1_bits_vc_sel_1_0,
  input        io_in_1_bits_vc_sel_1_1,
  input        io_in_1_bits_vc_sel_1_2,
  input        io_in_1_bits_vc_sel_1_3,
  input        io_in_1_bits_vc_sel_0_0,
  input        io_in_1_bits_vc_sel_0_1,
  input        io_in_1_bits_vc_sel_0_2,
  input        io_in_1_bits_vc_sel_0_3,
  input        io_in_1_bits_tail,
  output       io_in_2_ready,
  input        io_in_2_valid,
  input        io_in_2_bits_vc_sel_2_0,
  input        io_in_2_bits_vc_sel_1_0,
  input        io_in_2_bits_vc_sel_1_1,
  input        io_in_2_bits_vc_sel_1_2,
  input        io_in_2_bits_vc_sel_1_3,
  input        io_in_2_bits_vc_sel_0_0,
  input        io_in_2_bits_vc_sel_0_1,
  input        io_in_2_bits_vc_sel_0_2,
  input        io_in_2_bits_vc_sel_0_3,
  input        io_in_2_bits_tail,
  output       io_out_0_valid,
  output       io_out_0_bits_vc_sel_2_0,
  output       io_out_0_bits_vc_sel_1_0,
  output       io_out_0_bits_vc_sel_1_1,
  output       io_out_0_bits_vc_sel_1_2,
  output       io_out_0_bits_vc_sel_1_3,
  output       io_out_0_bits_vc_sel_0_0,
  output       io_out_0_bits_vc_sel_0_1,
  output       io_out_0_bits_vc_sel_0_2,
  output       io_out_0_bits_vc_sel_0_3,
  output       io_out_0_bits_tail,
  output [2:0] io_chosen_oh_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] lock_0; // @[SwitchAllocator.scala 24:38]
  wire [2:0] _unassigned_T = {io_in_2_valid,io_in_1_valid,io_in_0_valid}; // @[Cat.scala 33:92]
  wire [2:0] _unassigned_T_1 = ~lock_0; // @[SwitchAllocator.scala 25:54]
  wire [2:0] unassigned = _unassigned_T & _unassigned_T_1; // @[SwitchAllocator.scala 25:52]
  reg [2:0] mask; // @[SwitchAllocator.scala 27:21]
  wire [2:0] _GEN_5 = {{2'd0}, mask == 3'h0}; // @[SwitchAllocator.scala 30:58]
  wire [2:0] _sel_T_1 = unassigned & _GEN_5; // @[SwitchAllocator.scala 30:58]
  wire [5:0] _sel_T_2 = {unassigned,_sel_T_1}; // @[Cat.scala 33:92]
  wire [5:0] _sel_T_9 = _sel_T_2[5] ? 6'h20 : 6'h0; // @[Mux.scala 47:70]
  wire [5:0] _sel_T_10 = _sel_T_2[4] ? 6'h10 : _sel_T_9; // @[Mux.scala 47:70]
  wire [5:0] _sel_T_11 = _sel_T_2[3] ? 6'h8 : _sel_T_10; // @[Mux.scala 47:70]
  wire [5:0] _sel_T_12 = _sel_T_2[2] ? 6'h4 : _sel_T_11; // @[Mux.scala 47:70]
  wire [5:0] _sel_T_13 = _sel_T_2[1] ? 6'h2 : _sel_T_12; // @[Mux.scala 47:70]
  wire [5:0] sel = _sel_T_2[0] ? 6'h1 : _sel_T_13; // @[Mux.scala 47:70]
  wire [5:0] _GEN_6 = {{3'd0}, sel[5:3]}; // @[SwitchAllocator.scala 32:23]
  wire [5:0] _choices_0_T_1 = sel | _GEN_6; // @[SwitchAllocator.scala 32:23]
  wire [2:0] choices_0 = _choices_0_T_1[2:0]; // @[SwitchAllocator.scala 28:21 32:16]
  wire [2:0] in_tails = {io_in_2_bits_tail,io_in_1_bits_tail,io_in_0_bits_tail}; // @[Cat.scala 33:92]
  wire [2:0] _chosen_T = _unassigned_T & lock_0; // @[SwitchAllocator.scala 42:33]
  wire [2:0] chosen = |_chosen_T ? lock_0 : choices_0; // @[SwitchAllocator.scala 42:21]
  wire [2:0] _io_out_0_valid_T = _unassigned_T & chosen; // @[SwitchAllocator.scala 44:35]
  wire [2:0] _lock_0_T = ~in_tails; // @[SwitchAllocator.scala 53:27]
  wire [2:0] _lock_0_T_1 = chosen & _lock_0_T; // @[SwitchAllocator.scala 53:25]
  wire [2:0] _GEN_7 = {{1'd0}, io_chosen_oh_0[2:1]}; // @[SwitchAllocator.scala 58:71]
  wire [2:0] _mask_T_3 = io_chosen_oh_0 | _GEN_7; // @[SwitchAllocator.scala 58:71]
  wire [2:0] _GEN_8 = {{2'd0}, io_chosen_oh_0[2]}; // @[SwitchAllocator.scala 58:71]
  wire [2:0] _mask_T_4 = _mask_T_3 | _GEN_8; // @[SwitchAllocator.scala 58:71]
  wire [2:0] _mask_T_5 = ~mask; // @[SwitchAllocator.scala 60:17]
  wire [3:0] _mask_T_7 = {mask, 1'h0}; // @[SwitchAllocator.scala 60:43]
  wire [3:0] _mask_T_8 = _mask_T_7 | 4'h1; // @[SwitchAllocator.scala 60:49]
  wire [3:0] _mask_T_9 = _mask_T_5 == 3'h0 ? 4'h0 : _mask_T_8; // @[SwitchAllocator.scala 60:16]
  wire [3:0] _GEN_4 = io_out_0_valid ? {{1'd0}, _mask_T_4} : _mask_T_9; // @[SwitchAllocator.scala 57:27 58:10 60:10]
  wire [3:0] _GEN_9 = reset ? 4'h0 : _GEN_4; // @[SwitchAllocator.scala 27:{21,21}]
  assign io_in_0_ready = chosen[0]; // @[SwitchAllocator.scala 47:19]
  assign io_in_1_ready = chosen[1]; // @[SwitchAllocator.scala 47:19]
  assign io_in_2_ready = chosen[2]; // @[SwitchAllocator.scala 47:19]
  assign io_out_0_valid = |_io_out_0_valid_T; // @[SwitchAllocator.scala 44:45]
  assign io_out_0_bits_vc_sel_2_0 = chosen[0] & io_in_0_bits_vc_sel_2_0 | chosen[1] & io_in_1_bits_vc_sel_2_0 | chosen[2
    ] & io_in_2_bits_vc_sel_2_0; // @[Mux.scala 27:73]
  assign io_out_0_bits_vc_sel_1_0 = chosen[0] & io_in_0_bits_vc_sel_1_0 | chosen[1] & io_in_1_bits_vc_sel_1_0 | chosen[2
    ] & io_in_2_bits_vc_sel_1_0; // @[Mux.scala 27:73]
  assign io_out_0_bits_vc_sel_1_1 = chosen[0] & io_in_0_bits_vc_sel_1_1 | chosen[1] & io_in_1_bits_vc_sel_1_1 | chosen[2
    ] & io_in_2_bits_vc_sel_1_1; // @[Mux.scala 27:73]
  assign io_out_0_bits_vc_sel_1_2 = chosen[0] & io_in_0_bits_vc_sel_1_2 | chosen[1] & io_in_1_bits_vc_sel_1_2 | chosen[2
    ] & io_in_2_bits_vc_sel_1_2; // @[Mux.scala 27:73]
  assign io_out_0_bits_vc_sel_1_3 = chosen[0] & io_in_0_bits_vc_sel_1_3 | chosen[1] & io_in_1_bits_vc_sel_1_3 | chosen[2
    ] & io_in_2_bits_vc_sel_1_3; // @[Mux.scala 27:73]
  assign io_out_0_bits_vc_sel_0_0 = chosen[0] & io_in_0_bits_vc_sel_0_0 | chosen[1] & io_in_1_bits_vc_sel_0_0 | chosen[2
    ] & io_in_2_bits_vc_sel_0_0; // @[Mux.scala 27:73]
  assign io_out_0_bits_vc_sel_0_1 = chosen[0] & io_in_0_bits_vc_sel_0_1 | chosen[1] & io_in_1_bits_vc_sel_0_1 | chosen[2
    ] & io_in_2_bits_vc_sel_0_1; // @[Mux.scala 27:73]
  assign io_out_0_bits_vc_sel_0_2 = chosen[0] & io_in_0_bits_vc_sel_0_2 | chosen[1] & io_in_1_bits_vc_sel_0_2 | chosen[2
    ] & io_in_2_bits_vc_sel_0_2; // @[Mux.scala 27:73]
  assign io_out_0_bits_vc_sel_0_3 = chosen[0] & io_in_0_bits_vc_sel_0_3 | chosen[1] & io_in_1_bits_vc_sel_0_3 | chosen[2
    ] & io_in_2_bits_vc_sel_0_3; // @[Mux.scala 27:73]
  assign io_out_0_bits_tail = chosen[0] & io_in_0_bits_tail | chosen[1] & io_in_1_bits_tail | chosen[2] &
    io_in_2_bits_tail; // @[Mux.scala 27:73]
  assign io_chosen_oh_0 = |_chosen_T ? lock_0 : choices_0; // @[SwitchAllocator.scala 42:21]
  always @(posedge clock) begin
    if (reset) begin // @[SwitchAllocator.scala 24:38]
      lock_0 <= 3'h0; // @[SwitchAllocator.scala 24:38]
    end else if (io_out_0_valid) begin // @[SwitchAllocator.scala 52:29]
      lock_0 <= _lock_0_T_1; // @[SwitchAllocator.scala 53:15]
    end
    mask <= _GEN_9[2:0]; // @[SwitchAllocator.scala 27:{21,21}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lock_0 = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  mask = _RAND_1[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SwitchAllocator(
  input   clock,
  input   reset,
  output  io_req_2_0_ready,
  input   io_req_2_0_valid,
  input   io_req_2_0_bits_vc_sel_2_0,
  input   io_req_2_0_bits_vc_sel_1_0,
  input   io_req_2_0_bits_vc_sel_1_1,
  input   io_req_2_0_bits_vc_sel_1_2,
  input   io_req_2_0_bits_vc_sel_1_3,
  input   io_req_2_0_bits_vc_sel_0_0,
  input   io_req_2_0_bits_vc_sel_0_1,
  input   io_req_2_0_bits_vc_sel_0_2,
  input   io_req_2_0_bits_vc_sel_0_3,
  input   io_req_2_0_bits_tail,
  output  io_req_1_0_ready,
  input   io_req_1_0_valid,
  input   io_req_1_0_bits_vc_sel_2_0,
  input   io_req_1_0_bits_vc_sel_1_0,
  input   io_req_1_0_bits_vc_sel_1_1,
  input   io_req_1_0_bits_vc_sel_1_2,
  input   io_req_1_0_bits_vc_sel_1_3,
  input   io_req_1_0_bits_vc_sel_0_0,
  input   io_req_1_0_bits_vc_sel_0_1,
  input   io_req_1_0_bits_vc_sel_0_2,
  input   io_req_1_0_bits_vc_sel_0_3,
  input   io_req_1_0_bits_tail,
  output  io_req_0_0_ready,
  input   io_req_0_0_valid,
  input   io_req_0_0_bits_vc_sel_2_0,
  input   io_req_0_0_bits_vc_sel_1_0,
  input   io_req_0_0_bits_vc_sel_1_1,
  input   io_req_0_0_bits_vc_sel_1_2,
  input   io_req_0_0_bits_vc_sel_1_3,
  input   io_req_0_0_bits_vc_sel_0_0,
  input   io_req_0_0_bits_vc_sel_0_1,
  input   io_req_0_0_bits_vc_sel_0_2,
  input   io_req_0_0_bits_vc_sel_0_3,
  input   io_req_0_0_bits_tail,
  output  io_credit_alloc_2_0_alloc,
  output  io_credit_alloc_2_0_tail,
  output  io_credit_alloc_1_0_alloc,
  output  io_credit_alloc_1_1_alloc,
  output  io_credit_alloc_1_2_alloc,
  output  io_credit_alloc_1_3_alloc,
  output  io_credit_alloc_0_0_alloc,
  output  io_credit_alloc_0_1_alloc,
  output  io_credit_alloc_0_2_alloc,
  output  io_credit_alloc_0_3_alloc,
  output  io_switch_sel_2_0_2_0,
  output  io_switch_sel_2_0_1_0,
  output  io_switch_sel_2_0_0_0,
  output  io_switch_sel_1_0_2_0,
  output  io_switch_sel_1_0_1_0,
  output  io_switch_sel_1_0_0_0,
  output  io_switch_sel_0_0_2_0,
  output  io_switch_sel_0_0_1_0,
  output  io_switch_sel_0_0_0_0
);
  wire  arbs_0_clock; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_reset; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_0_ready; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_0_valid; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_0_bits_vc_sel_2_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_0_bits_vc_sel_1_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_0_bits_vc_sel_1_1; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_0_bits_vc_sel_1_2; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_0_bits_vc_sel_1_3; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_0_bits_vc_sel_0_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_0_bits_vc_sel_0_1; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_0_bits_vc_sel_0_2; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_0_bits_vc_sel_0_3; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_0_bits_tail; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_1_ready; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_1_valid; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_1_bits_vc_sel_2_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_1_bits_vc_sel_1_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_1_bits_vc_sel_1_1; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_1_bits_vc_sel_1_2; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_1_bits_vc_sel_1_3; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_1_bits_vc_sel_0_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_1_bits_vc_sel_0_1; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_1_bits_vc_sel_0_2; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_1_bits_vc_sel_0_3; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_1_bits_tail; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_2_ready; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_2_valid; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_2_bits_vc_sel_2_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_2_bits_vc_sel_1_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_2_bits_vc_sel_1_1; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_2_bits_vc_sel_1_2; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_2_bits_vc_sel_1_3; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_2_bits_vc_sel_0_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_2_bits_vc_sel_0_1; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_2_bits_vc_sel_0_2; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_2_bits_vc_sel_0_3; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_2_bits_tail; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_out_0_valid; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_out_0_bits_vc_sel_2_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_out_0_bits_vc_sel_1_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_out_0_bits_vc_sel_1_1; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_out_0_bits_vc_sel_1_2; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_out_0_bits_vc_sel_1_3; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_out_0_bits_vc_sel_0_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_out_0_bits_vc_sel_0_1; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_out_0_bits_vc_sel_0_2; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_out_0_bits_vc_sel_0_3; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_out_0_bits_tail; // @[SwitchAllocator.scala 83:45]
  wire [2:0] arbs_0_io_chosen_oh_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_clock; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_reset; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_0_ready; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_0_valid; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_0_bits_vc_sel_2_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_0_bits_vc_sel_1_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_0_bits_vc_sel_1_1; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_0_bits_vc_sel_1_2; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_0_bits_vc_sel_1_3; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_0_bits_vc_sel_0_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_0_bits_vc_sel_0_1; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_0_bits_vc_sel_0_2; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_0_bits_vc_sel_0_3; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_0_bits_tail; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_1_ready; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_1_valid; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_1_bits_vc_sel_2_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_1_bits_vc_sel_1_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_1_bits_vc_sel_1_1; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_1_bits_vc_sel_1_2; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_1_bits_vc_sel_1_3; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_1_bits_vc_sel_0_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_1_bits_vc_sel_0_1; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_1_bits_vc_sel_0_2; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_1_bits_vc_sel_0_3; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_1_bits_tail; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_2_ready; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_2_valid; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_2_bits_vc_sel_2_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_2_bits_vc_sel_1_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_2_bits_vc_sel_1_1; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_2_bits_vc_sel_1_2; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_2_bits_vc_sel_1_3; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_2_bits_vc_sel_0_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_2_bits_vc_sel_0_1; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_2_bits_vc_sel_0_2; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_2_bits_vc_sel_0_3; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_2_bits_tail; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_out_0_valid; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_out_0_bits_vc_sel_2_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_out_0_bits_vc_sel_1_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_out_0_bits_vc_sel_1_1; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_out_0_bits_vc_sel_1_2; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_out_0_bits_vc_sel_1_3; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_out_0_bits_vc_sel_0_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_out_0_bits_vc_sel_0_1; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_out_0_bits_vc_sel_0_2; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_out_0_bits_vc_sel_0_3; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_out_0_bits_tail; // @[SwitchAllocator.scala 83:45]
  wire [2:0] arbs_1_io_chosen_oh_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_clock; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_reset; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_in_0_ready; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_in_0_valid; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_in_0_bits_vc_sel_2_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_in_0_bits_vc_sel_1_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_in_0_bits_vc_sel_1_1; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_in_0_bits_vc_sel_1_2; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_in_0_bits_vc_sel_1_3; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_in_0_bits_vc_sel_0_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_in_0_bits_vc_sel_0_1; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_in_0_bits_vc_sel_0_2; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_in_0_bits_vc_sel_0_3; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_in_0_bits_tail; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_in_1_ready; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_in_1_valid; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_in_1_bits_vc_sel_2_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_in_1_bits_vc_sel_1_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_in_1_bits_vc_sel_1_1; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_in_1_bits_vc_sel_1_2; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_in_1_bits_vc_sel_1_3; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_in_1_bits_vc_sel_0_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_in_1_bits_vc_sel_0_1; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_in_1_bits_vc_sel_0_2; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_in_1_bits_vc_sel_0_3; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_in_1_bits_tail; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_in_2_ready; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_in_2_valid; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_in_2_bits_vc_sel_2_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_in_2_bits_vc_sel_1_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_in_2_bits_vc_sel_1_1; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_in_2_bits_vc_sel_1_2; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_in_2_bits_vc_sel_1_3; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_in_2_bits_vc_sel_0_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_in_2_bits_vc_sel_0_1; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_in_2_bits_vc_sel_0_2; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_in_2_bits_vc_sel_0_3; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_in_2_bits_tail; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_out_0_valid; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_out_0_bits_vc_sel_2_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_out_0_bits_vc_sel_1_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_out_0_bits_vc_sel_1_1; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_out_0_bits_vc_sel_1_2; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_out_0_bits_vc_sel_1_3; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_out_0_bits_vc_sel_0_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_out_0_bits_vc_sel_0_1; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_out_0_bits_vc_sel_0_2; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_out_0_bits_vc_sel_0_3; // @[SwitchAllocator.scala 83:45]
  wire  arbs_2_io_out_0_bits_tail; // @[SwitchAllocator.scala 83:45]
  wire [2:0] arbs_2_io_chosen_oh_0; // @[SwitchAllocator.scala 83:45]
  wire  fires__0 = arbs_0_io_in_0_ready & arbs_0_io_in_0_valid; // @[Decoupled.scala 51:35]
  wire  fires__1 = arbs_1_io_in_0_ready & arbs_1_io_in_0_valid; // @[Decoupled.scala 51:35]
  wire  fires__2 = arbs_2_io_in_0_ready & arbs_2_io_in_0_valid; // @[Decoupled.scala 51:35]
  wire  fires_1_0 = arbs_0_io_in_1_ready & arbs_0_io_in_1_valid; // @[Decoupled.scala 51:35]
  wire  fires_1_1 = arbs_1_io_in_1_ready & arbs_1_io_in_1_valid; // @[Decoupled.scala 51:35]
  wire  fires_1_2 = arbs_2_io_in_1_ready & arbs_2_io_in_1_valid; // @[Decoupled.scala 51:35]
  wire  fires_2_0 = arbs_0_io_in_2_ready & arbs_0_io_in_2_valid; // @[Decoupled.scala 51:35]
  wire  fires_2_1 = arbs_1_io_in_2_ready & arbs_1_io_in_2_valid; // @[Decoupled.scala 51:35]
  wire  fires_2_2 = arbs_2_io_in_2_ready & arbs_2_io_in_2_valid; // @[Decoupled.scala 51:35]
  SwitchArbiter_2 arbs_0 ( // @[SwitchAllocator.scala 83:45]
    .clock(arbs_0_clock),
    .reset(arbs_0_reset),
    .io_in_0_ready(arbs_0_io_in_0_ready),
    .io_in_0_valid(arbs_0_io_in_0_valid),
    .io_in_0_bits_vc_sel_2_0(arbs_0_io_in_0_bits_vc_sel_2_0),
    .io_in_0_bits_vc_sel_1_0(arbs_0_io_in_0_bits_vc_sel_1_0),
    .io_in_0_bits_vc_sel_1_1(arbs_0_io_in_0_bits_vc_sel_1_1),
    .io_in_0_bits_vc_sel_1_2(arbs_0_io_in_0_bits_vc_sel_1_2),
    .io_in_0_bits_vc_sel_1_3(arbs_0_io_in_0_bits_vc_sel_1_3),
    .io_in_0_bits_vc_sel_0_0(arbs_0_io_in_0_bits_vc_sel_0_0),
    .io_in_0_bits_vc_sel_0_1(arbs_0_io_in_0_bits_vc_sel_0_1),
    .io_in_0_bits_vc_sel_0_2(arbs_0_io_in_0_bits_vc_sel_0_2),
    .io_in_0_bits_vc_sel_0_3(arbs_0_io_in_0_bits_vc_sel_0_3),
    .io_in_0_bits_tail(arbs_0_io_in_0_bits_tail),
    .io_in_1_ready(arbs_0_io_in_1_ready),
    .io_in_1_valid(arbs_0_io_in_1_valid),
    .io_in_1_bits_vc_sel_2_0(arbs_0_io_in_1_bits_vc_sel_2_0),
    .io_in_1_bits_vc_sel_1_0(arbs_0_io_in_1_bits_vc_sel_1_0),
    .io_in_1_bits_vc_sel_1_1(arbs_0_io_in_1_bits_vc_sel_1_1),
    .io_in_1_bits_vc_sel_1_2(arbs_0_io_in_1_bits_vc_sel_1_2),
    .io_in_1_bits_vc_sel_1_3(arbs_0_io_in_1_bits_vc_sel_1_3),
    .io_in_1_bits_vc_sel_0_0(arbs_0_io_in_1_bits_vc_sel_0_0),
    .io_in_1_bits_vc_sel_0_1(arbs_0_io_in_1_bits_vc_sel_0_1),
    .io_in_1_bits_vc_sel_0_2(arbs_0_io_in_1_bits_vc_sel_0_2),
    .io_in_1_bits_vc_sel_0_3(arbs_0_io_in_1_bits_vc_sel_0_3),
    .io_in_1_bits_tail(arbs_0_io_in_1_bits_tail),
    .io_in_2_ready(arbs_0_io_in_2_ready),
    .io_in_2_valid(arbs_0_io_in_2_valid),
    .io_in_2_bits_vc_sel_2_0(arbs_0_io_in_2_bits_vc_sel_2_0),
    .io_in_2_bits_vc_sel_1_0(arbs_0_io_in_2_bits_vc_sel_1_0),
    .io_in_2_bits_vc_sel_1_1(arbs_0_io_in_2_bits_vc_sel_1_1),
    .io_in_2_bits_vc_sel_1_2(arbs_0_io_in_2_bits_vc_sel_1_2),
    .io_in_2_bits_vc_sel_1_3(arbs_0_io_in_2_bits_vc_sel_1_3),
    .io_in_2_bits_vc_sel_0_0(arbs_0_io_in_2_bits_vc_sel_0_0),
    .io_in_2_bits_vc_sel_0_1(arbs_0_io_in_2_bits_vc_sel_0_1),
    .io_in_2_bits_vc_sel_0_2(arbs_0_io_in_2_bits_vc_sel_0_2),
    .io_in_2_bits_vc_sel_0_3(arbs_0_io_in_2_bits_vc_sel_0_3),
    .io_in_2_bits_tail(arbs_0_io_in_2_bits_tail),
    .io_out_0_valid(arbs_0_io_out_0_valid),
    .io_out_0_bits_vc_sel_2_0(arbs_0_io_out_0_bits_vc_sel_2_0),
    .io_out_0_bits_vc_sel_1_0(arbs_0_io_out_0_bits_vc_sel_1_0),
    .io_out_0_bits_vc_sel_1_1(arbs_0_io_out_0_bits_vc_sel_1_1),
    .io_out_0_bits_vc_sel_1_2(arbs_0_io_out_0_bits_vc_sel_1_2),
    .io_out_0_bits_vc_sel_1_3(arbs_0_io_out_0_bits_vc_sel_1_3),
    .io_out_0_bits_vc_sel_0_0(arbs_0_io_out_0_bits_vc_sel_0_0),
    .io_out_0_bits_vc_sel_0_1(arbs_0_io_out_0_bits_vc_sel_0_1),
    .io_out_0_bits_vc_sel_0_2(arbs_0_io_out_0_bits_vc_sel_0_2),
    .io_out_0_bits_vc_sel_0_3(arbs_0_io_out_0_bits_vc_sel_0_3),
    .io_out_0_bits_tail(arbs_0_io_out_0_bits_tail),
    .io_chosen_oh_0(arbs_0_io_chosen_oh_0)
  );
  SwitchArbiter_2 arbs_1 ( // @[SwitchAllocator.scala 83:45]
    .clock(arbs_1_clock),
    .reset(arbs_1_reset),
    .io_in_0_ready(arbs_1_io_in_0_ready),
    .io_in_0_valid(arbs_1_io_in_0_valid),
    .io_in_0_bits_vc_sel_2_0(arbs_1_io_in_0_bits_vc_sel_2_0),
    .io_in_0_bits_vc_sel_1_0(arbs_1_io_in_0_bits_vc_sel_1_0),
    .io_in_0_bits_vc_sel_1_1(arbs_1_io_in_0_bits_vc_sel_1_1),
    .io_in_0_bits_vc_sel_1_2(arbs_1_io_in_0_bits_vc_sel_1_2),
    .io_in_0_bits_vc_sel_1_3(arbs_1_io_in_0_bits_vc_sel_1_3),
    .io_in_0_bits_vc_sel_0_0(arbs_1_io_in_0_bits_vc_sel_0_0),
    .io_in_0_bits_vc_sel_0_1(arbs_1_io_in_0_bits_vc_sel_0_1),
    .io_in_0_bits_vc_sel_0_2(arbs_1_io_in_0_bits_vc_sel_0_2),
    .io_in_0_bits_vc_sel_0_3(arbs_1_io_in_0_bits_vc_sel_0_3),
    .io_in_0_bits_tail(arbs_1_io_in_0_bits_tail),
    .io_in_1_ready(arbs_1_io_in_1_ready),
    .io_in_1_valid(arbs_1_io_in_1_valid),
    .io_in_1_bits_vc_sel_2_0(arbs_1_io_in_1_bits_vc_sel_2_0),
    .io_in_1_bits_vc_sel_1_0(arbs_1_io_in_1_bits_vc_sel_1_0),
    .io_in_1_bits_vc_sel_1_1(arbs_1_io_in_1_bits_vc_sel_1_1),
    .io_in_1_bits_vc_sel_1_2(arbs_1_io_in_1_bits_vc_sel_1_2),
    .io_in_1_bits_vc_sel_1_3(arbs_1_io_in_1_bits_vc_sel_1_3),
    .io_in_1_bits_vc_sel_0_0(arbs_1_io_in_1_bits_vc_sel_0_0),
    .io_in_1_bits_vc_sel_0_1(arbs_1_io_in_1_bits_vc_sel_0_1),
    .io_in_1_bits_vc_sel_0_2(arbs_1_io_in_1_bits_vc_sel_0_2),
    .io_in_1_bits_vc_sel_0_3(arbs_1_io_in_1_bits_vc_sel_0_3),
    .io_in_1_bits_tail(arbs_1_io_in_1_bits_tail),
    .io_in_2_ready(arbs_1_io_in_2_ready),
    .io_in_2_valid(arbs_1_io_in_2_valid),
    .io_in_2_bits_vc_sel_2_0(arbs_1_io_in_2_bits_vc_sel_2_0),
    .io_in_2_bits_vc_sel_1_0(arbs_1_io_in_2_bits_vc_sel_1_0),
    .io_in_2_bits_vc_sel_1_1(arbs_1_io_in_2_bits_vc_sel_1_1),
    .io_in_2_bits_vc_sel_1_2(arbs_1_io_in_2_bits_vc_sel_1_2),
    .io_in_2_bits_vc_sel_1_3(arbs_1_io_in_2_bits_vc_sel_1_3),
    .io_in_2_bits_vc_sel_0_0(arbs_1_io_in_2_bits_vc_sel_0_0),
    .io_in_2_bits_vc_sel_0_1(arbs_1_io_in_2_bits_vc_sel_0_1),
    .io_in_2_bits_vc_sel_0_2(arbs_1_io_in_2_bits_vc_sel_0_2),
    .io_in_2_bits_vc_sel_0_3(arbs_1_io_in_2_bits_vc_sel_0_3),
    .io_in_2_bits_tail(arbs_1_io_in_2_bits_tail),
    .io_out_0_valid(arbs_1_io_out_0_valid),
    .io_out_0_bits_vc_sel_2_0(arbs_1_io_out_0_bits_vc_sel_2_0),
    .io_out_0_bits_vc_sel_1_0(arbs_1_io_out_0_bits_vc_sel_1_0),
    .io_out_0_bits_vc_sel_1_1(arbs_1_io_out_0_bits_vc_sel_1_1),
    .io_out_0_bits_vc_sel_1_2(arbs_1_io_out_0_bits_vc_sel_1_2),
    .io_out_0_bits_vc_sel_1_3(arbs_1_io_out_0_bits_vc_sel_1_3),
    .io_out_0_bits_vc_sel_0_0(arbs_1_io_out_0_bits_vc_sel_0_0),
    .io_out_0_bits_vc_sel_0_1(arbs_1_io_out_0_bits_vc_sel_0_1),
    .io_out_0_bits_vc_sel_0_2(arbs_1_io_out_0_bits_vc_sel_0_2),
    .io_out_0_bits_vc_sel_0_3(arbs_1_io_out_0_bits_vc_sel_0_3),
    .io_out_0_bits_tail(arbs_1_io_out_0_bits_tail),
    .io_chosen_oh_0(arbs_1_io_chosen_oh_0)
  );
  SwitchArbiter_2 arbs_2 ( // @[SwitchAllocator.scala 83:45]
    .clock(arbs_2_clock),
    .reset(arbs_2_reset),
    .io_in_0_ready(arbs_2_io_in_0_ready),
    .io_in_0_valid(arbs_2_io_in_0_valid),
    .io_in_0_bits_vc_sel_2_0(arbs_2_io_in_0_bits_vc_sel_2_0),
    .io_in_0_bits_vc_sel_1_0(arbs_2_io_in_0_bits_vc_sel_1_0),
    .io_in_0_bits_vc_sel_1_1(arbs_2_io_in_0_bits_vc_sel_1_1),
    .io_in_0_bits_vc_sel_1_2(arbs_2_io_in_0_bits_vc_sel_1_2),
    .io_in_0_bits_vc_sel_1_3(arbs_2_io_in_0_bits_vc_sel_1_3),
    .io_in_0_bits_vc_sel_0_0(arbs_2_io_in_0_bits_vc_sel_0_0),
    .io_in_0_bits_vc_sel_0_1(arbs_2_io_in_0_bits_vc_sel_0_1),
    .io_in_0_bits_vc_sel_0_2(arbs_2_io_in_0_bits_vc_sel_0_2),
    .io_in_0_bits_vc_sel_0_3(arbs_2_io_in_0_bits_vc_sel_0_3),
    .io_in_0_bits_tail(arbs_2_io_in_0_bits_tail),
    .io_in_1_ready(arbs_2_io_in_1_ready),
    .io_in_1_valid(arbs_2_io_in_1_valid),
    .io_in_1_bits_vc_sel_2_0(arbs_2_io_in_1_bits_vc_sel_2_0),
    .io_in_1_bits_vc_sel_1_0(arbs_2_io_in_1_bits_vc_sel_1_0),
    .io_in_1_bits_vc_sel_1_1(arbs_2_io_in_1_bits_vc_sel_1_1),
    .io_in_1_bits_vc_sel_1_2(arbs_2_io_in_1_bits_vc_sel_1_2),
    .io_in_1_bits_vc_sel_1_3(arbs_2_io_in_1_bits_vc_sel_1_3),
    .io_in_1_bits_vc_sel_0_0(arbs_2_io_in_1_bits_vc_sel_0_0),
    .io_in_1_bits_vc_sel_0_1(arbs_2_io_in_1_bits_vc_sel_0_1),
    .io_in_1_bits_vc_sel_0_2(arbs_2_io_in_1_bits_vc_sel_0_2),
    .io_in_1_bits_vc_sel_0_3(arbs_2_io_in_1_bits_vc_sel_0_3),
    .io_in_1_bits_tail(arbs_2_io_in_1_bits_tail),
    .io_in_2_ready(arbs_2_io_in_2_ready),
    .io_in_2_valid(arbs_2_io_in_2_valid),
    .io_in_2_bits_vc_sel_2_0(arbs_2_io_in_2_bits_vc_sel_2_0),
    .io_in_2_bits_vc_sel_1_0(arbs_2_io_in_2_bits_vc_sel_1_0),
    .io_in_2_bits_vc_sel_1_1(arbs_2_io_in_2_bits_vc_sel_1_1),
    .io_in_2_bits_vc_sel_1_2(arbs_2_io_in_2_bits_vc_sel_1_2),
    .io_in_2_bits_vc_sel_1_3(arbs_2_io_in_2_bits_vc_sel_1_3),
    .io_in_2_bits_vc_sel_0_0(arbs_2_io_in_2_bits_vc_sel_0_0),
    .io_in_2_bits_vc_sel_0_1(arbs_2_io_in_2_bits_vc_sel_0_1),
    .io_in_2_bits_vc_sel_0_2(arbs_2_io_in_2_bits_vc_sel_0_2),
    .io_in_2_bits_vc_sel_0_3(arbs_2_io_in_2_bits_vc_sel_0_3),
    .io_in_2_bits_tail(arbs_2_io_in_2_bits_tail),
    .io_out_0_valid(arbs_2_io_out_0_valid),
    .io_out_0_bits_vc_sel_2_0(arbs_2_io_out_0_bits_vc_sel_2_0),
    .io_out_0_bits_vc_sel_1_0(arbs_2_io_out_0_bits_vc_sel_1_0),
    .io_out_0_bits_vc_sel_1_1(arbs_2_io_out_0_bits_vc_sel_1_1),
    .io_out_0_bits_vc_sel_1_2(arbs_2_io_out_0_bits_vc_sel_1_2),
    .io_out_0_bits_vc_sel_1_3(arbs_2_io_out_0_bits_vc_sel_1_3),
    .io_out_0_bits_vc_sel_0_0(arbs_2_io_out_0_bits_vc_sel_0_0),
    .io_out_0_bits_vc_sel_0_1(arbs_2_io_out_0_bits_vc_sel_0_1),
    .io_out_0_bits_vc_sel_0_2(arbs_2_io_out_0_bits_vc_sel_0_2),
    .io_out_0_bits_vc_sel_0_3(arbs_2_io_out_0_bits_vc_sel_0_3),
    .io_out_0_bits_tail(arbs_2_io_out_0_bits_tail),
    .io_chosen_oh_0(arbs_2_io_chosen_oh_0)
  );
  assign io_req_2_0_ready = fires_2_0 | fires_2_1 | fires_2_2; // @[SwitchAllocator.scala 99:30]
  assign io_req_1_0_ready = fires_1_0 | fires_1_1 | fires_1_2; // @[SwitchAllocator.scala 99:30]
  assign io_req_0_0_ready = fires__0 | fires__1 | fires__2; // @[SwitchAllocator.scala 99:30]
  assign io_credit_alloc_2_0_alloc = arbs_2_io_out_0_valid & arbs_2_io_out_0_bits_vc_sel_2_0; // @[SwitchAllocator.scala 120:33]
  assign io_credit_alloc_2_0_tail = arbs_2_io_out_0_valid & arbs_2_io_out_0_bits_vc_sel_2_0 & arbs_2_io_out_0_bits_tail; // @[SwitchAllocator.scala 120:67 122:21 116:44]
  assign io_credit_alloc_1_0_alloc = arbs_1_io_out_0_valid & arbs_1_io_out_0_bits_vc_sel_1_0; // @[SwitchAllocator.scala 120:33]
  assign io_credit_alloc_1_1_alloc = arbs_1_io_out_0_valid & arbs_1_io_out_0_bits_vc_sel_1_1; // @[SwitchAllocator.scala 120:33]
  assign io_credit_alloc_1_2_alloc = arbs_1_io_out_0_valid & arbs_1_io_out_0_bits_vc_sel_1_2; // @[SwitchAllocator.scala 120:33]
  assign io_credit_alloc_1_3_alloc = arbs_1_io_out_0_valid & arbs_1_io_out_0_bits_vc_sel_1_3; // @[SwitchAllocator.scala 120:33]
  assign io_credit_alloc_0_0_alloc = arbs_0_io_out_0_valid & arbs_0_io_out_0_bits_vc_sel_0_0; // @[SwitchAllocator.scala 120:33]
  assign io_credit_alloc_0_1_alloc = arbs_0_io_out_0_valid & arbs_0_io_out_0_bits_vc_sel_0_1; // @[SwitchAllocator.scala 120:33]
  assign io_credit_alloc_0_2_alloc = arbs_0_io_out_0_valid & arbs_0_io_out_0_bits_vc_sel_0_2; // @[SwitchAllocator.scala 120:33]
  assign io_credit_alloc_0_3_alloc = arbs_0_io_out_0_valid & arbs_0_io_out_0_bits_vc_sel_0_3; // @[SwitchAllocator.scala 120:33]
  assign io_switch_sel_2_0_2_0 = arbs_2_io_in_2_valid & arbs_2_io_chosen_oh_0[2] & arbs_2_io_out_0_valid; // @[SwitchAllocator.scala 108:97]
  assign io_switch_sel_2_0_1_0 = arbs_2_io_in_1_valid & arbs_2_io_chosen_oh_0[1] & arbs_2_io_out_0_valid; // @[SwitchAllocator.scala 108:97]
  assign io_switch_sel_2_0_0_0 = arbs_2_io_in_0_valid & arbs_2_io_chosen_oh_0[0] & arbs_2_io_out_0_valid; // @[SwitchAllocator.scala 108:97]
  assign io_switch_sel_1_0_2_0 = arbs_1_io_in_2_valid & arbs_1_io_chosen_oh_0[2] & arbs_1_io_out_0_valid; // @[SwitchAllocator.scala 108:97]
  assign io_switch_sel_1_0_1_0 = arbs_1_io_in_1_valid & arbs_1_io_chosen_oh_0[1] & arbs_1_io_out_0_valid; // @[SwitchAllocator.scala 108:97]
  assign io_switch_sel_1_0_0_0 = arbs_1_io_in_0_valid & arbs_1_io_chosen_oh_0[0] & arbs_1_io_out_0_valid; // @[SwitchAllocator.scala 108:97]
  assign io_switch_sel_0_0_2_0 = arbs_0_io_in_2_valid & arbs_0_io_chosen_oh_0[2] & arbs_0_io_out_0_valid; // @[SwitchAllocator.scala 108:97]
  assign io_switch_sel_0_0_1_0 = arbs_0_io_in_1_valid & arbs_0_io_chosen_oh_0[1] & arbs_0_io_out_0_valid; // @[SwitchAllocator.scala 108:97]
  assign io_switch_sel_0_0_0_0 = arbs_0_io_in_0_valid & arbs_0_io_chosen_oh_0[0] & arbs_0_io_out_0_valid; // @[SwitchAllocator.scala 108:97]
  assign arbs_0_clock = clock;
  assign arbs_0_reset = reset;
  assign arbs_0_io_in_0_valid = io_req_0_0_valid & (io_req_0_0_bits_vc_sel_0_0 | io_req_0_0_bits_vc_sel_0_1 |
    io_req_0_0_bits_vc_sel_0_2 | io_req_0_0_bits_vc_sel_0_3); // @[SwitchAllocator.scala 95:37]
  assign arbs_0_io_in_0_bits_vc_sel_2_0 = io_req_0_0_bits_vc_sel_2_0; // @[SwitchAllocator.scala 96:25]
  assign arbs_0_io_in_0_bits_vc_sel_1_0 = io_req_0_0_bits_vc_sel_1_0; // @[SwitchAllocator.scala 96:25]
  assign arbs_0_io_in_0_bits_vc_sel_1_1 = io_req_0_0_bits_vc_sel_1_1; // @[SwitchAllocator.scala 96:25]
  assign arbs_0_io_in_0_bits_vc_sel_1_2 = io_req_0_0_bits_vc_sel_1_2; // @[SwitchAllocator.scala 96:25]
  assign arbs_0_io_in_0_bits_vc_sel_1_3 = io_req_0_0_bits_vc_sel_1_3; // @[SwitchAllocator.scala 96:25]
  assign arbs_0_io_in_0_bits_vc_sel_0_0 = io_req_0_0_bits_vc_sel_0_0; // @[SwitchAllocator.scala 96:25]
  assign arbs_0_io_in_0_bits_vc_sel_0_1 = io_req_0_0_bits_vc_sel_0_1; // @[SwitchAllocator.scala 96:25]
  assign arbs_0_io_in_0_bits_vc_sel_0_2 = io_req_0_0_bits_vc_sel_0_2; // @[SwitchAllocator.scala 96:25]
  assign arbs_0_io_in_0_bits_vc_sel_0_3 = io_req_0_0_bits_vc_sel_0_3; // @[SwitchAllocator.scala 96:25]
  assign arbs_0_io_in_0_bits_tail = io_req_0_0_bits_tail; // @[SwitchAllocator.scala 96:25]
  assign arbs_0_io_in_1_valid = io_req_1_0_valid & (io_req_1_0_bits_vc_sel_0_0 | io_req_1_0_bits_vc_sel_0_1 |
    io_req_1_0_bits_vc_sel_0_2 | io_req_1_0_bits_vc_sel_0_3); // @[SwitchAllocator.scala 95:37]
  assign arbs_0_io_in_1_bits_vc_sel_2_0 = io_req_1_0_bits_vc_sel_2_0; // @[SwitchAllocator.scala 96:25]
  assign arbs_0_io_in_1_bits_vc_sel_1_0 = io_req_1_0_bits_vc_sel_1_0; // @[SwitchAllocator.scala 96:25]
  assign arbs_0_io_in_1_bits_vc_sel_1_1 = io_req_1_0_bits_vc_sel_1_1; // @[SwitchAllocator.scala 96:25]
  assign arbs_0_io_in_1_bits_vc_sel_1_2 = io_req_1_0_bits_vc_sel_1_2; // @[SwitchAllocator.scala 96:25]
  assign arbs_0_io_in_1_bits_vc_sel_1_3 = io_req_1_0_bits_vc_sel_1_3; // @[SwitchAllocator.scala 96:25]
  assign arbs_0_io_in_1_bits_vc_sel_0_0 = io_req_1_0_bits_vc_sel_0_0; // @[SwitchAllocator.scala 96:25]
  assign arbs_0_io_in_1_bits_vc_sel_0_1 = io_req_1_0_bits_vc_sel_0_1; // @[SwitchAllocator.scala 96:25]
  assign arbs_0_io_in_1_bits_vc_sel_0_2 = io_req_1_0_bits_vc_sel_0_2; // @[SwitchAllocator.scala 96:25]
  assign arbs_0_io_in_1_bits_vc_sel_0_3 = io_req_1_0_bits_vc_sel_0_3; // @[SwitchAllocator.scala 96:25]
  assign arbs_0_io_in_1_bits_tail = io_req_1_0_bits_tail; // @[SwitchAllocator.scala 96:25]
  assign arbs_0_io_in_2_valid = io_req_2_0_valid & (io_req_2_0_bits_vc_sel_0_0 | io_req_2_0_bits_vc_sel_0_1 |
    io_req_2_0_bits_vc_sel_0_2 | io_req_2_0_bits_vc_sel_0_3); // @[SwitchAllocator.scala 95:37]
  assign arbs_0_io_in_2_bits_vc_sel_2_0 = io_req_2_0_bits_vc_sel_2_0; // @[SwitchAllocator.scala 96:25]
  assign arbs_0_io_in_2_bits_vc_sel_1_0 = io_req_2_0_bits_vc_sel_1_0; // @[SwitchAllocator.scala 96:25]
  assign arbs_0_io_in_2_bits_vc_sel_1_1 = io_req_2_0_bits_vc_sel_1_1; // @[SwitchAllocator.scala 96:25]
  assign arbs_0_io_in_2_bits_vc_sel_1_2 = io_req_2_0_bits_vc_sel_1_2; // @[SwitchAllocator.scala 96:25]
  assign arbs_0_io_in_2_bits_vc_sel_1_3 = io_req_2_0_bits_vc_sel_1_3; // @[SwitchAllocator.scala 96:25]
  assign arbs_0_io_in_2_bits_vc_sel_0_0 = io_req_2_0_bits_vc_sel_0_0; // @[SwitchAllocator.scala 96:25]
  assign arbs_0_io_in_2_bits_vc_sel_0_1 = io_req_2_0_bits_vc_sel_0_1; // @[SwitchAllocator.scala 96:25]
  assign arbs_0_io_in_2_bits_vc_sel_0_2 = io_req_2_0_bits_vc_sel_0_2; // @[SwitchAllocator.scala 96:25]
  assign arbs_0_io_in_2_bits_vc_sel_0_3 = io_req_2_0_bits_vc_sel_0_3; // @[SwitchAllocator.scala 96:25]
  assign arbs_0_io_in_2_bits_tail = io_req_2_0_bits_tail; // @[SwitchAllocator.scala 96:25]
  assign arbs_1_clock = clock;
  assign arbs_1_reset = reset;
  assign arbs_1_io_in_0_valid = io_req_0_0_valid & (io_req_0_0_bits_vc_sel_1_0 | io_req_0_0_bits_vc_sel_1_1 |
    io_req_0_0_bits_vc_sel_1_2 | io_req_0_0_bits_vc_sel_1_3); // @[SwitchAllocator.scala 95:37]
  assign arbs_1_io_in_0_bits_vc_sel_2_0 = io_req_0_0_bits_vc_sel_2_0; // @[SwitchAllocator.scala 96:25]
  assign arbs_1_io_in_0_bits_vc_sel_1_0 = io_req_0_0_bits_vc_sel_1_0; // @[SwitchAllocator.scala 96:25]
  assign arbs_1_io_in_0_bits_vc_sel_1_1 = io_req_0_0_bits_vc_sel_1_1; // @[SwitchAllocator.scala 96:25]
  assign arbs_1_io_in_0_bits_vc_sel_1_2 = io_req_0_0_bits_vc_sel_1_2; // @[SwitchAllocator.scala 96:25]
  assign arbs_1_io_in_0_bits_vc_sel_1_3 = io_req_0_0_bits_vc_sel_1_3; // @[SwitchAllocator.scala 96:25]
  assign arbs_1_io_in_0_bits_vc_sel_0_0 = io_req_0_0_bits_vc_sel_0_0; // @[SwitchAllocator.scala 96:25]
  assign arbs_1_io_in_0_bits_vc_sel_0_1 = io_req_0_0_bits_vc_sel_0_1; // @[SwitchAllocator.scala 96:25]
  assign arbs_1_io_in_0_bits_vc_sel_0_2 = io_req_0_0_bits_vc_sel_0_2; // @[SwitchAllocator.scala 96:25]
  assign arbs_1_io_in_0_bits_vc_sel_0_3 = io_req_0_0_bits_vc_sel_0_3; // @[SwitchAllocator.scala 96:25]
  assign arbs_1_io_in_0_bits_tail = io_req_0_0_bits_tail; // @[SwitchAllocator.scala 96:25]
  assign arbs_1_io_in_1_valid = io_req_1_0_valid & (io_req_1_0_bits_vc_sel_1_0 | io_req_1_0_bits_vc_sel_1_1 |
    io_req_1_0_bits_vc_sel_1_2 | io_req_1_0_bits_vc_sel_1_3); // @[SwitchAllocator.scala 95:37]
  assign arbs_1_io_in_1_bits_vc_sel_2_0 = io_req_1_0_bits_vc_sel_2_0; // @[SwitchAllocator.scala 96:25]
  assign arbs_1_io_in_1_bits_vc_sel_1_0 = io_req_1_0_bits_vc_sel_1_0; // @[SwitchAllocator.scala 96:25]
  assign arbs_1_io_in_1_bits_vc_sel_1_1 = io_req_1_0_bits_vc_sel_1_1; // @[SwitchAllocator.scala 96:25]
  assign arbs_1_io_in_1_bits_vc_sel_1_2 = io_req_1_0_bits_vc_sel_1_2; // @[SwitchAllocator.scala 96:25]
  assign arbs_1_io_in_1_bits_vc_sel_1_3 = io_req_1_0_bits_vc_sel_1_3; // @[SwitchAllocator.scala 96:25]
  assign arbs_1_io_in_1_bits_vc_sel_0_0 = io_req_1_0_bits_vc_sel_0_0; // @[SwitchAllocator.scala 96:25]
  assign arbs_1_io_in_1_bits_vc_sel_0_1 = io_req_1_0_bits_vc_sel_0_1; // @[SwitchAllocator.scala 96:25]
  assign arbs_1_io_in_1_bits_vc_sel_0_2 = io_req_1_0_bits_vc_sel_0_2; // @[SwitchAllocator.scala 96:25]
  assign arbs_1_io_in_1_bits_vc_sel_0_3 = io_req_1_0_bits_vc_sel_0_3; // @[SwitchAllocator.scala 96:25]
  assign arbs_1_io_in_1_bits_tail = io_req_1_0_bits_tail; // @[SwitchAllocator.scala 96:25]
  assign arbs_1_io_in_2_valid = io_req_2_0_valid & (io_req_2_0_bits_vc_sel_1_0 | io_req_2_0_bits_vc_sel_1_1 |
    io_req_2_0_bits_vc_sel_1_2 | io_req_2_0_bits_vc_sel_1_3); // @[SwitchAllocator.scala 95:37]
  assign arbs_1_io_in_2_bits_vc_sel_2_0 = io_req_2_0_bits_vc_sel_2_0; // @[SwitchAllocator.scala 96:25]
  assign arbs_1_io_in_2_bits_vc_sel_1_0 = io_req_2_0_bits_vc_sel_1_0; // @[SwitchAllocator.scala 96:25]
  assign arbs_1_io_in_2_bits_vc_sel_1_1 = io_req_2_0_bits_vc_sel_1_1; // @[SwitchAllocator.scala 96:25]
  assign arbs_1_io_in_2_bits_vc_sel_1_2 = io_req_2_0_bits_vc_sel_1_2; // @[SwitchAllocator.scala 96:25]
  assign arbs_1_io_in_2_bits_vc_sel_1_3 = io_req_2_0_bits_vc_sel_1_3; // @[SwitchAllocator.scala 96:25]
  assign arbs_1_io_in_2_bits_vc_sel_0_0 = io_req_2_0_bits_vc_sel_0_0; // @[SwitchAllocator.scala 96:25]
  assign arbs_1_io_in_2_bits_vc_sel_0_1 = io_req_2_0_bits_vc_sel_0_1; // @[SwitchAllocator.scala 96:25]
  assign arbs_1_io_in_2_bits_vc_sel_0_2 = io_req_2_0_bits_vc_sel_0_2; // @[SwitchAllocator.scala 96:25]
  assign arbs_1_io_in_2_bits_vc_sel_0_3 = io_req_2_0_bits_vc_sel_0_3; // @[SwitchAllocator.scala 96:25]
  assign arbs_1_io_in_2_bits_tail = io_req_2_0_bits_tail; // @[SwitchAllocator.scala 96:25]
  assign arbs_2_clock = clock;
  assign arbs_2_reset = reset;
  assign arbs_2_io_in_0_valid = io_req_0_0_valid & io_req_0_0_bits_vc_sel_2_0; // @[SwitchAllocator.scala 95:37]
  assign arbs_2_io_in_0_bits_vc_sel_2_0 = io_req_0_0_bits_vc_sel_2_0; // @[SwitchAllocator.scala 96:25]
  assign arbs_2_io_in_0_bits_vc_sel_1_0 = io_req_0_0_bits_vc_sel_1_0; // @[SwitchAllocator.scala 96:25]
  assign arbs_2_io_in_0_bits_vc_sel_1_1 = io_req_0_0_bits_vc_sel_1_1; // @[SwitchAllocator.scala 96:25]
  assign arbs_2_io_in_0_bits_vc_sel_1_2 = io_req_0_0_bits_vc_sel_1_2; // @[SwitchAllocator.scala 96:25]
  assign arbs_2_io_in_0_bits_vc_sel_1_3 = io_req_0_0_bits_vc_sel_1_3; // @[SwitchAllocator.scala 96:25]
  assign arbs_2_io_in_0_bits_vc_sel_0_0 = io_req_0_0_bits_vc_sel_0_0; // @[SwitchAllocator.scala 96:25]
  assign arbs_2_io_in_0_bits_vc_sel_0_1 = io_req_0_0_bits_vc_sel_0_1; // @[SwitchAllocator.scala 96:25]
  assign arbs_2_io_in_0_bits_vc_sel_0_2 = io_req_0_0_bits_vc_sel_0_2; // @[SwitchAllocator.scala 96:25]
  assign arbs_2_io_in_0_bits_vc_sel_0_3 = io_req_0_0_bits_vc_sel_0_3; // @[SwitchAllocator.scala 96:25]
  assign arbs_2_io_in_0_bits_tail = io_req_0_0_bits_tail; // @[SwitchAllocator.scala 96:25]
  assign arbs_2_io_in_1_valid = io_req_1_0_valid & io_req_1_0_bits_vc_sel_2_0; // @[SwitchAllocator.scala 95:37]
  assign arbs_2_io_in_1_bits_vc_sel_2_0 = io_req_1_0_bits_vc_sel_2_0; // @[SwitchAllocator.scala 96:25]
  assign arbs_2_io_in_1_bits_vc_sel_1_0 = io_req_1_0_bits_vc_sel_1_0; // @[SwitchAllocator.scala 96:25]
  assign arbs_2_io_in_1_bits_vc_sel_1_1 = io_req_1_0_bits_vc_sel_1_1; // @[SwitchAllocator.scala 96:25]
  assign arbs_2_io_in_1_bits_vc_sel_1_2 = io_req_1_0_bits_vc_sel_1_2; // @[SwitchAllocator.scala 96:25]
  assign arbs_2_io_in_1_bits_vc_sel_1_3 = io_req_1_0_bits_vc_sel_1_3; // @[SwitchAllocator.scala 96:25]
  assign arbs_2_io_in_1_bits_vc_sel_0_0 = io_req_1_0_bits_vc_sel_0_0; // @[SwitchAllocator.scala 96:25]
  assign arbs_2_io_in_1_bits_vc_sel_0_1 = io_req_1_0_bits_vc_sel_0_1; // @[SwitchAllocator.scala 96:25]
  assign arbs_2_io_in_1_bits_vc_sel_0_2 = io_req_1_0_bits_vc_sel_0_2; // @[SwitchAllocator.scala 96:25]
  assign arbs_2_io_in_1_bits_vc_sel_0_3 = io_req_1_0_bits_vc_sel_0_3; // @[SwitchAllocator.scala 96:25]
  assign arbs_2_io_in_1_bits_tail = io_req_1_0_bits_tail; // @[SwitchAllocator.scala 96:25]
  assign arbs_2_io_in_2_valid = io_req_2_0_valid & io_req_2_0_bits_vc_sel_2_0; // @[SwitchAllocator.scala 95:37]
  assign arbs_2_io_in_2_bits_vc_sel_2_0 = io_req_2_0_bits_vc_sel_2_0; // @[SwitchAllocator.scala 96:25]
  assign arbs_2_io_in_2_bits_vc_sel_1_0 = io_req_2_0_bits_vc_sel_1_0; // @[SwitchAllocator.scala 96:25]
  assign arbs_2_io_in_2_bits_vc_sel_1_1 = io_req_2_0_bits_vc_sel_1_1; // @[SwitchAllocator.scala 96:25]
  assign arbs_2_io_in_2_bits_vc_sel_1_2 = io_req_2_0_bits_vc_sel_1_2; // @[SwitchAllocator.scala 96:25]
  assign arbs_2_io_in_2_bits_vc_sel_1_3 = io_req_2_0_bits_vc_sel_1_3; // @[SwitchAllocator.scala 96:25]
  assign arbs_2_io_in_2_bits_vc_sel_0_0 = io_req_2_0_bits_vc_sel_0_0; // @[SwitchAllocator.scala 96:25]
  assign arbs_2_io_in_2_bits_vc_sel_0_1 = io_req_2_0_bits_vc_sel_0_1; // @[SwitchAllocator.scala 96:25]
  assign arbs_2_io_in_2_bits_vc_sel_0_2 = io_req_2_0_bits_vc_sel_0_2; // @[SwitchAllocator.scala 96:25]
  assign arbs_2_io_in_2_bits_vc_sel_0_3 = io_req_2_0_bits_vc_sel_0_3; // @[SwitchAllocator.scala 96:25]
  assign arbs_2_io_in_2_bits_tail = io_req_2_0_bits_tail; // @[SwitchAllocator.scala 96:25]
endmodule
module RotatingSingleVCAllocator(
  input   clock,
  input   reset,
  output  io_req_2_ready,
  input   io_req_2_valid,
  input   io_req_2_bits_vc_sel_2_0,
  input   io_req_2_bits_vc_sel_1_0,
  input   io_req_2_bits_vc_sel_1_1,
  input   io_req_2_bits_vc_sel_1_2,
  input   io_req_2_bits_vc_sel_1_3,
  input   io_req_2_bits_vc_sel_0_0,
  input   io_req_2_bits_vc_sel_0_1,
  input   io_req_2_bits_vc_sel_0_2,
  input   io_req_2_bits_vc_sel_0_3,
  output  io_req_1_ready,
  input   io_req_1_valid,
  input   io_req_1_bits_vc_sel_2_0,
  input   io_req_1_bits_vc_sel_1_0,
  input   io_req_1_bits_vc_sel_1_1,
  input   io_req_1_bits_vc_sel_1_2,
  input   io_req_1_bits_vc_sel_1_3,
  input   io_req_1_bits_vc_sel_0_0,
  input   io_req_1_bits_vc_sel_0_1,
  input   io_req_1_bits_vc_sel_0_2,
  input   io_req_1_bits_vc_sel_0_3,
  output  io_req_0_ready,
  input   io_req_0_valid,
  input   io_req_0_bits_vc_sel_2_0,
  input   io_req_0_bits_vc_sel_1_0,
  input   io_req_0_bits_vc_sel_1_1,
  input   io_req_0_bits_vc_sel_1_2,
  input   io_req_0_bits_vc_sel_1_3,
  input   io_req_0_bits_vc_sel_0_0,
  input   io_req_0_bits_vc_sel_0_1,
  input   io_req_0_bits_vc_sel_0_2,
  input   io_req_0_bits_vc_sel_0_3,
  output  io_resp_2_vc_sel_2_0,
  output  io_resp_2_vc_sel_1_0,
  output  io_resp_2_vc_sel_1_1,
  output  io_resp_2_vc_sel_1_2,
  output  io_resp_2_vc_sel_1_3,
  output  io_resp_2_vc_sel_0_0,
  output  io_resp_2_vc_sel_0_1,
  output  io_resp_2_vc_sel_0_2,
  output  io_resp_2_vc_sel_0_3,
  output  io_resp_1_vc_sel_2_0,
  output  io_resp_1_vc_sel_1_0,
  output  io_resp_1_vc_sel_1_1,
  output  io_resp_1_vc_sel_1_2,
  output  io_resp_1_vc_sel_1_3,
  output  io_resp_1_vc_sel_0_0,
  output  io_resp_1_vc_sel_0_1,
  output  io_resp_1_vc_sel_0_2,
  output  io_resp_1_vc_sel_0_3,
  output  io_resp_0_vc_sel_2_0,
  output  io_resp_0_vc_sel_1_0,
  output  io_resp_0_vc_sel_1_1,
  output  io_resp_0_vc_sel_1_2,
  output  io_resp_0_vc_sel_1_3,
  output  io_resp_0_vc_sel_0_0,
  output  io_resp_0_vc_sel_0_1,
  output  io_resp_0_vc_sel_0_2,
  output  io_resp_0_vc_sel_0_3,
  input   io_channel_status_2_0_occupied,
  input   io_channel_status_1_0_occupied,
  input   io_channel_status_1_1_occupied,
  input   io_channel_status_1_2_occupied,
  input   io_channel_status_1_3_occupied,
  input   io_channel_status_0_0_occupied,
  input   io_channel_status_0_1_occupied,
  input   io_channel_status_0_2_occupied,
  input   io_channel_status_0_3_occupied,
  output  io_out_allocs_2_0_alloc,
  output  io_out_allocs_1_0_alloc,
  output  io_out_allocs_1_1_alloc,
  output  io_out_allocs_1_2_alloc,
  output  io_out_allocs_1_3_alloc,
  output  io_out_allocs_0_0_alloc,
  output  io_out_allocs_0_1_alloc,
  output  io_out_allocs_0_2_alloc,
  output  io_out_allocs_0_3_alloc
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] mask; // @[SingleVCAllocator.scala 16:21]
  wire  in_arb_reqs_2_0_0 = io_req_2_bits_vc_sel_0_0 & ~io_channel_status_0_0_occupied; // @[SingleVCAllocator.scala 28:61]
  wire  in_arb_reqs_2_0_1 = io_req_2_bits_vc_sel_0_1 & ~io_channel_status_0_1_occupied; // @[SingleVCAllocator.scala 28:61]
  wire  in_arb_reqs_2_0_2 = io_req_2_bits_vc_sel_0_2 & ~io_channel_status_0_2_occupied; // @[SingleVCAllocator.scala 28:61]
  wire  in_arb_reqs_2_0_3 = io_req_2_bits_vc_sel_0_3 & ~io_channel_status_0_3_occupied; // @[SingleVCAllocator.scala 28:61]
  wire  in_arb_reqs_2_1_0 = io_req_2_bits_vc_sel_1_0 & ~io_channel_status_1_0_occupied; // @[SingleVCAllocator.scala 28:61]
  wire  in_arb_reqs_2_1_1 = io_req_2_bits_vc_sel_1_1 & ~io_channel_status_1_1_occupied; // @[SingleVCAllocator.scala 28:61]
  wire  in_arb_reqs_2_1_2 = io_req_2_bits_vc_sel_1_2 & ~io_channel_status_1_2_occupied; // @[SingleVCAllocator.scala 28:61]
  wire  in_arb_reqs_2_1_3 = io_req_2_bits_vc_sel_1_3 & ~io_channel_status_1_3_occupied; // @[SingleVCAllocator.scala 28:61]
  wire  in_arb_reqs_2_2_0 = io_req_2_bits_vc_sel_2_0 & ~io_channel_status_2_0_occupied; // @[SingleVCAllocator.scala 28:61]
  wire  _in_arb_vals_2_T_7 = in_arb_reqs_2_0_0 | in_arb_reqs_2_0_1 | in_arb_reqs_2_0_2 | in_arb_reqs_2_0_3 | (
    in_arb_reqs_2_1_0 | in_arb_reqs_2_1_1 | in_arb_reqs_2_1_2 | in_arb_reqs_2_1_3) | in_arb_reqs_2_2_0; // @[package.scala 73:59]
  wire  in_arb_vals_2 = io_req_2_valid & _in_arb_vals_2_T_7; // @[SingleVCAllocator.scala 32:39]
  wire  in_arb_reqs_1_0_0 = io_req_1_bits_vc_sel_0_0 & ~io_channel_status_0_0_occupied; // @[SingleVCAllocator.scala 28:61]
  wire  in_arb_reqs_1_0_1 = io_req_1_bits_vc_sel_0_1 & ~io_channel_status_0_1_occupied; // @[SingleVCAllocator.scala 28:61]
  wire  in_arb_reqs_1_0_2 = io_req_1_bits_vc_sel_0_2 & ~io_channel_status_0_2_occupied; // @[SingleVCAllocator.scala 28:61]
  wire  in_arb_reqs_1_0_3 = io_req_1_bits_vc_sel_0_3 & ~io_channel_status_0_3_occupied; // @[SingleVCAllocator.scala 28:61]
  wire  in_arb_reqs_1_1_0 = io_req_1_bits_vc_sel_1_0 & ~io_channel_status_1_0_occupied; // @[SingleVCAllocator.scala 28:61]
  wire  in_arb_reqs_1_1_1 = io_req_1_bits_vc_sel_1_1 & ~io_channel_status_1_1_occupied; // @[SingleVCAllocator.scala 28:61]
  wire  in_arb_reqs_1_1_2 = io_req_1_bits_vc_sel_1_2 & ~io_channel_status_1_2_occupied; // @[SingleVCAllocator.scala 28:61]
  wire  in_arb_reqs_1_1_3 = io_req_1_bits_vc_sel_1_3 & ~io_channel_status_1_3_occupied; // @[SingleVCAllocator.scala 28:61]
  wire  in_arb_reqs_1_2_0 = io_req_1_bits_vc_sel_2_0 & ~io_channel_status_2_0_occupied; // @[SingleVCAllocator.scala 28:61]
  wire  _in_arb_vals_1_T_7 = in_arb_reqs_1_0_0 | in_arb_reqs_1_0_1 | in_arb_reqs_1_0_2 | in_arb_reqs_1_0_3 | (
    in_arb_reqs_1_1_0 | in_arb_reqs_1_1_1 | in_arb_reqs_1_1_2 | in_arb_reqs_1_1_3) | in_arb_reqs_1_2_0; // @[package.scala 73:59]
  wire  in_arb_vals_1 = io_req_1_valid & _in_arb_vals_1_T_7; // @[SingleVCAllocator.scala 32:39]
  wire  in_arb_reqs_0_0_0 = io_req_0_bits_vc_sel_0_0 & ~io_channel_status_0_0_occupied; // @[SingleVCAllocator.scala 28:61]
  wire  in_arb_reqs_0_0_1 = io_req_0_bits_vc_sel_0_1 & ~io_channel_status_0_1_occupied; // @[SingleVCAllocator.scala 28:61]
  wire  in_arb_reqs_0_0_2 = io_req_0_bits_vc_sel_0_2 & ~io_channel_status_0_2_occupied; // @[SingleVCAllocator.scala 28:61]
  wire  in_arb_reqs_0_0_3 = io_req_0_bits_vc_sel_0_3 & ~io_channel_status_0_3_occupied; // @[SingleVCAllocator.scala 28:61]
  wire  in_arb_reqs_0_1_0 = io_req_0_bits_vc_sel_1_0 & ~io_channel_status_1_0_occupied; // @[SingleVCAllocator.scala 28:61]
  wire  in_arb_reqs_0_1_1 = io_req_0_bits_vc_sel_1_1 & ~io_channel_status_1_1_occupied; // @[SingleVCAllocator.scala 28:61]
  wire  in_arb_reqs_0_1_2 = io_req_0_bits_vc_sel_1_2 & ~io_channel_status_1_2_occupied; // @[SingleVCAllocator.scala 28:61]
  wire  in_arb_reqs_0_1_3 = io_req_0_bits_vc_sel_1_3 & ~io_channel_status_1_3_occupied; // @[SingleVCAllocator.scala 28:61]
  wire  in_arb_reqs_0_2_0 = io_req_0_bits_vc_sel_2_0 & ~io_channel_status_2_0_occupied; // @[SingleVCAllocator.scala 28:61]
  wire  _in_arb_vals_0_T_7 = in_arb_reqs_0_0_0 | in_arb_reqs_0_0_1 | in_arb_reqs_0_0_2 | in_arb_reqs_0_0_3 | (
    in_arb_reqs_0_1_0 | in_arb_reqs_0_1_1 | in_arb_reqs_0_1_2 | in_arb_reqs_0_1_3) | in_arb_reqs_0_2_0; // @[package.scala 73:59]
  wire  in_arb_vals_0 = io_req_0_valid & _in_arb_vals_0_T_7; // @[SingleVCAllocator.scala 32:39]
  wire [2:0] _in_arb_filter_T = {in_arb_vals_2,in_arb_vals_1,in_arb_vals_0}; // @[SingleVCAllocator.scala 19:57]
  wire [2:0] _in_arb_filter_T_2 = ~mask; // @[SingleVCAllocator.scala 19:86]
  wire [2:0] _in_arb_filter_T_3 = _in_arb_filter_T & _in_arb_filter_T_2; // @[SingleVCAllocator.scala 19:84]
  wire [5:0] _in_arb_filter_T_4 = {in_arb_vals_2,in_arb_vals_1,in_arb_vals_0,_in_arb_filter_T_3}; // @[Cat.scala 33:92]
  wire [5:0] _in_arb_filter_T_11 = _in_arb_filter_T_4[5] ? 6'h20 : 6'h0; // @[Mux.scala 47:70]
  wire [5:0] _in_arb_filter_T_12 = _in_arb_filter_T_4[4] ? 6'h10 : _in_arb_filter_T_11; // @[Mux.scala 47:70]
  wire [5:0] _in_arb_filter_T_13 = _in_arb_filter_T_4[3] ? 6'h8 : _in_arb_filter_T_12; // @[Mux.scala 47:70]
  wire [5:0] _in_arb_filter_T_14 = _in_arb_filter_T_4[2] ? 6'h4 : _in_arb_filter_T_13; // @[Mux.scala 47:70]
  wire [5:0] _in_arb_filter_T_15 = _in_arb_filter_T_4[1] ? 6'h2 : _in_arb_filter_T_14; // @[Mux.scala 47:70]
  wire [5:0] in_arb_filter = _in_arb_filter_T_4[0] ? 6'h1 : _in_arb_filter_T_15; // @[Mux.scala 47:70]
  wire [2:0] in_arb_sel = in_arb_filter[2:0] | in_arb_filter[5:3]; // @[SingleVCAllocator.scala 20:57]
  wire  _T_1 = in_arb_vals_0 | in_arb_vals_1 | in_arb_vals_2; // @[package.scala 73:59]
  wire [1:0] _mask_T_7 = in_arb_sel[1] ? 2'h3 : 2'h0; // @[Mux.scala 27:73]
  wire [2:0] _mask_T_8 = in_arb_sel[2] ? 3'h7 : 3'h0; // @[Mux.scala 27:73]
  wire [1:0] _GEN_2 = {{1'd0}, in_arb_sel[0]}; // @[Mux.scala 27:73]
  wire [1:0] _mask_T_9 = _GEN_2 | _mask_T_7; // @[Mux.scala 27:73]
  wire [2:0] _GEN_3 = {{1'd0}, _mask_T_9}; // @[Mux.scala 27:73]
  wire [2:0] _mask_T_10 = _GEN_3 | _mask_T_8; // @[Mux.scala 27:73]
  wire  in_vc_sel_0_0 = in_arb_sel[0] & in_arb_reqs_0_0_0 | in_arb_sel[1] & in_arb_reqs_1_0_0 | in_arb_sel[2] &
    in_arb_reqs_2_0_0; // @[Mux.scala 27:73]
  wire  in_vc_sel_0_1 = in_arb_sel[0] & in_arb_reqs_0_0_1 | in_arb_sel[1] & in_arb_reqs_1_0_1 | in_arb_sel[2] &
    in_arb_reqs_2_0_1; // @[Mux.scala 27:73]
  wire  in_vc_sel_0_2 = in_arb_sel[0] & in_arb_reqs_0_0_2 | in_arb_sel[1] & in_arb_reqs_1_0_2 | in_arb_sel[2] &
    in_arb_reqs_2_0_2; // @[Mux.scala 27:73]
  wire  in_vc_sel_0_3 = in_arb_sel[0] & in_arb_reqs_0_0_3 | in_arb_sel[1] & in_arb_reqs_1_0_3 | in_arb_sel[2] &
    in_arb_reqs_2_0_3; // @[Mux.scala 27:73]
  wire  in_vc_sel_1_0 = in_arb_sel[0] & in_arb_reqs_0_1_0 | in_arb_sel[1] & in_arb_reqs_1_1_0 | in_arb_sel[2] &
    in_arb_reqs_2_1_0; // @[Mux.scala 27:73]
  wire  in_vc_sel_1_1 = in_arb_sel[0] & in_arb_reqs_0_1_1 | in_arb_sel[1] & in_arb_reqs_1_1_1 | in_arb_sel[2] &
    in_arb_reqs_2_1_1; // @[Mux.scala 27:73]
  wire  in_vc_sel_1_2 = in_arb_sel[0] & in_arb_reqs_0_1_2 | in_arb_sel[1] & in_arb_reqs_1_1_2 | in_arb_sel[2] &
    in_arb_reqs_2_1_2; // @[Mux.scala 27:73]
  wire  in_vc_sel_1_3 = in_arb_sel[0] & in_arb_reqs_0_1_3 | in_arb_sel[1] & in_arb_reqs_1_1_3 | in_arb_sel[2] &
    in_arb_reqs_2_1_3; // @[Mux.scala 27:73]
  wire  in_vc_sel_2_0 = in_arb_sel[0] & in_arb_reqs_0_2_0 | in_arb_sel[1] & in_arb_reqs_1_2_0 | in_arb_sel[2] &
    in_arb_reqs_2_2_0; // @[Mux.scala 27:73]
  wire  _in_alloc_T_6 = io_req_0_ready & io_req_0_valid; // @[Decoupled.scala 51:35]
  wire  _in_alloc_T_7 = io_req_1_ready & io_req_1_valid; // @[Decoupled.scala 51:35]
  wire  _in_alloc_T_8 = io_req_2_ready & io_req_2_valid; // @[Decoupled.scala 51:35]
  wire  _in_alloc_T_10 = _in_alloc_T_6 | _in_alloc_T_7 | _in_alloc_T_8; // @[package.scala 73:59]
  wire [8:0] _in_alloc_T_11 = {in_vc_sel_2_0,in_vc_sel_1_3,in_vc_sel_1_2,in_vc_sel_1_1,in_vc_sel_1_0,in_vc_sel_0_3,
    in_vc_sel_0_2,in_vc_sel_0_1,in_vc_sel_0_0}; // @[ISLIP.scala 33:18]
  reg [8:0] in_alloc_mask; // @[ISLIP.scala 17:25]
  wire [8:0] _in_alloc_full_T = ~in_alloc_mask; // @[ISLIP.scala 18:31]
  wire [8:0] _in_alloc_full_T_1 = _in_alloc_T_11 & _in_alloc_full_T; // @[ISLIP.scala 18:29]
  wire [17:0] in_alloc_full = {in_vc_sel_2_0,in_vc_sel_1_3,in_vc_sel_1_2,in_vc_sel_1_1,in_vc_sel_1_0,in_vc_sel_0_3,
    in_vc_sel_0_2,in_vc_sel_0_1,in_vc_sel_0_0,_in_alloc_full_T_1}; // @[Cat.scala 33:92]
  wire [17:0] _in_alloc_oh_T_18 = in_alloc_full[17] ? 18'h20000 : 18'h0; // @[Mux.scala 47:70]
  wire [17:0] _in_alloc_oh_T_19 = in_alloc_full[16] ? 18'h10000 : _in_alloc_oh_T_18; // @[Mux.scala 47:70]
  wire [17:0] _in_alloc_oh_T_20 = in_alloc_full[15] ? 18'h8000 : _in_alloc_oh_T_19; // @[Mux.scala 47:70]
  wire [17:0] _in_alloc_oh_T_21 = in_alloc_full[14] ? 18'h4000 : _in_alloc_oh_T_20; // @[Mux.scala 47:70]
  wire [17:0] _in_alloc_oh_T_22 = in_alloc_full[13] ? 18'h2000 : _in_alloc_oh_T_21; // @[Mux.scala 47:70]
  wire [17:0] _in_alloc_oh_T_23 = in_alloc_full[12] ? 18'h1000 : _in_alloc_oh_T_22; // @[Mux.scala 47:70]
  wire [17:0] _in_alloc_oh_T_24 = in_alloc_full[11] ? 18'h800 : _in_alloc_oh_T_23; // @[Mux.scala 47:70]
  wire [17:0] _in_alloc_oh_T_25 = in_alloc_full[10] ? 18'h400 : _in_alloc_oh_T_24; // @[Mux.scala 47:70]
  wire [17:0] _in_alloc_oh_T_26 = in_alloc_full[9] ? 18'h200 : _in_alloc_oh_T_25; // @[Mux.scala 47:70]
  wire [17:0] _in_alloc_oh_T_27 = in_alloc_full[8] ? 18'h100 : _in_alloc_oh_T_26; // @[Mux.scala 47:70]
  wire [17:0] _in_alloc_oh_T_28 = in_alloc_full[7] ? 18'h80 : _in_alloc_oh_T_27; // @[Mux.scala 47:70]
  wire [17:0] _in_alloc_oh_T_29 = in_alloc_full[6] ? 18'h40 : _in_alloc_oh_T_28; // @[Mux.scala 47:70]
  wire [17:0] _in_alloc_oh_T_30 = in_alloc_full[5] ? 18'h20 : _in_alloc_oh_T_29; // @[Mux.scala 47:70]
  wire [17:0] _in_alloc_oh_T_31 = in_alloc_full[4] ? 18'h10 : _in_alloc_oh_T_30; // @[Mux.scala 47:70]
  wire [17:0] _in_alloc_oh_T_32 = in_alloc_full[3] ? 18'h8 : _in_alloc_oh_T_31; // @[Mux.scala 47:70]
  wire [17:0] _in_alloc_oh_T_33 = in_alloc_full[2] ? 18'h4 : _in_alloc_oh_T_32; // @[Mux.scala 47:70]
  wire [17:0] _in_alloc_oh_T_34 = in_alloc_full[1] ? 18'h2 : _in_alloc_oh_T_33; // @[Mux.scala 47:70]
  wire [17:0] in_alloc_oh = in_alloc_full[0] ? 18'h1 : _in_alloc_oh_T_34; // @[Mux.scala 47:70]
  wire [8:0] in_alloc_sel = in_alloc_oh[8:0] | in_alloc_oh[17:9]; // @[ISLIP.scala 20:28]
  wire [8:0] _in_alloc_mask_T_18 = in_alloc_sel[8] ? 9'h1ff : 9'h0; // @[Mux.scala 101:16]
  wire [8:0] _in_alloc_mask_T_19 = in_alloc_sel[7] ? 9'hff : _in_alloc_mask_T_18; // @[Mux.scala 101:16]
  wire [8:0] _in_alloc_mask_T_20 = in_alloc_sel[6] ? 9'h7f : _in_alloc_mask_T_19; // @[Mux.scala 101:16]
  wire [8:0] _in_alloc_mask_T_21 = in_alloc_sel[5] ? 9'h3f : _in_alloc_mask_T_20; // @[Mux.scala 101:16]
  wire [8:0] _in_alloc_mask_T_22 = in_alloc_sel[4] ? 9'h1f : _in_alloc_mask_T_21; // @[Mux.scala 101:16]
  wire [8:0] _in_alloc_mask_T_23 = in_alloc_sel[3] ? 9'hf : _in_alloc_mask_T_22; // @[Mux.scala 101:16]
  wire [8:0] _in_alloc_mask_T_24 = in_alloc_sel[2] ? 9'h7 : _in_alloc_mask_T_23; // @[Mux.scala 101:16]
  wire [8:0] _T_2 = {io_resp_0_vc_sel_2_0,io_resp_0_vc_sel_1_3,io_resp_0_vc_sel_1_2,io_resp_0_vc_sel_1_1,
    io_resp_0_vc_sel_1_0,io_resp_0_vc_sel_0_3,io_resp_0_vc_sel_0_2,io_resp_0_vc_sel_0_1,io_resp_0_vc_sel_0_0}; // @[SingleVCAllocator.scala 53:39]
  wire [1:0] _T_12 = _T_2[0] + _T_2[1]; // @[Bitwise.scala 51:90]
  wire [1:0] _T_14 = _T_2[2] + _T_2[3]; // @[Bitwise.scala 51:90]
  wire [2:0] _T_16 = _T_12 + _T_14; // @[Bitwise.scala 51:90]
  wire [1:0] _T_18 = _T_2[4] + _T_2[5]; // @[Bitwise.scala 51:90]
  wire [1:0] _T_20 = _T_2[7] + _T_2[8]; // @[Bitwise.scala 51:90]
  wire [1:0] _GEN_5 = {{1'd0}, _T_2[6]}; // @[Bitwise.scala 51:90]
  wire [2:0] _T_22 = _GEN_5 + _T_20; // @[Bitwise.scala 51:90]
  wire [2:0] _T_24 = _T_18 + _T_22[1:0]; // @[Bitwise.scala 51:90]
  wire [3:0] _T_26 = _T_16 + _T_24; // @[Bitwise.scala 51:90]
  wire [8:0] _T_32 = {io_resp_1_vc_sel_2_0,io_resp_1_vc_sel_1_3,io_resp_1_vc_sel_1_2,io_resp_1_vc_sel_1_1,
    io_resp_1_vc_sel_1_0,io_resp_1_vc_sel_0_3,io_resp_1_vc_sel_0_2,io_resp_1_vc_sel_0_1,io_resp_1_vc_sel_0_0}; // @[SingleVCAllocator.scala 53:39]
  wire [1:0] _T_42 = _T_32[0] + _T_32[1]; // @[Bitwise.scala 51:90]
  wire [1:0] _T_44 = _T_32[2] + _T_32[3]; // @[Bitwise.scala 51:90]
  wire [2:0] _T_46 = _T_42 + _T_44; // @[Bitwise.scala 51:90]
  wire [1:0] _T_48 = _T_32[4] + _T_32[5]; // @[Bitwise.scala 51:90]
  wire [1:0] _T_50 = _T_32[7] + _T_32[8]; // @[Bitwise.scala 51:90]
  wire [1:0] _GEN_6 = {{1'd0}, _T_32[6]}; // @[Bitwise.scala 51:90]
  wire [2:0] _T_52 = _GEN_6 + _T_50; // @[Bitwise.scala 51:90]
  wire [2:0] _T_54 = _T_48 + _T_52[1:0]; // @[Bitwise.scala 51:90]
  wire [3:0] _T_56 = _T_46 + _T_54; // @[Bitwise.scala 51:90]
  wire [8:0] _T_62 = {io_resp_2_vc_sel_2_0,io_resp_2_vc_sel_1_3,io_resp_2_vc_sel_1_2,io_resp_2_vc_sel_1_1,
    io_resp_2_vc_sel_1_0,io_resp_2_vc_sel_0_3,io_resp_2_vc_sel_0_2,io_resp_2_vc_sel_0_1,io_resp_2_vc_sel_0_0}; // @[SingleVCAllocator.scala 53:39]
  wire [1:0] _T_72 = _T_62[0] + _T_62[1]; // @[Bitwise.scala 51:90]
  wire [1:0] _T_74 = _T_62[2] + _T_62[3]; // @[Bitwise.scala 51:90]
  wire [2:0] _T_76 = _T_72 + _T_74; // @[Bitwise.scala 51:90]
  wire [1:0] _T_78 = _T_62[4] + _T_62[5]; // @[Bitwise.scala 51:90]
  wire [1:0] _T_80 = _T_62[7] + _T_62[8]; // @[Bitwise.scala 51:90]
  wire [1:0] _GEN_7 = {{1'd0}, _T_62[6]}; // @[Bitwise.scala 51:90]
  wire [2:0] _T_82 = _GEN_7 + _T_80; // @[Bitwise.scala 51:90]
  wire [2:0] _T_84 = _T_78 + _T_82[1:0]; // @[Bitwise.scala 51:90]
  wire [3:0] _T_86 = _T_76 + _T_84; // @[Bitwise.scala 51:90]
  assign io_req_2_ready = in_arb_sel[2]; // @[SingleVCAllocator.scala 47:34]
  assign io_req_1_ready = in_arb_sel[1]; // @[SingleVCAllocator.scala 47:34]
  assign io_req_0_ready = in_arb_sel[0]; // @[SingleVCAllocator.scala 47:34]
  assign io_resp_2_vc_sel_2_0 = _T_1 & in_alloc_sel[8]; // @[SingleVCAllocator.scala 41:18]
  assign io_resp_2_vc_sel_1_0 = _T_1 & in_alloc_sel[4]; // @[SingleVCAllocator.scala 41:18]
  assign io_resp_2_vc_sel_1_1 = _T_1 & in_alloc_sel[5]; // @[SingleVCAllocator.scala 41:18]
  assign io_resp_2_vc_sel_1_2 = _T_1 & in_alloc_sel[6]; // @[SingleVCAllocator.scala 41:18]
  assign io_resp_2_vc_sel_1_3 = _T_1 & in_alloc_sel[7]; // @[SingleVCAllocator.scala 41:18]
  assign io_resp_2_vc_sel_0_0 = _T_1 & in_alloc_sel[0]; // @[SingleVCAllocator.scala 41:18]
  assign io_resp_2_vc_sel_0_1 = _T_1 & in_alloc_sel[1]; // @[SingleVCAllocator.scala 41:18]
  assign io_resp_2_vc_sel_0_2 = _T_1 & in_alloc_sel[2]; // @[SingleVCAllocator.scala 41:18]
  assign io_resp_2_vc_sel_0_3 = _T_1 & in_alloc_sel[3]; // @[SingleVCAllocator.scala 41:18]
  assign io_resp_1_vc_sel_2_0 = _T_1 & in_alloc_sel[8]; // @[SingleVCAllocator.scala 41:18]
  assign io_resp_1_vc_sel_1_0 = _T_1 & in_alloc_sel[4]; // @[SingleVCAllocator.scala 41:18]
  assign io_resp_1_vc_sel_1_1 = _T_1 & in_alloc_sel[5]; // @[SingleVCAllocator.scala 41:18]
  assign io_resp_1_vc_sel_1_2 = _T_1 & in_alloc_sel[6]; // @[SingleVCAllocator.scala 41:18]
  assign io_resp_1_vc_sel_1_3 = _T_1 & in_alloc_sel[7]; // @[SingleVCAllocator.scala 41:18]
  assign io_resp_1_vc_sel_0_0 = _T_1 & in_alloc_sel[0]; // @[SingleVCAllocator.scala 41:18]
  assign io_resp_1_vc_sel_0_1 = _T_1 & in_alloc_sel[1]; // @[SingleVCAllocator.scala 41:18]
  assign io_resp_1_vc_sel_0_2 = _T_1 & in_alloc_sel[2]; // @[SingleVCAllocator.scala 41:18]
  assign io_resp_1_vc_sel_0_3 = _T_1 & in_alloc_sel[3]; // @[SingleVCAllocator.scala 41:18]
  assign io_resp_0_vc_sel_2_0 = _T_1 & in_alloc_sel[8]; // @[SingleVCAllocator.scala 41:18]
  assign io_resp_0_vc_sel_1_0 = _T_1 & in_alloc_sel[4]; // @[SingleVCAllocator.scala 41:18]
  assign io_resp_0_vc_sel_1_1 = _T_1 & in_alloc_sel[5]; // @[SingleVCAllocator.scala 41:18]
  assign io_resp_0_vc_sel_1_2 = _T_1 & in_alloc_sel[6]; // @[SingleVCAllocator.scala 41:18]
  assign io_resp_0_vc_sel_1_3 = _T_1 & in_alloc_sel[7]; // @[SingleVCAllocator.scala 41:18]
  assign io_resp_0_vc_sel_0_0 = _T_1 & in_alloc_sel[0]; // @[SingleVCAllocator.scala 41:18]
  assign io_resp_0_vc_sel_0_1 = _T_1 & in_alloc_sel[1]; // @[SingleVCAllocator.scala 41:18]
  assign io_resp_0_vc_sel_0_2 = _T_1 & in_alloc_sel[2]; // @[SingleVCAllocator.scala 41:18]
  assign io_resp_0_vc_sel_0_3 = _T_1 & in_alloc_sel[3]; // @[SingleVCAllocator.scala 41:18]
  assign io_out_allocs_2_0_alloc = _T_1 & in_alloc_sel[8]; // @[SingleVCAllocator.scala 41:18]
  assign io_out_allocs_1_0_alloc = _T_1 & in_alloc_sel[4]; // @[SingleVCAllocator.scala 41:18]
  assign io_out_allocs_1_1_alloc = _T_1 & in_alloc_sel[5]; // @[SingleVCAllocator.scala 41:18]
  assign io_out_allocs_1_2_alloc = _T_1 & in_alloc_sel[6]; // @[SingleVCAllocator.scala 41:18]
  assign io_out_allocs_1_3_alloc = _T_1 & in_alloc_sel[7]; // @[SingleVCAllocator.scala 41:18]
  assign io_out_allocs_0_0_alloc = _T_1 & in_alloc_sel[0]; // @[SingleVCAllocator.scala 41:18]
  assign io_out_allocs_0_1_alloc = _T_1 & in_alloc_sel[1]; // @[SingleVCAllocator.scala 41:18]
  assign io_out_allocs_0_2_alloc = _T_1 & in_alloc_sel[2]; // @[SingleVCAllocator.scala 41:18]
  assign io_out_allocs_0_3_alloc = _T_1 & in_alloc_sel[3]; // @[SingleVCAllocator.scala 41:18]
  always @(posedge clock) begin
    if (reset) begin // @[SingleVCAllocator.scala 16:21]
      mask <= 3'h0; // @[SingleVCAllocator.scala 16:21]
    end else if (_T_1) begin // @[SingleVCAllocator.scala 21:26]
      mask <= _mask_T_10; // @[SingleVCAllocator.scala 22:10]
    end
    if (reset) begin // @[ISLIP.scala 17:25]
      in_alloc_mask <= 9'h0; // @[ISLIP.scala 17:25]
    end else if (_in_alloc_T_10) begin // @[ISLIP.scala 21:19]
      if (in_alloc_sel[0]) begin // @[Mux.scala 101:16]
        in_alloc_mask <= 9'h1;
      end else if (in_alloc_sel[1]) begin // @[Mux.scala 101:16]
        in_alloc_mask <= 9'h3;
      end else begin
        in_alloc_mask <= _in_alloc_mask_T_24;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(_T_26 <= 4'h1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at SingleVCAllocator.scala:53 assert(PopCount(io.resp(i).vc_sel.asUInt) <= 1.U)\n"); // @[SingleVCAllocator.scala 53:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(_T_56 <= 4'h1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at SingleVCAllocator.scala:53 assert(PopCount(io.resp(i).vc_sel.asUInt) <= 1.U)\n"); // @[SingleVCAllocator.scala 53:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(_T_86 <= 4'h1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at SingleVCAllocator.scala:53 assert(PopCount(io.resp(i).vc_sel.asUInt) <= 1.U)\n"); // @[SingleVCAllocator.scala 53:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mask = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  in_alloc_mask = _RAND_1[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(_T_26 <= 4'h1); // @[SingleVCAllocator.scala 53:11]
    end
    //
    if (~reset) begin
      assert(_T_56 <= 4'h1); // @[SingleVCAllocator.scala 53:11]
    end
    //
    if (~reset) begin
      assert(_T_86 <= 4'h1); // @[SingleVCAllocator.scala 53:11]
    end
  end
endmodule
module RouteComputer(
  input  [1:0] io_req_2_bits_flow_ingress_node,
  input  [1:0] io_req_2_bits_flow_egress_node,
  input  [1:0] io_req_1_bits_src_virt_id,
  input  [1:0] io_req_1_bits_flow_ingress_node,
  input  [1:0] io_req_1_bits_flow_egress_node,
  input  [1:0] io_req_0_bits_src_virt_id,
  input  [1:0] io_req_0_bits_flow_ingress_node,
  input  [1:0] io_req_0_bits_flow_egress_node,
  output       io_resp_2_vc_sel_1_0,
  output       io_resp_2_vc_sel_1_1,
  output       io_resp_2_vc_sel_1_2,
  output       io_resp_2_vc_sel_1_3,
  output       io_resp_2_vc_sel_0_0,
  output       io_resp_2_vc_sel_0_1,
  output       io_resp_2_vc_sel_0_2,
  output       io_resp_2_vc_sel_0_3,
  output       io_resp_1_vc_sel_1_0,
  output       io_resp_1_vc_sel_1_1,
  output       io_resp_1_vc_sel_1_2,
  output       io_resp_1_vc_sel_0_0,
  output       io_resp_1_vc_sel_0_1,
  output       io_resp_1_vc_sel_0_2,
  output       io_resp_1_vc_sel_0_3,
  output       io_resp_0_vc_sel_1_0,
  output       io_resp_0_vc_sel_1_1,
  output       io_resp_0_vc_sel_1_2,
  output       io_resp_0_vc_sel_0_0,
  output       io_resp_0_vc_sel_0_1,
  output       io_resp_0_vc_sel_0_2,
  output       io_resp_0_vc_sel_0_3
);
  wire [5:0] addr = {io_req_0_bits_src_virt_id,io_req_0_bits_flow_ingress_node,io_req_0_bits_flow_egress_node}; // @[RouteComputer.scala 74:27]
  wire [5:0] decoded_invInputs = ~addr; // @[pla.scala 78:21]
  wire  decoded_andMatrixInput_0 = decoded_invInputs[0]; // @[pla.scala 91:29]
  wire  decoded_andMatrixInput_1 = decoded_invInputs[1]; // @[pla.scala 91:29]
  wire [1:0] _decoded_T = {decoded_andMatrixInput_0,decoded_andMatrixInput_1}; // @[Cat.scala 33:92]
  wire  _decoded_T_1 = &_decoded_T; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_0_1 = addr[0]; // @[pla.scala 90:45]
  wire  decoded_andMatrixInput_1_1 = addr[1]; // @[pla.scala 90:45]
  wire [1:0] _decoded_T_2 = {decoded_andMatrixInput_0_1,decoded_andMatrixInput_1_1}; // @[Cat.scala 33:92]
  wire  _decoded_T_3 = &_decoded_T_2; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_1_2 = addr[2]; // @[pla.scala 90:45]
  wire  decoded_andMatrixInput_2 = decoded_invInputs[3]; // @[pla.scala 91:29]
  wire  decoded_andMatrixInput_3 = decoded_invInputs[4]; // @[pla.scala 91:29]
  wire  decoded_andMatrixInput_4 = decoded_invInputs[5]; // @[pla.scala 91:29]
  wire [4:0] _decoded_T_4 = {decoded_andMatrixInput_1,decoded_andMatrixInput_1_2,decoded_andMatrixInput_2,
    decoded_andMatrixInput_3,decoded_andMatrixInput_4}; // @[Cat.scala 33:92]
  wire  _decoded_T_5 = &_decoded_T_4; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_0_3 = addr[3]; // @[pla.scala 90:45]
  wire [2:0] _decoded_T_6 = {decoded_andMatrixInput_0_3,decoded_andMatrixInput_3,decoded_andMatrixInput_4}; // @[Cat.scala 33:92]
  wire  _decoded_T_7 = &_decoded_T_6; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_1_4 = addr[4]; // @[pla.scala 90:45]
  wire [1:0] _decoded_T_8 = {decoded_andMatrixInput_0,decoded_andMatrixInput_1_4}; // @[Cat.scala 33:92]
  wire  _decoded_T_9 = &_decoded_T_8; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_1_5 = addr[5]; // @[pla.scala 90:45]
  wire [1:0] _decoded_T_10 = {decoded_andMatrixInput_0,decoded_andMatrixInput_1_5}; // @[Cat.scala 33:92]
  wire  _decoded_T_11 = &_decoded_T_10; // @[pla.scala 98:74]
  wire [1:0] _decoded_T_12 = {decoded_andMatrixInput_1_2,decoded_andMatrixInput_1_5}; // @[Cat.scala 33:92]
  wire  _decoded_T_13 = &_decoded_T_12; // @[pla.scala 98:74]
  wire [1:0] _decoded_T_14 = {decoded_andMatrixInput_1_4,decoded_andMatrixInput_1_5}; // @[Cat.scala 33:92]
  wire  _decoded_T_15 = &_decoded_T_14; // @[pla.scala 98:74]
  wire [4:0] _decoded_T_16 = {decoded_andMatrixInput_1,decoded_andMatrixInput_1_2,decoded_andMatrixInput_2,
    decoded_andMatrixInput_1_4,decoded_andMatrixInput_1_5}; // @[Cat.scala 33:92]
  wire  _decoded_T_17 = &_decoded_T_16; // @[pla.scala 98:74]
  wire [2:0] _decoded_T_18 = {decoded_andMatrixInput_0_3,decoded_andMatrixInput_1_4,decoded_andMatrixInput_1_5}; // @[Cat.scala 33:92]
  wire  _decoded_T_19 = &_decoded_T_18; // @[pla.scala 98:74]
  wire  _decoded_orMatrixOutputs_T = |_decoded_T_15; // @[pla.scala 114:39]
  wire [1:0] _decoded_orMatrixOutputs_T_1 = {_decoded_T_11,_decoded_T_13}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_2 = |_decoded_orMatrixOutputs_T_1; // @[pla.scala 114:39]
  wire [1:0] _decoded_orMatrixOutputs_T_3 = {_decoded_T_1,_decoded_T_3}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_4 = |_decoded_orMatrixOutputs_T_3; // @[pla.scala 114:39]
  wire [1:0] _decoded_orMatrixOutputs_T_5 = {_decoded_T_17,_decoded_T_19}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_6 = |_decoded_orMatrixOutputs_T_5; // @[pla.scala 114:39]
  wire  _decoded_orMatrixOutputs_T_7 = |_decoded_T_11; // @[pla.scala 114:39]
  wire [1:0] _decoded_orMatrixOutputs_T_8 = {_decoded_T_9,_decoded_T_11}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_9 = |_decoded_orMatrixOutputs_T_8; // @[pla.scala 114:39]
  wire [1:0] _decoded_orMatrixOutputs_T_10 = {_decoded_T_5,_decoded_T_7}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_11 = |_decoded_orMatrixOutputs_T_10; // @[pla.scala 114:39]
  wire [7:0] decoded_orMatrixOutputs = {_decoded_orMatrixOutputs_T_11,_decoded_orMatrixOutputs_T_9,
    _decoded_orMatrixOutputs_T_7,_decoded_orMatrixOutputs_T_6,_decoded_orMatrixOutputs_T_4,_decoded_orMatrixOutputs_T_2,
    _decoded_orMatrixOutputs_T,1'h0}; // @[Cat.scala 33:92]
  wire [7:0] decoded_invMatrixOutputs = {decoded_orMatrixOutputs[7],decoded_orMatrixOutputs[6],decoded_orMatrixOutputs[5
    ],decoded_orMatrixOutputs[4],decoded_orMatrixOutputs[3],decoded_orMatrixOutputs[2],decoded_orMatrixOutputs[1],
    decoded_orMatrixOutputs[0]}; // @[Cat.scala 33:92]
  wire [7:0] _GEN_0 = {{4'd0}, decoded_invMatrixOutputs[7:4]}; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_23 = _GEN_0 & 8'hf; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_25 = {decoded_invMatrixOutputs[3:0], 4'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _decoded_T_27 = _decoded_T_25 & 8'hf0; // @[Bitwise.scala 108:80]
  wire [7:0] _decoded_T_28 = _decoded_T_23 | _decoded_T_27; // @[Bitwise.scala 108:39]
  wire [7:0] _GEN_1 = {{2'd0}, _decoded_T_28[7:2]}; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_33 = _GEN_1 & 8'h33; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_35 = {_decoded_T_28[5:0], 2'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _decoded_T_37 = _decoded_T_35 & 8'hcc; // @[Bitwise.scala 108:80]
  wire [7:0] _decoded_T_38 = _decoded_T_33 | _decoded_T_37; // @[Bitwise.scala 108:39]
  wire [7:0] _GEN_2 = {{1'd0}, _decoded_T_38[7:1]}; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_43 = _GEN_2 & 8'h55; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_45 = {_decoded_T_38[6:0], 1'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _decoded_T_47 = _decoded_T_45 & 8'haa; // @[Bitwise.scala 108:80]
  wire [7:0] decoded = _decoded_T_43 | _decoded_T_47; // @[Bitwise.scala 108:39]
  wire [5:0] addr_1 = {io_req_1_bits_src_virt_id,io_req_1_bits_flow_ingress_node,io_req_1_bits_flow_egress_node}; // @[RouteComputer.scala 74:27]
  wire [5:0] decoded_invInputs_1 = ~addr_1; // @[pla.scala 78:21]
  wire  decoded_andMatrixInput_0_10 = decoded_invInputs_1[0]; // @[pla.scala 91:29]
  wire  decoded_andMatrixInput_1_10 = decoded_invInputs_1[1]; // @[pla.scala 91:29]
  wire [1:0] _decoded_T_48 = {decoded_andMatrixInput_0_10,decoded_andMatrixInput_1_10}; // @[Cat.scala 33:92]
  wire  _decoded_T_49 = &_decoded_T_48; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_0_11 = decoded_invInputs_1[4]; // @[pla.scala 91:29]
  wire  decoded_andMatrixInput_1_11 = decoded_invInputs_1[5]; // @[pla.scala 91:29]
  wire [1:0] _decoded_T_50 = {decoded_andMatrixInput_0_11,decoded_andMatrixInput_1_11}; // @[Cat.scala 33:92]
  wire  _decoded_T_51 = &_decoded_T_50; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_0_12 = addr_1[0]; // @[pla.scala 90:45]
  wire [1:0] _decoded_T_52 = {decoded_andMatrixInput_0_12,decoded_andMatrixInput_1_10}; // @[Cat.scala 33:92]
  wire  _decoded_T_53 = &_decoded_T_52; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_1_13 = addr_1[4]; // @[pla.scala 90:45]
  wire [1:0] _decoded_T_54 = {decoded_andMatrixInput_1_10,decoded_andMatrixInput_1_13}; // @[Cat.scala 33:92]
  wire  _decoded_T_55 = &_decoded_T_54; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_1_14 = addr_1[5]; // @[pla.scala 90:45]
  wire [1:0] _decoded_T_56 = {decoded_andMatrixInput_1_10,decoded_andMatrixInput_1_14}; // @[Cat.scala 33:92]
  wire  _decoded_T_57 = &_decoded_T_56; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_2_4 = addr_1[3]; // @[pla.scala 90:45]
  wire [3:0] _decoded_T_58 = {decoded_andMatrixInput_0_10,decoded_andMatrixInput_1_10,decoded_andMatrixInput_2_4,
    decoded_andMatrixInput_1_14}; // @[Cat.scala 33:92]
  wire  _decoded_T_59 = &_decoded_T_58; // @[pla.scala 98:74]
  wire [1:0] _decoded_T_60 = {decoded_andMatrixInput_1_13,decoded_andMatrixInput_1_14}; // @[Cat.scala 33:92]
  wire  _decoded_T_61 = &_decoded_T_60; // @[pla.scala 98:74]
  wire [3:0] _decoded_T_62 = {decoded_andMatrixInput_0_10,decoded_andMatrixInput_2_4,decoded_andMatrixInput_1_13,
    decoded_andMatrixInput_1_14}; // @[Cat.scala 33:92]
  wire  _decoded_T_63 = &_decoded_T_62; // @[pla.scala 98:74]
  wire  _decoded_orMatrixOutputs_T_12 = |_decoded_T_63; // @[pla.scala 114:39]
  wire  _decoded_orMatrixOutputs_T_13 = |_decoded_T_59; // @[pla.scala 114:39]
  wire  _decoded_orMatrixOutputs_T_14 = |_decoded_T_49; // @[pla.scala 114:39]
  wire  _decoded_orMatrixOutputs_T_15 = |_decoded_T_61; // @[pla.scala 114:39]
  wire  _decoded_orMatrixOutputs_T_16 = |_decoded_T_57; // @[pla.scala 114:39]
  wire [1:0] _decoded_orMatrixOutputs_T_17 = {_decoded_T_55,_decoded_T_57}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_18 = |_decoded_orMatrixOutputs_T_17; // @[pla.scala 114:39]
  wire [1:0] _decoded_orMatrixOutputs_T_19 = {_decoded_T_51,_decoded_T_53}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_20 = |_decoded_orMatrixOutputs_T_19; // @[pla.scala 114:39]
  wire [7:0] decoded_orMatrixOutputs_1 = {_decoded_orMatrixOutputs_T_20,_decoded_orMatrixOutputs_T_18,
    _decoded_orMatrixOutputs_T_16,_decoded_orMatrixOutputs_T_15,_decoded_orMatrixOutputs_T_14,
    _decoded_orMatrixOutputs_T_13,_decoded_orMatrixOutputs_T_12,1'h0}; // @[Cat.scala 33:92]
  wire [7:0] decoded_invMatrixOutputs_1 = {decoded_orMatrixOutputs_1[7],decoded_orMatrixOutputs_1[6],
    decoded_orMatrixOutputs_1[5],decoded_orMatrixOutputs_1[4],decoded_orMatrixOutputs_1[3],decoded_orMatrixOutputs_1[2],
    decoded_orMatrixOutputs_1[1],decoded_orMatrixOutputs_1[0]}; // @[Cat.scala 33:92]
  wire [7:0] _GEN_3 = {{4'd0}, decoded_invMatrixOutputs_1[7:4]}; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_67 = _GEN_3 & 8'hf; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_69 = {decoded_invMatrixOutputs_1[3:0], 4'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _decoded_T_71 = _decoded_T_69 & 8'hf0; // @[Bitwise.scala 108:80]
  wire [7:0] _decoded_T_72 = _decoded_T_67 | _decoded_T_71; // @[Bitwise.scala 108:39]
  wire [7:0] _GEN_4 = {{2'd0}, _decoded_T_72[7:2]}; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_77 = _GEN_4 & 8'h33; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_79 = {_decoded_T_72[5:0], 2'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _decoded_T_81 = _decoded_T_79 & 8'hcc; // @[Bitwise.scala 108:80]
  wire [7:0] _decoded_T_82 = _decoded_T_77 | _decoded_T_81; // @[Bitwise.scala 108:39]
  wire [7:0] _GEN_5 = {{1'd0}, _decoded_T_82[7:1]}; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_87 = _GEN_5 & 8'h55; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_89 = {_decoded_T_82[6:0], 1'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _decoded_T_91 = _decoded_T_89 & 8'haa; // @[Bitwise.scala 108:80]
  wire [7:0] decoded_1 = _decoded_T_87 | _decoded_T_91; // @[Bitwise.scala 108:39]
  wire [5:0] addr_2 = {2'h0,io_req_2_bits_flow_ingress_node,io_req_2_bits_flow_egress_node}; // @[RouteComputer.scala 74:27]
  wire [5:0] decoded_invInputs_2 = ~addr_2; // @[pla.scala 78:21]
  wire  decoded_andMatrixInput_0_18 = decoded_invInputs_2[0]; // @[pla.scala 91:29]
  wire  decoded_andMatrixInput_1_18 = decoded_invInputs_2[2]; // @[pla.scala 91:29]
  wire  decoded_andMatrixInput_2_6 = decoded_invInputs_2[3]; // @[pla.scala 91:29]
  wire  decoded_andMatrixInput_3_4 = decoded_invInputs_2[4]; // @[pla.scala 91:29]
  wire  decoded_andMatrixInput_4_2 = decoded_invInputs_2[5]; // @[pla.scala 91:29]
  wire [4:0] _decoded_T_92 = {decoded_andMatrixInput_0_18,decoded_andMatrixInput_1_18,decoded_andMatrixInput_2_6,
    decoded_andMatrixInput_3_4,decoded_andMatrixInput_4_2}; // @[Cat.scala 33:92]
  wire  _decoded_T_93 = &_decoded_T_92; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_0_19 = decoded_invInputs_2[1]; // @[pla.scala 91:29]
  wire [4:0] _decoded_T_94 = {decoded_andMatrixInput_0_19,decoded_andMatrixInput_1_18,decoded_andMatrixInput_2_6,
    decoded_andMatrixInput_3_4,decoded_andMatrixInput_4_2}; // @[Cat.scala 33:92]
  wire  _decoded_T_95 = &_decoded_T_94; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_0_20 = addr_2[1]; // @[pla.scala 90:45]
  wire [4:0] _decoded_T_96 = {decoded_andMatrixInput_0_20,decoded_andMatrixInput_1_18,decoded_andMatrixInput_2_6,
    decoded_andMatrixInput_3_4,decoded_andMatrixInput_4_2}; // @[Cat.scala 33:92]
  wire  _decoded_T_97 = &_decoded_T_96; // @[pla.scala 98:74]
  wire [1:0] _decoded_orMatrixOutputs_T_21 = {_decoded_T_93,_decoded_T_97}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_22 = |_decoded_orMatrixOutputs_T_21; // @[pla.scala 114:39]
  wire [1:0] _decoded_orMatrixOutputs_T_27 = {_decoded_T_93,_decoded_T_95}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_28 = |_decoded_orMatrixOutputs_T_27; // @[pla.scala 114:39]
  wire [7:0] decoded_orMatrixOutputs_2 = {1'h0,_decoded_orMatrixOutputs_T_28,_decoded_orMatrixOutputs_T_28,
    _decoded_orMatrixOutputs_T_28,1'h0,_decoded_orMatrixOutputs_T_22,_decoded_orMatrixOutputs_T_22,
    _decoded_orMatrixOutputs_T_22}; // @[Cat.scala 33:92]
  wire [7:0] decoded_invMatrixOutputs_2 = {decoded_orMatrixOutputs_2[7],decoded_orMatrixOutputs_2[6],
    decoded_orMatrixOutputs_2[5],decoded_orMatrixOutputs_2[4],decoded_orMatrixOutputs_2[3],decoded_orMatrixOutputs_2[2],
    decoded_orMatrixOutputs_2[1],decoded_orMatrixOutputs_2[0]}; // @[Cat.scala 33:92]
  wire [7:0] _GEN_6 = {{4'd0}, decoded_invMatrixOutputs_2[7:4]}; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_101 = _GEN_6 & 8'hf; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_103 = {decoded_invMatrixOutputs_2[3:0], 4'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _decoded_T_105 = _decoded_T_103 & 8'hf0; // @[Bitwise.scala 108:80]
  wire [7:0] _decoded_T_106 = _decoded_T_101 | _decoded_T_105; // @[Bitwise.scala 108:39]
  wire [7:0] _GEN_7 = {{2'd0}, _decoded_T_106[7:2]}; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_111 = _GEN_7 & 8'h33; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_113 = {_decoded_T_106[5:0], 2'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _decoded_T_115 = _decoded_T_113 & 8'hcc; // @[Bitwise.scala 108:80]
  wire [7:0] _decoded_T_116 = _decoded_T_111 | _decoded_T_115; // @[Bitwise.scala 108:39]
  wire [7:0] _GEN_8 = {{1'd0}, _decoded_T_116[7:1]}; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_121 = _GEN_8 & 8'h55; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_123 = {_decoded_T_116[6:0], 1'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _decoded_T_125 = _decoded_T_123 & 8'haa; // @[Bitwise.scala 108:80]
  wire [7:0] decoded_2 = _decoded_T_121 | _decoded_T_125; // @[Bitwise.scala 108:39]
  assign io_resp_2_vc_sel_1_0 = decoded_2[4]; // @[RouteComputer.scala 90:46]
  assign io_resp_2_vc_sel_1_1 = decoded_2[5]; // @[RouteComputer.scala 90:46]
  assign io_resp_2_vc_sel_1_2 = decoded_2[6]; // @[RouteComputer.scala 90:46]
  assign io_resp_2_vc_sel_1_3 = decoded_2[7]; // @[RouteComputer.scala 90:46]
  assign io_resp_2_vc_sel_0_0 = decoded_2[0]; // @[RouteComputer.scala 90:46]
  assign io_resp_2_vc_sel_0_1 = decoded_2[1]; // @[RouteComputer.scala 90:46]
  assign io_resp_2_vc_sel_0_2 = decoded_2[2]; // @[RouteComputer.scala 90:46]
  assign io_resp_2_vc_sel_0_3 = decoded_2[3]; // @[RouteComputer.scala 90:46]
  assign io_resp_1_vc_sel_1_0 = decoded_1[4]; // @[RouteComputer.scala 90:46]
  assign io_resp_1_vc_sel_1_1 = decoded_1[5]; // @[RouteComputer.scala 90:46]
  assign io_resp_1_vc_sel_1_2 = decoded_1[6]; // @[RouteComputer.scala 90:46]
  assign io_resp_1_vc_sel_0_0 = decoded_1[0]; // @[RouteComputer.scala 90:46]
  assign io_resp_1_vc_sel_0_1 = decoded_1[1]; // @[RouteComputer.scala 90:46]
  assign io_resp_1_vc_sel_0_2 = decoded_1[2]; // @[RouteComputer.scala 90:46]
  assign io_resp_1_vc_sel_0_3 = decoded_1[3]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_1_0 = decoded[4]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_1_1 = decoded[5]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_1_2 = decoded[6]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_0_0 = decoded[0]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_0_1 = decoded[1]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_0_2 = decoded[2]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_0_3 = decoded[3]; // @[RouteComputer.scala 90:46]
endmodule
module Router(
  input         clock,
  input         reset,
  output [1:0]  auto_debug_out_va_stall_0,
  output [1:0]  auto_debug_out_va_stall_1,
  output [1:0]  auto_debug_out_sa_stall_0,
  output [1:0]  auto_debug_out_sa_stall_1,
  output        auto_egress_nodes_out_flit_valid,
  output        auto_egress_nodes_out_flit_bits_head,
  output        auto_egress_nodes_out_flit_bits_tail,
  output [63:0] auto_egress_nodes_out_flit_bits_payload,
  output [1:0]  auto_egress_nodes_out_flit_bits_ingress_id,
  output        auto_ingress_nodes_in_flit_ready,
  input         auto_ingress_nodes_in_flit_valid,
  input         auto_ingress_nodes_in_flit_bits_head,
  input         auto_ingress_nodes_in_flit_bits_tail,
  input  [63:0] auto_ingress_nodes_in_flit_bits_payload,
  input  [1:0]  auto_ingress_nodes_in_flit_bits_egress_id,
  output        auto_source_nodes_out_1_flit_0_valid,
  output        auto_source_nodes_out_1_flit_0_bits_head,
  output        auto_source_nodes_out_1_flit_0_bits_tail,
  output [63:0] auto_source_nodes_out_1_flit_0_bits_payload,
  output [1:0]  auto_source_nodes_out_1_flit_0_bits_flow_ingress_node,
  output [1:0]  auto_source_nodes_out_1_flit_0_bits_flow_egress_node,
  output [1:0]  auto_source_nodes_out_1_flit_0_bits_virt_channel_id,
  input  [3:0]  auto_source_nodes_out_1_credit_return,
  input  [3:0]  auto_source_nodes_out_1_vc_free,
  output        auto_source_nodes_out_0_flit_0_valid,
  output        auto_source_nodes_out_0_flit_0_bits_head,
  output        auto_source_nodes_out_0_flit_0_bits_tail,
  output [63:0] auto_source_nodes_out_0_flit_0_bits_payload,
  output [1:0]  auto_source_nodes_out_0_flit_0_bits_flow_ingress_node,
  output [1:0]  auto_source_nodes_out_0_flit_0_bits_flow_egress_node,
  output [1:0]  auto_source_nodes_out_0_flit_0_bits_virt_channel_id,
  input  [3:0]  auto_source_nodes_out_0_credit_return,
  input  [3:0]  auto_source_nodes_out_0_vc_free,
  input         auto_dest_nodes_in_1_flit_0_valid,
  input         auto_dest_nodes_in_1_flit_0_bits_head,
  input         auto_dest_nodes_in_1_flit_0_bits_tail,
  input  [63:0] auto_dest_nodes_in_1_flit_0_bits_payload,
  input  [1:0]  auto_dest_nodes_in_1_flit_0_bits_flow_ingress_node,
  input  [1:0]  auto_dest_nodes_in_1_flit_0_bits_flow_egress_node,
  input  [1:0]  auto_dest_nodes_in_1_flit_0_bits_virt_channel_id,
  output [3:0]  auto_dest_nodes_in_1_credit_return,
  output [3:0]  auto_dest_nodes_in_1_vc_free,
  input         auto_dest_nodes_in_0_flit_0_valid,
  input         auto_dest_nodes_in_0_flit_0_bits_head,
  input         auto_dest_nodes_in_0_flit_0_bits_tail,
  input  [63:0] auto_dest_nodes_in_0_flit_0_bits_payload,
  input  [1:0]  auto_dest_nodes_in_0_flit_0_bits_flow_ingress_node,
  input  [1:0]  auto_dest_nodes_in_0_flit_0_bits_flow_egress_node,
  input  [1:0]  auto_dest_nodes_in_0_flit_0_bits_virt_channel_id,
  output [3:0]  auto_dest_nodes_in_0_credit_return,
  output [3:0]  auto_dest_nodes_in_0_vc_free
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_REG_INIT
  wire  monitor_clock; // @[Nodes.scala 24:25]
  wire  monitor_reset; // @[Nodes.scala 24:25]
  wire  monitor_io_in_flit_0_valid; // @[Nodes.scala 24:25]
  wire  monitor_io_in_flit_0_bits_head; // @[Nodes.scala 24:25]
  wire  monitor_io_in_flit_0_bits_tail; // @[Nodes.scala 24:25]
  wire [1:0] monitor_io_in_flit_0_bits_flow_ingress_node; // @[Nodes.scala 24:25]
  wire [1:0] monitor_io_in_flit_0_bits_flow_egress_node; // @[Nodes.scala 24:25]
  wire [1:0] monitor_io_in_flit_0_bits_virt_channel_id; // @[Nodes.scala 24:25]
  wire  monitor_1_clock; // @[Nodes.scala 24:25]
  wire  monitor_1_reset; // @[Nodes.scala 24:25]
  wire  monitor_1_io_in_flit_0_valid; // @[Nodes.scala 24:25]
  wire  monitor_1_io_in_flit_0_bits_head; // @[Nodes.scala 24:25]
  wire  monitor_1_io_in_flit_0_bits_tail; // @[Nodes.scala 24:25]
  wire [1:0] monitor_1_io_in_flit_0_bits_flow_ingress_node; // @[Nodes.scala 24:25]
  wire [1:0] monitor_1_io_in_flit_0_bits_flow_egress_node; // @[Nodes.scala 24:25]
  wire [1:0] monitor_1_io_in_flit_0_bits_virt_channel_id; // @[Nodes.scala 24:25]
  wire  input_unit_0_from_1_clock; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_reset; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_router_req_valid; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_1_io_router_req_bits_src_virt_id; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_1_io_router_req_bits_flow_ingress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_1_io_router_req_bits_flow_egress_node; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_router_resp_vc_sel_1_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_router_resp_vc_sel_1_1; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_router_resp_vc_sel_1_2; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_router_resp_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_router_resp_vc_sel_0_1; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_router_resp_vc_sel_0_2; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_router_resp_vc_sel_0_3; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_vcalloc_req_ready; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_vcalloc_req_valid; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_2_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_1_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_1_1; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_1_2; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_0_1; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_0_2; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_0_3; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_vcalloc_resp_vc_sel_2_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_vcalloc_resp_vc_sel_1_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_vcalloc_resp_vc_sel_1_1; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_vcalloc_resp_vc_sel_1_2; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_vcalloc_resp_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_vcalloc_resp_vc_sel_0_1; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_vcalloc_resp_vc_sel_0_2; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_vcalloc_resp_vc_sel_0_3; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_out_credit_available_2_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_out_credit_available_1_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_out_credit_available_1_1; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_out_credit_available_1_2; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_out_credit_available_1_3; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_out_credit_available_0_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_out_credit_available_0_1; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_out_credit_available_0_2; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_out_credit_available_0_3; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_salloc_req_0_ready; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_salloc_req_0_valid; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_2_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_1_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_1_1; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_1_2; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_1_3; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_0_1; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_0_2; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_0_3; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_salloc_req_0_bits_tail; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_out_0_valid; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_out_0_bits_flit_head; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_out_0_bits_flit_tail; // @[Router.scala 112:13]
  wire [63:0] input_unit_0_from_1_io_out_0_bits_flit_payload; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_1_io_out_0_bits_flit_flow_ingress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_1_io_out_0_bits_flit_flow_egress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_1_io_out_0_bits_out_virt_channel; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_1_io_debug_va_stall; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_1_io_debug_sa_stall; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_in_flit_0_valid; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_in_flit_0_bits_head; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_in_flit_0_bits_tail; // @[Router.scala 112:13]
  wire [63:0] input_unit_0_from_1_io_in_flit_0_bits_payload; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_1_io_in_flit_0_bits_flow_ingress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_1_io_in_flit_0_bits_flow_egress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_1_io_in_flit_0_bits_virt_channel_id; // @[Router.scala 112:13]
  wire [3:0] input_unit_0_from_1_io_in_credit_return; // @[Router.scala 112:13]
  wire [3:0] input_unit_0_from_1_io_in_vc_free; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_clock; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_reset; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_router_req_valid; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_3_io_router_req_bits_src_virt_id; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_3_io_router_req_bits_flow_ingress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_3_io_router_req_bits_flow_egress_node; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_router_resp_vc_sel_1_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_router_resp_vc_sel_1_1; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_router_resp_vc_sel_1_2; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_router_resp_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_router_resp_vc_sel_0_1; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_router_resp_vc_sel_0_2; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_router_resp_vc_sel_0_3; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_vcalloc_req_ready; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_vcalloc_req_valid; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_2_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_1_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_1_1; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_1_2; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_0_1; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_0_2; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_0_3; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_vcalloc_resp_vc_sel_2_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_vcalloc_resp_vc_sel_1_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_vcalloc_resp_vc_sel_1_1; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_vcalloc_resp_vc_sel_1_2; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_vcalloc_resp_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_vcalloc_resp_vc_sel_0_1; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_vcalloc_resp_vc_sel_0_2; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_vcalloc_resp_vc_sel_0_3; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_out_credit_available_2_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_out_credit_available_1_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_out_credit_available_1_1; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_out_credit_available_1_2; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_out_credit_available_1_3; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_out_credit_available_0_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_out_credit_available_0_1; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_out_credit_available_0_2; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_out_credit_available_0_3; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_salloc_req_0_ready; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_salloc_req_0_valid; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_2_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_1_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_1_1; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_1_2; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_1_3; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_0_1; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_0_2; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_0_3; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_salloc_req_0_bits_tail; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_out_0_valid; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_out_0_bits_flit_head; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_out_0_bits_flit_tail; // @[Router.scala 112:13]
  wire [63:0] input_unit_1_from_3_io_out_0_bits_flit_payload; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_3_io_out_0_bits_flit_flow_ingress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_3_io_out_0_bits_flit_flow_egress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_3_io_out_0_bits_out_virt_channel; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_3_io_debug_va_stall; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_3_io_debug_sa_stall; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_in_flit_0_valid; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_in_flit_0_bits_head; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_in_flit_0_bits_tail; // @[Router.scala 112:13]
  wire [63:0] input_unit_1_from_3_io_in_flit_0_bits_payload; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_3_io_in_flit_0_bits_flow_ingress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_3_io_in_flit_0_bits_flow_egress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_3_io_in_flit_0_bits_virt_channel_id; // @[Router.scala 112:13]
  wire [3:0] input_unit_1_from_3_io_in_credit_return; // @[Router.scala 112:13]
  wire [3:0] input_unit_1_from_3_io_in_vc_free; // @[Router.scala 112:13]
  wire  ingress_unit_2_from_0_clock; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_reset; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_router_req_valid; // @[Router.scala 116:13]
  wire [1:0] ingress_unit_2_from_0_io_router_req_bits_flow_ingress_node; // @[Router.scala 116:13]
  wire [1:0] ingress_unit_2_from_0_io_router_req_bits_flow_egress_node; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_router_resp_vc_sel_1_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_router_resp_vc_sel_1_1; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_router_resp_vc_sel_1_2; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_router_resp_vc_sel_1_3; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_router_resp_vc_sel_0_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_router_resp_vc_sel_0_1; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_router_resp_vc_sel_0_2; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_router_resp_vc_sel_0_3; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_vcalloc_req_ready; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_vcalloc_req_valid; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_vcalloc_req_bits_vc_sel_2_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_vcalloc_req_bits_vc_sel_1_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_vcalloc_req_bits_vc_sel_1_1; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_vcalloc_req_bits_vc_sel_1_2; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_vcalloc_req_bits_vc_sel_1_3; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_vcalloc_req_bits_vc_sel_0_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_vcalloc_req_bits_vc_sel_0_1; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_vcalloc_req_bits_vc_sel_0_2; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_vcalloc_req_bits_vc_sel_0_3; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_vcalloc_resp_vc_sel_2_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_vcalloc_resp_vc_sel_1_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_vcalloc_resp_vc_sel_1_1; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_vcalloc_resp_vc_sel_1_2; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_vcalloc_resp_vc_sel_1_3; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_vcalloc_resp_vc_sel_0_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_vcalloc_resp_vc_sel_0_1; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_vcalloc_resp_vc_sel_0_2; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_vcalloc_resp_vc_sel_0_3; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_out_credit_available_2_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_out_credit_available_1_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_out_credit_available_1_1; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_out_credit_available_1_2; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_out_credit_available_1_3; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_out_credit_available_0_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_out_credit_available_0_1; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_out_credit_available_0_2; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_out_credit_available_0_3; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_salloc_req_0_ready; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_salloc_req_0_valid; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_salloc_req_0_bits_vc_sel_2_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_salloc_req_0_bits_vc_sel_1_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_salloc_req_0_bits_vc_sel_1_1; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_salloc_req_0_bits_vc_sel_1_2; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_salloc_req_0_bits_vc_sel_1_3; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_salloc_req_0_bits_vc_sel_0_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_salloc_req_0_bits_vc_sel_0_1; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_salloc_req_0_bits_vc_sel_0_2; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_salloc_req_0_bits_vc_sel_0_3; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_salloc_req_0_bits_tail; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_out_0_valid; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_out_0_bits_flit_head; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_out_0_bits_flit_tail; // @[Router.scala 116:13]
  wire [63:0] ingress_unit_2_from_0_io_out_0_bits_flit_payload; // @[Router.scala 116:13]
  wire [1:0] ingress_unit_2_from_0_io_out_0_bits_flit_flow_ingress_node; // @[Router.scala 116:13]
  wire [1:0] ingress_unit_2_from_0_io_out_0_bits_flit_flow_egress_node; // @[Router.scala 116:13]
  wire [1:0] ingress_unit_2_from_0_io_out_0_bits_out_virt_channel; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_in_ready; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_in_valid; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_in_bits_head; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_0_io_in_bits_tail; // @[Router.scala 116:13]
  wire [63:0] ingress_unit_2_from_0_io_in_bits_payload; // @[Router.scala 116:13]
  wire [1:0] ingress_unit_2_from_0_io_in_bits_egress_id; // @[Router.scala 116:13]
  wire  output_unit_0_to_1_clock; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_reset; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_in_0_valid; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_in_0_bits_head; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_in_0_bits_tail; // @[Router.scala 122:13]
  wire [63:0] output_unit_0_to_1_io_in_0_bits_payload; // @[Router.scala 122:13]
  wire [1:0] output_unit_0_to_1_io_in_0_bits_flow_ingress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_0_to_1_io_in_0_bits_flow_egress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_0_to_1_io_in_0_bits_virt_channel_id; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_credit_available_0; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_credit_available_1; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_credit_available_2; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_credit_available_3; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_channel_status_0_occupied; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_channel_status_1_occupied; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_channel_status_2_occupied; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_channel_status_3_occupied; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_allocs_0_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_allocs_1_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_allocs_2_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_allocs_3_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_credit_alloc_0_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_credit_alloc_1_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_credit_alloc_2_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_credit_alloc_3_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_out_flit_0_valid; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_out_flit_0_bits_head; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_out_flit_0_bits_tail; // @[Router.scala 122:13]
  wire [63:0] output_unit_0_to_1_io_out_flit_0_bits_payload; // @[Router.scala 122:13]
  wire [1:0] output_unit_0_to_1_io_out_flit_0_bits_flow_ingress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_0_to_1_io_out_flit_0_bits_flow_egress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_0_to_1_io_out_flit_0_bits_virt_channel_id; // @[Router.scala 122:13]
  wire [3:0] output_unit_0_to_1_io_out_credit_return; // @[Router.scala 122:13]
  wire [3:0] output_unit_0_to_1_io_out_vc_free; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_clock; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_reset; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_in_0_valid; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_in_0_bits_head; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_in_0_bits_tail; // @[Router.scala 122:13]
  wire [63:0] output_unit_1_to_3_io_in_0_bits_payload; // @[Router.scala 122:13]
  wire [1:0] output_unit_1_to_3_io_in_0_bits_flow_ingress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_1_to_3_io_in_0_bits_flow_egress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_1_to_3_io_in_0_bits_virt_channel_id; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_credit_available_0; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_credit_available_1; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_credit_available_2; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_credit_available_3; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_channel_status_0_occupied; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_channel_status_1_occupied; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_channel_status_2_occupied; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_channel_status_3_occupied; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_allocs_0_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_allocs_1_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_allocs_2_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_allocs_3_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_credit_alloc_0_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_credit_alloc_1_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_credit_alloc_2_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_credit_alloc_3_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_out_flit_0_valid; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_out_flit_0_bits_head; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_out_flit_0_bits_tail; // @[Router.scala 122:13]
  wire [63:0] output_unit_1_to_3_io_out_flit_0_bits_payload; // @[Router.scala 122:13]
  wire [1:0] output_unit_1_to_3_io_out_flit_0_bits_flow_ingress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_1_to_3_io_out_flit_0_bits_flow_egress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_1_to_3_io_out_flit_0_bits_virt_channel_id; // @[Router.scala 122:13]
  wire [3:0] output_unit_1_to_3_io_out_credit_return; // @[Router.scala 122:13]
  wire [3:0] output_unit_1_to_3_io_out_vc_free; // @[Router.scala 122:13]
  wire  egress_unit_2_to_0_clock; // @[Router.scala 125:13]
  wire  egress_unit_2_to_0_reset; // @[Router.scala 125:13]
  wire  egress_unit_2_to_0_io_in_0_valid; // @[Router.scala 125:13]
  wire  egress_unit_2_to_0_io_in_0_bits_head; // @[Router.scala 125:13]
  wire  egress_unit_2_to_0_io_in_0_bits_tail; // @[Router.scala 125:13]
  wire [63:0] egress_unit_2_to_0_io_in_0_bits_payload; // @[Router.scala 125:13]
  wire [1:0] egress_unit_2_to_0_io_in_0_bits_flow_ingress_node; // @[Router.scala 125:13]
  wire  egress_unit_2_to_0_io_credit_available_0; // @[Router.scala 125:13]
  wire  egress_unit_2_to_0_io_channel_status_0_occupied; // @[Router.scala 125:13]
  wire  egress_unit_2_to_0_io_allocs_0_alloc; // @[Router.scala 125:13]
  wire  egress_unit_2_to_0_io_credit_alloc_0_alloc; // @[Router.scala 125:13]
  wire  egress_unit_2_to_0_io_credit_alloc_0_tail; // @[Router.scala 125:13]
  wire  egress_unit_2_to_0_io_out_valid; // @[Router.scala 125:13]
  wire  egress_unit_2_to_0_io_out_bits_head; // @[Router.scala 125:13]
  wire  egress_unit_2_to_0_io_out_bits_tail; // @[Router.scala 125:13]
  wire [63:0] egress_unit_2_to_0_io_out_bits_payload; // @[Router.scala 125:13]
  wire [1:0] egress_unit_2_to_0_io_out_bits_ingress_id; // @[Router.scala 125:13]
  wire  switch_clock; // @[Router.scala 129:24]
  wire  switch_reset; // @[Router.scala 129:24]
  wire  switch_io_in_2_0_valid; // @[Router.scala 129:24]
  wire  switch_io_in_2_0_bits_flit_head; // @[Router.scala 129:24]
  wire  switch_io_in_2_0_bits_flit_tail; // @[Router.scala 129:24]
  wire [63:0] switch_io_in_2_0_bits_flit_payload; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_2_0_bits_flit_flow_ingress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_2_0_bits_flit_flow_egress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_2_0_bits_out_virt_channel; // @[Router.scala 129:24]
  wire  switch_io_in_1_0_valid; // @[Router.scala 129:24]
  wire  switch_io_in_1_0_bits_flit_head; // @[Router.scala 129:24]
  wire  switch_io_in_1_0_bits_flit_tail; // @[Router.scala 129:24]
  wire [63:0] switch_io_in_1_0_bits_flit_payload; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_1_0_bits_flit_flow_ingress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_1_0_bits_flit_flow_egress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_1_0_bits_out_virt_channel; // @[Router.scala 129:24]
  wire  switch_io_in_0_0_valid; // @[Router.scala 129:24]
  wire  switch_io_in_0_0_bits_flit_head; // @[Router.scala 129:24]
  wire  switch_io_in_0_0_bits_flit_tail; // @[Router.scala 129:24]
  wire [63:0] switch_io_in_0_0_bits_flit_payload; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_0_0_bits_flit_flow_ingress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_0_0_bits_flit_flow_egress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_0_0_bits_out_virt_channel; // @[Router.scala 129:24]
  wire  switch_io_out_2_0_valid; // @[Router.scala 129:24]
  wire  switch_io_out_2_0_bits_head; // @[Router.scala 129:24]
  wire  switch_io_out_2_0_bits_tail; // @[Router.scala 129:24]
  wire [63:0] switch_io_out_2_0_bits_payload; // @[Router.scala 129:24]
  wire [1:0] switch_io_out_2_0_bits_flow_ingress_node; // @[Router.scala 129:24]
  wire  switch_io_out_1_0_valid; // @[Router.scala 129:24]
  wire  switch_io_out_1_0_bits_head; // @[Router.scala 129:24]
  wire  switch_io_out_1_0_bits_tail; // @[Router.scala 129:24]
  wire [63:0] switch_io_out_1_0_bits_payload; // @[Router.scala 129:24]
  wire [1:0] switch_io_out_1_0_bits_flow_ingress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_out_1_0_bits_flow_egress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_out_1_0_bits_virt_channel_id; // @[Router.scala 129:24]
  wire  switch_io_out_0_0_valid; // @[Router.scala 129:24]
  wire  switch_io_out_0_0_bits_head; // @[Router.scala 129:24]
  wire  switch_io_out_0_0_bits_tail; // @[Router.scala 129:24]
  wire [63:0] switch_io_out_0_0_bits_payload; // @[Router.scala 129:24]
  wire [1:0] switch_io_out_0_0_bits_flow_ingress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_out_0_0_bits_flow_egress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_out_0_0_bits_virt_channel_id; // @[Router.scala 129:24]
  wire  switch_io_sel_2_0_2_0; // @[Router.scala 129:24]
  wire  switch_io_sel_2_0_1_0; // @[Router.scala 129:24]
  wire  switch_io_sel_2_0_0_0; // @[Router.scala 129:24]
  wire  switch_io_sel_1_0_2_0; // @[Router.scala 129:24]
  wire  switch_io_sel_1_0_1_0; // @[Router.scala 129:24]
  wire  switch_io_sel_1_0_0_0; // @[Router.scala 129:24]
  wire  switch_io_sel_0_0_2_0; // @[Router.scala 129:24]
  wire  switch_io_sel_0_0_1_0; // @[Router.scala 129:24]
  wire  switch_io_sel_0_0_0_0; // @[Router.scala 129:24]
  wire  switch_allocator_clock; // @[Router.scala 130:34]
  wire  switch_allocator_reset; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_ready; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_valid; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_bits_vc_sel_2_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_bits_vc_sel_1_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_bits_vc_sel_1_1; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_bits_vc_sel_1_2; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_bits_vc_sel_1_3; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_bits_vc_sel_0_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_bits_vc_sel_0_1; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_bits_vc_sel_0_2; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_bits_vc_sel_0_3; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_bits_tail; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_ready; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_valid; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_vc_sel_2_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_vc_sel_1_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_vc_sel_1_1; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_vc_sel_1_2; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_vc_sel_1_3; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_vc_sel_0_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_vc_sel_0_1; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_vc_sel_0_2; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_vc_sel_0_3; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_tail; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_ready; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_valid; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_2_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_1_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_1_1; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_1_2; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_1_3; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_0_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_0_1; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_0_2; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_0_3; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_tail; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_2_0_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_2_0_tail; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_1_0_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_1_1_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_1_2_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_1_3_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_0_0_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_0_1_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_0_2_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_0_3_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_2_0_2_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_2_0_1_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_2_0_0_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_1_0_2_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_1_0_1_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_1_0_0_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_0_0_2_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_0_0_1_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_0_0_0_0; // @[Router.scala 130:34]
  wire  vc_allocator_clock; // @[Router.scala 131:30]
  wire  vc_allocator_reset; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_ready; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_valid; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_bits_vc_sel_2_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_bits_vc_sel_1_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_bits_vc_sel_1_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_bits_vc_sel_1_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_bits_vc_sel_1_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_bits_vc_sel_0_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_bits_vc_sel_0_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_bits_vc_sel_0_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_bits_vc_sel_0_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_ready; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_valid; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_bits_vc_sel_2_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_bits_vc_sel_1_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_bits_vc_sel_1_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_bits_vc_sel_1_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_bits_vc_sel_1_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_bits_vc_sel_0_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_bits_vc_sel_0_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_bits_vc_sel_0_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_bits_vc_sel_0_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_ready; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_valid; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_2_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_1_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_1_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_1_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_1_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_0_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_0_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_0_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_0_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_2_vc_sel_2_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_2_vc_sel_1_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_2_vc_sel_1_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_2_vc_sel_1_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_2_vc_sel_1_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_2_vc_sel_0_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_2_vc_sel_0_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_2_vc_sel_0_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_2_vc_sel_0_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_1_vc_sel_2_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_1_vc_sel_1_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_1_vc_sel_1_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_1_vc_sel_1_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_1_vc_sel_1_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_1_vc_sel_0_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_1_vc_sel_0_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_1_vc_sel_0_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_1_vc_sel_0_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_2_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_1_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_1_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_1_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_1_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_0_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_0_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_0_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_0_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_2_0_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_1_0_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_1_1_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_1_2_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_1_3_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_0_0_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_0_1_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_0_2_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_0_3_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_2_0_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_1_0_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_1_1_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_1_2_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_1_3_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_0_0_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_0_1_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_0_2_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_0_3_alloc; // @[Router.scala 131:30]
  wire [1:0] route_computer_io_req_2_bits_flow_ingress_node; // @[Router.scala 134:32]
  wire [1:0] route_computer_io_req_2_bits_flow_egress_node; // @[Router.scala 134:32]
  wire [1:0] route_computer_io_req_1_bits_src_virt_id; // @[Router.scala 134:32]
  wire [1:0] route_computer_io_req_1_bits_flow_ingress_node; // @[Router.scala 134:32]
  wire [1:0] route_computer_io_req_1_bits_flow_egress_node; // @[Router.scala 134:32]
  wire [1:0] route_computer_io_req_0_bits_src_virt_id; // @[Router.scala 134:32]
  wire [1:0] route_computer_io_req_0_bits_flow_ingress_node; // @[Router.scala 134:32]
  wire [1:0] route_computer_io_req_0_bits_flow_egress_node; // @[Router.scala 134:32]
  wire  route_computer_io_resp_2_vc_sel_1_0; // @[Router.scala 134:32]
  wire  route_computer_io_resp_2_vc_sel_1_1; // @[Router.scala 134:32]
  wire  route_computer_io_resp_2_vc_sel_1_2; // @[Router.scala 134:32]
  wire  route_computer_io_resp_2_vc_sel_1_3; // @[Router.scala 134:32]
  wire  route_computer_io_resp_2_vc_sel_0_0; // @[Router.scala 134:32]
  wire  route_computer_io_resp_2_vc_sel_0_1; // @[Router.scala 134:32]
  wire  route_computer_io_resp_2_vc_sel_0_2; // @[Router.scala 134:32]
  wire  route_computer_io_resp_2_vc_sel_0_3; // @[Router.scala 134:32]
  wire  route_computer_io_resp_1_vc_sel_1_0; // @[Router.scala 134:32]
  wire  route_computer_io_resp_1_vc_sel_1_1; // @[Router.scala 134:32]
  wire  route_computer_io_resp_1_vc_sel_1_2; // @[Router.scala 134:32]
  wire  route_computer_io_resp_1_vc_sel_0_0; // @[Router.scala 134:32]
  wire  route_computer_io_resp_1_vc_sel_0_1; // @[Router.scala 134:32]
  wire  route_computer_io_resp_1_vc_sel_0_2; // @[Router.scala 134:32]
  wire  route_computer_io_resp_1_vc_sel_0_3; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_1_0; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_1_1; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_1_2; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_0_0; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_0_1; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_0_2; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_0_3; // @[Router.scala 134:32]
  wire [19:0] plusarg_reader_out; // @[PlusArg.scala 80:11]
  wire  _fires_count_T = vc_allocator_io_req_0_ready & vc_allocator_io_req_0_valid; // @[Decoupled.scala 51:35]
  wire  _fires_count_T_1 = vc_allocator_io_req_1_ready & vc_allocator_io_req_1_valid; // @[Decoupled.scala 51:35]
  wire  _fires_count_T_2 = vc_allocator_io_req_2_ready & vc_allocator_io_req_2_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _fires_count_T_3 = _fires_count_T_1 + _fires_count_T_2; // @[Bitwise.scala 51:90]
  wire [1:0] _GEN_5 = {{1'd0}, _fires_count_T}; // @[Bitwise.scala 51:90]
  wire [2:0] _fires_count_T_5 = _GEN_5 + _fires_count_T_3; // @[Bitwise.scala 51:90]
  reg  switch_io_sel_REG_2_0_2_0; // @[Router.scala 176:14]
  reg  switch_io_sel_REG_2_0_1_0; // @[Router.scala 176:14]
  reg  switch_io_sel_REG_2_0_0_0; // @[Router.scala 176:14]
  reg  switch_io_sel_REG_1_0_2_0; // @[Router.scala 176:14]
  reg  switch_io_sel_REG_1_0_1_0; // @[Router.scala 176:14]
  reg  switch_io_sel_REG_1_0_0_0; // @[Router.scala 176:14]
  reg  switch_io_sel_REG_0_0_2_0; // @[Router.scala 176:14]
  reg  switch_io_sel_REG_0_0_1_0; // @[Router.scala 176:14]
  reg  switch_io_sel_REG_0_0_0_0; // @[Router.scala 176:14]
  reg [63:0] debug_tsc; // @[Router.scala 193:28]
  wire [63:0] _debug_tsc_T_1 = debug_tsc + 64'h1; // @[Router.scala 194:28]
  reg [63:0] debug_sample; // @[Router.scala 195:31]
  wire [63:0] _debug_sample_T_1 = debug_sample + 64'h1; // @[Router.scala 196:34]
  wire [19:0] _T_1 = plusarg_reader_out - 20'h1; // @[Router.scala 198:40]
  wire [63:0] _GEN_6 = {{44'd0}, _T_1}; // @[Router.scala 198:24]
  wire  _T_2 = debug_sample == _GEN_6; // @[Router.scala 198:24]
  reg [63:0] util_ctr; // @[Router.scala 201:29]
  reg  fired; // @[Router.scala 202:26]
  wire [63:0] _GEN_7 = {{63'd0}, auto_dest_nodes_in_0_flit_0_valid}; // @[Router.scala 203:28]
  wire [63:0] _util_ctr_T_1 = util_ctr + _GEN_7; // @[Router.scala 203:28]
  wire  _T_8 = plusarg_reader_out != 20'h0 & _T_2 & fired; // @[Router.scala 205:71]
  reg [63:0] util_ctr_1; // @[Router.scala 201:29]
  reg  fired_1; // @[Router.scala 202:26]
  wire [63:0] _GEN_9 = {{63'd0}, auto_dest_nodes_in_1_flit_0_valid}; // @[Router.scala 203:28]
  wire [63:0] _util_ctr_T_3 = util_ctr_1 + _GEN_9; // @[Router.scala 203:28]
  wire  _T_16 = plusarg_reader_out != 20'h0 & _T_2 & fired_1; // @[Router.scala 205:71]
  wire  bundleIn_0_2_flit_ready = ingress_unit_2_from_0_io_in_ready; // @[Nodes.scala 1215:84 Router.scala 142:68]
  wire  _T_19 = bundleIn_0_2_flit_ready & auto_ingress_nodes_in_flit_valid; // @[Decoupled.scala 51:35]
  reg [63:0] util_ctr_2; // @[Router.scala 201:29]
  reg  fired_2; // @[Router.scala 202:26]
  wire [63:0] _GEN_11 = {{63'd0}, _T_19}; // @[Router.scala 203:28]
  wire [63:0] _util_ctr_T_5 = util_ctr_2 + _GEN_11; // @[Router.scala 203:28]
  wire  _T_25 = plusarg_reader_out != 20'h0 & _T_2 & fired_2; // @[Router.scala 205:71]
  wire  x1_2_flit_valid = egress_unit_2_to_0_io_out_valid; // @[Nodes.scala 1212:84 Router.scala 144:65]
  reg [63:0] util_ctr_3; // @[Router.scala 201:29]
  reg  fired_3; // @[Router.scala 202:26]
  wire [63:0] _GEN_13 = {{63'd0}, x1_2_flit_valid}; // @[Router.scala 203:28]
  wire [63:0] _util_ctr_T_7 = util_ctr_3 + _GEN_13; // @[Router.scala 203:28]
  wire  _T_34 = plusarg_reader_out != 20'h0 & _T_2 & fired_3; // @[Router.scala 205:71]
  wire [1:0] fires_count = _fires_count_T_5[1:0]; // @[Bitwise.scala 51:90]
  NoCMonitor monitor ( // @[Nodes.scala 24:25]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_flit_0_valid(monitor_io_in_flit_0_valid),
    .io_in_flit_0_bits_head(monitor_io_in_flit_0_bits_head),
    .io_in_flit_0_bits_tail(monitor_io_in_flit_0_bits_tail),
    .io_in_flit_0_bits_flow_ingress_node(monitor_io_in_flit_0_bits_flow_ingress_node),
    .io_in_flit_0_bits_flow_egress_node(monitor_io_in_flit_0_bits_flow_egress_node),
    .io_in_flit_0_bits_virt_channel_id(monitor_io_in_flit_0_bits_virt_channel_id)
  );
  NoCMonitor_1 monitor_1 ( // @[Nodes.scala 24:25]
    .clock(monitor_1_clock),
    .reset(monitor_1_reset),
    .io_in_flit_0_valid(monitor_1_io_in_flit_0_valid),
    .io_in_flit_0_bits_head(monitor_1_io_in_flit_0_bits_head),
    .io_in_flit_0_bits_tail(monitor_1_io_in_flit_0_bits_tail),
    .io_in_flit_0_bits_flow_ingress_node(monitor_1_io_in_flit_0_bits_flow_ingress_node),
    .io_in_flit_0_bits_flow_egress_node(monitor_1_io_in_flit_0_bits_flow_egress_node),
    .io_in_flit_0_bits_virt_channel_id(monitor_1_io_in_flit_0_bits_virt_channel_id)
  );
  InputUnit input_unit_0_from_1 ( // @[Router.scala 112:13]
    .clock(input_unit_0_from_1_clock),
    .reset(input_unit_0_from_1_reset),
    .io_router_req_valid(input_unit_0_from_1_io_router_req_valid),
    .io_router_req_bits_src_virt_id(input_unit_0_from_1_io_router_req_bits_src_virt_id),
    .io_router_req_bits_flow_ingress_node(input_unit_0_from_1_io_router_req_bits_flow_ingress_node),
    .io_router_req_bits_flow_egress_node(input_unit_0_from_1_io_router_req_bits_flow_egress_node),
    .io_router_resp_vc_sel_1_0(input_unit_0_from_1_io_router_resp_vc_sel_1_0),
    .io_router_resp_vc_sel_1_1(input_unit_0_from_1_io_router_resp_vc_sel_1_1),
    .io_router_resp_vc_sel_1_2(input_unit_0_from_1_io_router_resp_vc_sel_1_2),
    .io_router_resp_vc_sel_0_0(input_unit_0_from_1_io_router_resp_vc_sel_0_0),
    .io_router_resp_vc_sel_0_1(input_unit_0_from_1_io_router_resp_vc_sel_0_1),
    .io_router_resp_vc_sel_0_2(input_unit_0_from_1_io_router_resp_vc_sel_0_2),
    .io_router_resp_vc_sel_0_3(input_unit_0_from_1_io_router_resp_vc_sel_0_3),
    .io_vcalloc_req_ready(input_unit_0_from_1_io_vcalloc_req_ready),
    .io_vcalloc_req_valid(input_unit_0_from_1_io_vcalloc_req_valid),
    .io_vcalloc_req_bits_vc_sel_2_0(input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_2_0),
    .io_vcalloc_req_bits_vc_sel_1_0(input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_1_0),
    .io_vcalloc_req_bits_vc_sel_1_1(input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_1_1),
    .io_vcalloc_req_bits_vc_sel_1_2(input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_1_2),
    .io_vcalloc_req_bits_vc_sel_0_0(input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_0_0),
    .io_vcalloc_req_bits_vc_sel_0_1(input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_0_1),
    .io_vcalloc_req_bits_vc_sel_0_2(input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_0_2),
    .io_vcalloc_req_bits_vc_sel_0_3(input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_0_3),
    .io_vcalloc_resp_vc_sel_2_0(input_unit_0_from_1_io_vcalloc_resp_vc_sel_2_0),
    .io_vcalloc_resp_vc_sel_1_0(input_unit_0_from_1_io_vcalloc_resp_vc_sel_1_0),
    .io_vcalloc_resp_vc_sel_1_1(input_unit_0_from_1_io_vcalloc_resp_vc_sel_1_1),
    .io_vcalloc_resp_vc_sel_1_2(input_unit_0_from_1_io_vcalloc_resp_vc_sel_1_2),
    .io_vcalloc_resp_vc_sel_0_0(input_unit_0_from_1_io_vcalloc_resp_vc_sel_0_0),
    .io_vcalloc_resp_vc_sel_0_1(input_unit_0_from_1_io_vcalloc_resp_vc_sel_0_1),
    .io_vcalloc_resp_vc_sel_0_2(input_unit_0_from_1_io_vcalloc_resp_vc_sel_0_2),
    .io_vcalloc_resp_vc_sel_0_3(input_unit_0_from_1_io_vcalloc_resp_vc_sel_0_3),
    .io_out_credit_available_2_0(input_unit_0_from_1_io_out_credit_available_2_0),
    .io_out_credit_available_1_0(input_unit_0_from_1_io_out_credit_available_1_0),
    .io_out_credit_available_1_1(input_unit_0_from_1_io_out_credit_available_1_1),
    .io_out_credit_available_1_2(input_unit_0_from_1_io_out_credit_available_1_2),
    .io_out_credit_available_1_3(input_unit_0_from_1_io_out_credit_available_1_3),
    .io_out_credit_available_0_0(input_unit_0_from_1_io_out_credit_available_0_0),
    .io_out_credit_available_0_1(input_unit_0_from_1_io_out_credit_available_0_1),
    .io_out_credit_available_0_2(input_unit_0_from_1_io_out_credit_available_0_2),
    .io_out_credit_available_0_3(input_unit_0_from_1_io_out_credit_available_0_3),
    .io_salloc_req_0_ready(input_unit_0_from_1_io_salloc_req_0_ready),
    .io_salloc_req_0_valid(input_unit_0_from_1_io_salloc_req_0_valid),
    .io_salloc_req_0_bits_vc_sel_2_0(input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_2_0),
    .io_salloc_req_0_bits_vc_sel_1_0(input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_1_0),
    .io_salloc_req_0_bits_vc_sel_1_1(input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_1_1),
    .io_salloc_req_0_bits_vc_sel_1_2(input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_1_2),
    .io_salloc_req_0_bits_vc_sel_1_3(input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_1_3),
    .io_salloc_req_0_bits_vc_sel_0_0(input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_0_0),
    .io_salloc_req_0_bits_vc_sel_0_1(input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_0_1),
    .io_salloc_req_0_bits_vc_sel_0_2(input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_0_2),
    .io_salloc_req_0_bits_vc_sel_0_3(input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_0_3),
    .io_salloc_req_0_bits_tail(input_unit_0_from_1_io_salloc_req_0_bits_tail),
    .io_out_0_valid(input_unit_0_from_1_io_out_0_valid),
    .io_out_0_bits_flit_head(input_unit_0_from_1_io_out_0_bits_flit_head),
    .io_out_0_bits_flit_tail(input_unit_0_from_1_io_out_0_bits_flit_tail),
    .io_out_0_bits_flit_payload(input_unit_0_from_1_io_out_0_bits_flit_payload),
    .io_out_0_bits_flit_flow_ingress_node(input_unit_0_from_1_io_out_0_bits_flit_flow_ingress_node),
    .io_out_0_bits_flit_flow_egress_node(input_unit_0_from_1_io_out_0_bits_flit_flow_egress_node),
    .io_out_0_bits_out_virt_channel(input_unit_0_from_1_io_out_0_bits_out_virt_channel),
    .io_debug_va_stall(input_unit_0_from_1_io_debug_va_stall),
    .io_debug_sa_stall(input_unit_0_from_1_io_debug_sa_stall),
    .io_in_flit_0_valid(input_unit_0_from_1_io_in_flit_0_valid),
    .io_in_flit_0_bits_head(input_unit_0_from_1_io_in_flit_0_bits_head),
    .io_in_flit_0_bits_tail(input_unit_0_from_1_io_in_flit_0_bits_tail),
    .io_in_flit_0_bits_payload(input_unit_0_from_1_io_in_flit_0_bits_payload),
    .io_in_flit_0_bits_flow_ingress_node(input_unit_0_from_1_io_in_flit_0_bits_flow_ingress_node),
    .io_in_flit_0_bits_flow_egress_node(input_unit_0_from_1_io_in_flit_0_bits_flow_egress_node),
    .io_in_flit_0_bits_virt_channel_id(input_unit_0_from_1_io_in_flit_0_bits_virt_channel_id),
    .io_in_credit_return(input_unit_0_from_1_io_in_credit_return),
    .io_in_vc_free(input_unit_0_from_1_io_in_vc_free)
  );
  InputUnit_1 input_unit_1_from_3 ( // @[Router.scala 112:13]
    .clock(input_unit_1_from_3_clock),
    .reset(input_unit_1_from_3_reset),
    .io_router_req_valid(input_unit_1_from_3_io_router_req_valid),
    .io_router_req_bits_src_virt_id(input_unit_1_from_3_io_router_req_bits_src_virt_id),
    .io_router_req_bits_flow_ingress_node(input_unit_1_from_3_io_router_req_bits_flow_ingress_node),
    .io_router_req_bits_flow_egress_node(input_unit_1_from_3_io_router_req_bits_flow_egress_node),
    .io_router_resp_vc_sel_1_0(input_unit_1_from_3_io_router_resp_vc_sel_1_0),
    .io_router_resp_vc_sel_1_1(input_unit_1_from_3_io_router_resp_vc_sel_1_1),
    .io_router_resp_vc_sel_1_2(input_unit_1_from_3_io_router_resp_vc_sel_1_2),
    .io_router_resp_vc_sel_0_0(input_unit_1_from_3_io_router_resp_vc_sel_0_0),
    .io_router_resp_vc_sel_0_1(input_unit_1_from_3_io_router_resp_vc_sel_0_1),
    .io_router_resp_vc_sel_0_2(input_unit_1_from_3_io_router_resp_vc_sel_0_2),
    .io_router_resp_vc_sel_0_3(input_unit_1_from_3_io_router_resp_vc_sel_0_3),
    .io_vcalloc_req_ready(input_unit_1_from_3_io_vcalloc_req_ready),
    .io_vcalloc_req_valid(input_unit_1_from_3_io_vcalloc_req_valid),
    .io_vcalloc_req_bits_vc_sel_2_0(input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_2_0),
    .io_vcalloc_req_bits_vc_sel_1_0(input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_1_0),
    .io_vcalloc_req_bits_vc_sel_1_1(input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_1_1),
    .io_vcalloc_req_bits_vc_sel_1_2(input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_1_2),
    .io_vcalloc_req_bits_vc_sel_0_0(input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_0_0),
    .io_vcalloc_req_bits_vc_sel_0_1(input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_0_1),
    .io_vcalloc_req_bits_vc_sel_0_2(input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_0_2),
    .io_vcalloc_req_bits_vc_sel_0_3(input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_0_3),
    .io_vcalloc_resp_vc_sel_2_0(input_unit_1_from_3_io_vcalloc_resp_vc_sel_2_0),
    .io_vcalloc_resp_vc_sel_1_0(input_unit_1_from_3_io_vcalloc_resp_vc_sel_1_0),
    .io_vcalloc_resp_vc_sel_1_1(input_unit_1_from_3_io_vcalloc_resp_vc_sel_1_1),
    .io_vcalloc_resp_vc_sel_1_2(input_unit_1_from_3_io_vcalloc_resp_vc_sel_1_2),
    .io_vcalloc_resp_vc_sel_0_0(input_unit_1_from_3_io_vcalloc_resp_vc_sel_0_0),
    .io_vcalloc_resp_vc_sel_0_1(input_unit_1_from_3_io_vcalloc_resp_vc_sel_0_1),
    .io_vcalloc_resp_vc_sel_0_2(input_unit_1_from_3_io_vcalloc_resp_vc_sel_0_2),
    .io_vcalloc_resp_vc_sel_0_3(input_unit_1_from_3_io_vcalloc_resp_vc_sel_0_3),
    .io_out_credit_available_2_0(input_unit_1_from_3_io_out_credit_available_2_0),
    .io_out_credit_available_1_0(input_unit_1_from_3_io_out_credit_available_1_0),
    .io_out_credit_available_1_1(input_unit_1_from_3_io_out_credit_available_1_1),
    .io_out_credit_available_1_2(input_unit_1_from_3_io_out_credit_available_1_2),
    .io_out_credit_available_1_3(input_unit_1_from_3_io_out_credit_available_1_3),
    .io_out_credit_available_0_0(input_unit_1_from_3_io_out_credit_available_0_0),
    .io_out_credit_available_0_1(input_unit_1_from_3_io_out_credit_available_0_1),
    .io_out_credit_available_0_2(input_unit_1_from_3_io_out_credit_available_0_2),
    .io_out_credit_available_0_3(input_unit_1_from_3_io_out_credit_available_0_3),
    .io_salloc_req_0_ready(input_unit_1_from_3_io_salloc_req_0_ready),
    .io_salloc_req_0_valid(input_unit_1_from_3_io_salloc_req_0_valid),
    .io_salloc_req_0_bits_vc_sel_2_0(input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_2_0),
    .io_salloc_req_0_bits_vc_sel_1_0(input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_1_0),
    .io_salloc_req_0_bits_vc_sel_1_1(input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_1_1),
    .io_salloc_req_0_bits_vc_sel_1_2(input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_1_2),
    .io_salloc_req_0_bits_vc_sel_1_3(input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_1_3),
    .io_salloc_req_0_bits_vc_sel_0_0(input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_0_0),
    .io_salloc_req_0_bits_vc_sel_0_1(input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_0_1),
    .io_salloc_req_0_bits_vc_sel_0_2(input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_0_2),
    .io_salloc_req_0_bits_vc_sel_0_3(input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_0_3),
    .io_salloc_req_0_bits_tail(input_unit_1_from_3_io_salloc_req_0_bits_tail),
    .io_out_0_valid(input_unit_1_from_3_io_out_0_valid),
    .io_out_0_bits_flit_head(input_unit_1_from_3_io_out_0_bits_flit_head),
    .io_out_0_bits_flit_tail(input_unit_1_from_3_io_out_0_bits_flit_tail),
    .io_out_0_bits_flit_payload(input_unit_1_from_3_io_out_0_bits_flit_payload),
    .io_out_0_bits_flit_flow_ingress_node(input_unit_1_from_3_io_out_0_bits_flit_flow_ingress_node),
    .io_out_0_bits_flit_flow_egress_node(input_unit_1_from_3_io_out_0_bits_flit_flow_egress_node),
    .io_out_0_bits_out_virt_channel(input_unit_1_from_3_io_out_0_bits_out_virt_channel),
    .io_debug_va_stall(input_unit_1_from_3_io_debug_va_stall),
    .io_debug_sa_stall(input_unit_1_from_3_io_debug_sa_stall),
    .io_in_flit_0_valid(input_unit_1_from_3_io_in_flit_0_valid),
    .io_in_flit_0_bits_head(input_unit_1_from_3_io_in_flit_0_bits_head),
    .io_in_flit_0_bits_tail(input_unit_1_from_3_io_in_flit_0_bits_tail),
    .io_in_flit_0_bits_payload(input_unit_1_from_3_io_in_flit_0_bits_payload),
    .io_in_flit_0_bits_flow_ingress_node(input_unit_1_from_3_io_in_flit_0_bits_flow_ingress_node),
    .io_in_flit_0_bits_flow_egress_node(input_unit_1_from_3_io_in_flit_0_bits_flow_egress_node),
    .io_in_flit_0_bits_virt_channel_id(input_unit_1_from_3_io_in_flit_0_bits_virt_channel_id),
    .io_in_credit_return(input_unit_1_from_3_io_in_credit_return),
    .io_in_vc_free(input_unit_1_from_3_io_in_vc_free)
  );
  IngressUnit ingress_unit_2_from_0 ( // @[Router.scala 116:13]
    .clock(ingress_unit_2_from_0_clock),
    .reset(ingress_unit_2_from_0_reset),
    .io_router_req_valid(ingress_unit_2_from_0_io_router_req_valid),
    .io_router_req_bits_flow_ingress_node(ingress_unit_2_from_0_io_router_req_bits_flow_ingress_node),
    .io_router_req_bits_flow_egress_node(ingress_unit_2_from_0_io_router_req_bits_flow_egress_node),
    .io_router_resp_vc_sel_1_0(ingress_unit_2_from_0_io_router_resp_vc_sel_1_0),
    .io_router_resp_vc_sel_1_1(ingress_unit_2_from_0_io_router_resp_vc_sel_1_1),
    .io_router_resp_vc_sel_1_2(ingress_unit_2_from_0_io_router_resp_vc_sel_1_2),
    .io_router_resp_vc_sel_1_3(ingress_unit_2_from_0_io_router_resp_vc_sel_1_3),
    .io_router_resp_vc_sel_0_0(ingress_unit_2_from_0_io_router_resp_vc_sel_0_0),
    .io_router_resp_vc_sel_0_1(ingress_unit_2_from_0_io_router_resp_vc_sel_0_1),
    .io_router_resp_vc_sel_0_2(ingress_unit_2_from_0_io_router_resp_vc_sel_0_2),
    .io_router_resp_vc_sel_0_3(ingress_unit_2_from_0_io_router_resp_vc_sel_0_3),
    .io_vcalloc_req_ready(ingress_unit_2_from_0_io_vcalloc_req_ready),
    .io_vcalloc_req_valid(ingress_unit_2_from_0_io_vcalloc_req_valid),
    .io_vcalloc_req_bits_vc_sel_2_0(ingress_unit_2_from_0_io_vcalloc_req_bits_vc_sel_2_0),
    .io_vcalloc_req_bits_vc_sel_1_0(ingress_unit_2_from_0_io_vcalloc_req_bits_vc_sel_1_0),
    .io_vcalloc_req_bits_vc_sel_1_1(ingress_unit_2_from_0_io_vcalloc_req_bits_vc_sel_1_1),
    .io_vcalloc_req_bits_vc_sel_1_2(ingress_unit_2_from_0_io_vcalloc_req_bits_vc_sel_1_2),
    .io_vcalloc_req_bits_vc_sel_1_3(ingress_unit_2_from_0_io_vcalloc_req_bits_vc_sel_1_3),
    .io_vcalloc_req_bits_vc_sel_0_0(ingress_unit_2_from_0_io_vcalloc_req_bits_vc_sel_0_0),
    .io_vcalloc_req_bits_vc_sel_0_1(ingress_unit_2_from_0_io_vcalloc_req_bits_vc_sel_0_1),
    .io_vcalloc_req_bits_vc_sel_0_2(ingress_unit_2_from_0_io_vcalloc_req_bits_vc_sel_0_2),
    .io_vcalloc_req_bits_vc_sel_0_3(ingress_unit_2_from_0_io_vcalloc_req_bits_vc_sel_0_3),
    .io_vcalloc_resp_vc_sel_2_0(ingress_unit_2_from_0_io_vcalloc_resp_vc_sel_2_0),
    .io_vcalloc_resp_vc_sel_1_0(ingress_unit_2_from_0_io_vcalloc_resp_vc_sel_1_0),
    .io_vcalloc_resp_vc_sel_1_1(ingress_unit_2_from_0_io_vcalloc_resp_vc_sel_1_1),
    .io_vcalloc_resp_vc_sel_1_2(ingress_unit_2_from_0_io_vcalloc_resp_vc_sel_1_2),
    .io_vcalloc_resp_vc_sel_1_3(ingress_unit_2_from_0_io_vcalloc_resp_vc_sel_1_3),
    .io_vcalloc_resp_vc_sel_0_0(ingress_unit_2_from_0_io_vcalloc_resp_vc_sel_0_0),
    .io_vcalloc_resp_vc_sel_0_1(ingress_unit_2_from_0_io_vcalloc_resp_vc_sel_0_1),
    .io_vcalloc_resp_vc_sel_0_2(ingress_unit_2_from_0_io_vcalloc_resp_vc_sel_0_2),
    .io_vcalloc_resp_vc_sel_0_3(ingress_unit_2_from_0_io_vcalloc_resp_vc_sel_0_3),
    .io_out_credit_available_2_0(ingress_unit_2_from_0_io_out_credit_available_2_0),
    .io_out_credit_available_1_0(ingress_unit_2_from_0_io_out_credit_available_1_0),
    .io_out_credit_available_1_1(ingress_unit_2_from_0_io_out_credit_available_1_1),
    .io_out_credit_available_1_2(ingress_unit_2_from_0_io_out_credit_available_1_2),
    .io_out_credit_available_1_3(ingress_unit_2_from_0_io_out_credit_available_1_3),
    .io_out_credit_available_0_0(ingress_unit_2_from_0_io_out_credit_available_0_0),
    .io_out_credit_available_0_1(ingress_unit_2_from_0_io_out_credit_available_0_1),
    .io_out_credit_available_0_2(ingress_unit_2_from_0_io_out_credit_available_0_2),
    .io_out_credit_available_0_3(ingress_unit_2_from_0_io_out_credit_available_0_3),
    .io_salloc_req_0_ready(ingress_unit_2_from_0_io_salloc_req_0_ready),
    .io_salloc_req_0_valid(ingress_unit_2_from_0_io_salloc_req_0_valid),
    .io_salloc_req_0_bits_vc_sel_2_0(ingress_unit_2_from_0_io_salloc_req_0_bits_vc_sel_2_0),
    .io_salloc_req_0_bits_vc_sel_1_0(ingress_unit_2_from_0_io_salloc_req_0_bits_vc_sel_1_0),
    .io_salloc_req_0_bits_vc_sel_1_1(ingress_unit_2_from_0_io_salloc_req_0_bits_vc_sel_1_1),
    .io_salloc_req_0_bits_vc_sel_1_2(ingress_unit_2_from_0_io_salloc_req_0_bits_vc_sel_1_2),
    .io_salloc_req_0_bits_vc_sel_1_3(ingress_unit_2_from_0_io_salloc_req_0_bits_vc_sel_1_3),
    .io_salloc_req_0_bits_vc_sel_0_0(ingress_unit_2_from_0_io_salloc_req_0_bits_vc_sel_0_0),
    .io_salloc_req_0_bits_vc_sel_0_1(ingress_unit_2_from_0_io_salloc_req_0_bits_vc_sel_0_1),
    .io_salloc_req_0_bits_vc_sel_0_2(ingress_unit_2_from_0_io_salloc_req_0_bits_vc_sel_0_2),
    .io_salloc_req_0_bits_vc_sel_0_3(ingress_unit_2_from_0_io_salloc_req_0_bits_vc_sel_0_3),
    .io_salloc_req_0_bits_tail(ingress_unit_2_from_0_io_salloc_req_0_bits_tail),
    .io_out_0_valid(ingress_unit_2_from_0_io_out_0_valid),
    .io_out_0_bits_flit_head(ingress_unit_2_from_0_io_out_0_bits_flit_head),
    .io_out_0_bits_flit_tail(ingress_unit_2_from_0_io_out_0_bits_flit_tail),
    .io_out_0_bits_flit_payload(ingress_unit_2_from_0_io_out_0_bits_flit_payload),
    .io_out_0_bits_flit_flow_ingress_node(ingress_unit_2_from_0_io_out_0_bits_flit_flow_ingress_node),
    .io_out_0_bits_flit_flow_egress_node(ingress_unit_2_from_0_io_out_0_bits_flit_flow_egress_node),
    .io_out_0_bits_out_virt_channel(ingress_unit_2_from_0_io_out_0_bits_out_virt_channel),
    .io_in_ready(ingress_unit_2_from_0_io_in_ready),
    .io_in_valid(ingress_unit_2_from_0_io_in_valid),
    .io_in_bits_head(ingress_unit_2_from_0_io_in_bits_head),
    .io_in_bits_tail(ingress_unit_2_from_0_io_in_bits_tail),
    .io_in_bits_payload(ingress_unit_2_from_0_io_in_bits_payload),
    .io_in_bits_egress_id(ingress_unit_2_from_0_io_in_bits_egress_id)
  );
  OutputUnit output_unit_0_to_1 ( // @[Router.scala 122:13]
    .clock(output_unit_0_to_1_clock),
    .reset(output_unit_0_to_1_reset),
    .io_in_0_valid(output_unit_0_to_1_io_in_0_valid),
    .io_in_0_bits_head(output_unit_0_to_1_io_in_0_bits_head),
    .io_in_0_bits_tail(output_unit_0_to_1_io_in_0_bits_tail),
    .io_in_0_bits_payload(output_unit_0_to_1_io_in_0_bits_payload),
    .io_in_0_bits_flow_ingress_node(output_unit_0_to_1_io_in_0_bits_flow_ingress_node),
    .io_in_0_bits_flow_egress_node(output_unit_0_to_1_io_in_0_bits_flow_egress_node),
    .io_in_0_bits_virt_channel_id(output_unit_0_to_1_io_in_0_bits_virt_channel_id),
    .io_credit_available_0(output_unit_0_to_1_io_credit_available_0),
    .io_credit_available_1(output_unit_0_to_1_io_credit_available_1),
    .io_credit_available_2(output_unit_0_to_1_io_credit_available_2),
    .io_credit_available_3(output_unit_0_to_1_io_credit_available_3),
    .io_channel_status_0_occupied(output_unit_0_to_1_io_channel_status_0_occupied),
    .io_channel_status_1_occupied(output_unit_0_to_1_io_channel_status_1_occupied),
    .io_channel_status_2_occupied(output_unit_0_to_1_io_channel_status_2_occupied),
    .io_channel_status_3_occupied(output_unit_0_to_1_io_channel_status_3_occupied),
    .io_allocs_0_alloc(output_unit_0_to_1_io_allocs_0_alloc),
    .io_allocs_1_alloc(output_unit_0_to_1_io_allocs_1_alloc),
    .io_allocs_2_alloc(output_unit_0_to_1_io_allocs_2_alloc),
    .io_allocs_3_alloc(output_unit_0_to_1_io_allocs_3_alloc),
    .io_credit_alloc_0_alloc(output_unit_0_to_1_io_credit_alloc_0_alloc),
    .io_credit_alloc_1_alloc(output_unit_0_to_1_io_credit_alloc_1_alloc),
    .io_credit_alloc_2_alloc(output_unit_0_to_1_io_credit_alloc_2_alloc),
    .io_credit_alloc_3_alloc(output_unit_0_to_1_io_credit_alloc_3_alloc),
    .io_out_flit_0_valid(output_unit_0_to_1_io_out_flit_0_valid),
    .io_out_flit_0_bits_head(output_unit_0_to_1_io_out_flit_0_bits_head),
    .io_out_flit_0_bits_tail(output_unit_0_to_1_io_out_flit_0_bits_tail),
    .io_out_flit_0_bits_payload(output_unit_0_to_1_io_out_flit_0_bits_payload),
    .io_out_flit_0_bits_flow_ingress_node(output_unit_0_to_1_io_out_flit_0_bits_flow_ingress_node),
    .io_out_flit_0_bits_flow_egress_node(output_unit_0_to_1_io_out_flit_0_bits_flow_egress_node),
    .io_out_flit_0_bits_virt_channel_id(output_unit_0_to_1_io_out_flit_0_bits_virt_channel_id),
    .io_out_credit_return(output_unit_0_to_1_io_out_credit_return),
    .io_out_vc_free(output_unit_0_to_1_io_out_vc_free)
  );
  OutputUnit output_unit_1_to_3 ( // @[Router.scala 122:13]
    .clock(output_unit_1_to_3_clock),
    .reset(output_unit_1_to_3_reset),
    .io_in_0_valid(output_unit_1_to_3_io_in_0_valid),
    .io_in_0_bits_head(output_unit_1_to_3_io_in_0_bits_head),
    .io_in_0_bits_tail(output_unit_1_to_3_io_in_0_bits_tail),
    .io_in_0_bits_payload(output_unit_1_to_3_io_in_0_bits_payload),
    .io_in_0_bits_flow_ingress_node(output_unit_1_to_3_io_in_0_bits_flow_ingress_node),
    .io_in_0_bits_flow_egress_node(output_unit_1_to_3_io_in_0_bits_flow_egress_node),
    .io_in_0_bits_virt_channel_id(output_unit_1_to_3_io_in_0_bits_virt_channel_id),
    .io_credit_available_0(output_unit_1_to_3_io_credit_available_0),
    .io_credit_available_1(output_unit_1_to_3_io_credit_available_1),
    .io_credit_available_2(output_unit_1_to_3_io_credit_available_2),
    .io_credit_available_3(output_unit_1_to_3_io_credit_available_3),
    .io_channel_status_0_occupied(output_unit_1_to_3_io_channel_status_0_occupied),
    .io_channel_status_1_occupied(output_unit_1_to_3_io_channel_status_1_occupied),
    .io_channel_status_2_occupied(output_unit_1_to_3_io_channel_status_2_occupied),
    .io_channel_status_3_occupied(output_unit_1_to_3_io_channel_status_3_occupied),
    .io_allocs_0_alloc(output_unit_1_to_3_io_allocs_0_alloc),
    .io_allocs_1_alloc(output_unit_1_to_3_io_allocs_1_alloc),
    .io_allocs_2_alloc(output_unit_1_to_3_io_allocs_2_alloc),
    .io_allocs_3_alloc(output_unit_1_to_3_io_allocs_3_alloc),
    .io_credit_alloc_0_alloc(output_unit_1_to_3_io_credit_alloc_0_alloc),
    .io_credit_alloc_1_alloc(output_unit_1_to_3_io_credit_alloc_1_alloc),
    .io_credit_alloc_2_alloc(output_unit_1_to_3_io_credit_alloc_2_alloc),
    .io_credit_alloc_3_alloc(output_unit_1_to_3_io_credit_alloc_3_alloc),
    .io_out_flit_0_valid(output_unit_1_to_3_io_out_flit_0_valid),
    .io_out_flit_0_bits_head(output_unit_1_to_3_io_out_flit_0_bits_head),
    .io_out_flit_0_bits_tail(output_unit_1_to_3_io_out_flit_0_bits_tail),
    .io_out_flit_0_bits_payload(output_unit_1_to_3_io_out_flit_0_bits_payload),
    .io_out_flit_0_bits_flow_ingress_node(output_unit_1_to_3_io_out_flit_0_bits_flow_ingress_node),
    .io_out_flit_0_bits_flow_egress_node(output_unit_1_to_3_io_out_flit_0_bits_flow_egress_node),
    .io_out_flit_0_bits_virt_channel_id(output_unit_1_to_3_io_out_flit_0_bits_virt_channel_id),
    .io_out_credit_return(output_unit_1_to_3_io_out_credit_return),
    .io_out_vc_free(output_unit_1_to_3_io_out_vc_free)
  );
  EgressUnit egress_unit_2_to_0 ( // @[Router.scala 125:13]
    .clock(egress_unit_2_to_0_clock),
    .reset(egress_unit_2_to_0_reset),
    .io_in_0_valid(egress_unit_2_to_0_io_in_0_valid),
    .io_in_0_bits_head(egress_unit_2_to_0_io_in_0_bits_head),
    .io_in_0_bits_tail(egress_unit_2_to_0_io_in_0_bits_tail),
    .io_in_0_bits_payload(egress_unit_2_to_0_io_in_0_bits_payload),
    .io_in_0_bits_flow_ingress_node(egress_unit_2_to_0_io_in_0_bits_flow_ingress_node),
    .io_credit_available_0(egress_unit_2_to_0_io_credit_available_0),
    .io_channel_status_0_occupied(egress_unit_2_to_0_io_channel_status_0_occupied),
    .io_allocs_0_alloc(egress_unit_2_to_0_io_allocs_0_alloc),
    .io_credit_alloc_0_alloc(egress_unit_2_to_0_io_credit_alloc_0_alloc),
    .io_credit_alloc_0_tail(egress_unit_2_to_0_io_credit_alloc_0_tail),
    .io_out_valid(egress_unit_2_to_0_io_out_valid),
    .io_out_bits_head(egress_unit_2_to_0_io_out_bits_head),
    .io_out_bits_tail(egress_unit_2_to_0_io_out_bits_tail),
    .io_out_bits_payload(egress_unit_2_to_0_io_out_bits_payload),
    .io_out_bits_ingress_id(egress_unit_2_to_0_io_out_bits_ingress_id)
  );
  Switch switch ( // @[Router.scala 129:24]
    .clock(switch_clock),
    .reset(switch_reset),
    .io_in_2_0_valid(switch_io_in_2_0_valid),
    .io_in_2_0_bits_flit_head(switch_io_in_2_0_bits_flit_head),
    .io_in_2_0_bits_flit_tail(switch_io_in_2_0_bits_flit_tail),
    .io_in_2_0_bits_flit_payload(switch_io_in_2_0_bits_flit_payload),
    .io_in_2_0_bits_flit_flow_ingress_node(switch_io_in_2_0_bits_flit_flow_ingress_node),
    .io_in_2_0_bits_flit_flow_egress_node(switch_io_in_2_0_bits_flit_flow_egress_node),
    .io_in_2_0_bits_out_virt_channel(switch_io_in_2_0_bits_out_virt_channel),
    .io_in_1_0_valid(switch_io_in_1_0_valid),
    .io_in_1_0_bits_flit_head(switch_io_in_1_0_bits_flit_head),
    .io_in_1_0_bits_flit_tail(switch_io_in_1_0_bits_flit_tail),
    .io_in_1_0_bits_flit_payload(switch_io_in_1_0_bits_flit_payload),
    .io_in_1_0_bits_flit_flow_ingress_node(switch_io_in_1_0_bits_flit_flow_ingress_node),
    .io_in_1_0_bits_flit_flow_egress_node(switch_io_in_1_0_bits_flit_flow_egress_node),
    .io_in_1_0_bits_out_virt_channel(switch_io_in_1_0_bits_out_virt_channel),
    .io_in_0_0_valid(switch_io_in_0_0_valid),
    .io_in_0_0_bits_flit_head(switch_io_in_0_0_bits_flit_head),
    .io_in_0_0_bits_flit_tail(switch_io_in_0_0_bits_flit_tail),
    .io_in_0_0_bits_flit_payload(switch_io_in_0_0_bits_flit_payload),
    .io_in_0_0_bits_flit_flow_ingress_node(switch_io_in_0_0_bits_flit_flow_ingress_node),
    .io_in_0_0_bits_flit_flow_egress_node(switch_io_in_0_0_bits_flit_flow_egress_node),
    .io_in_0_0_bits_out_virt_channel(switch_io_in_0_0_bits_out_virt_channel),
    .io_out_2_0_valid(switch_io_out_2_0_valid),
    .io_out_2_0_bits_head(switch_io_out_2_0_bits_head),
    .io_out_2_0_bits_tail(switch_io_out_2_0_bits_tail),
    .io_out_2_0_bits_payload(switch_io_out_2_0_bits_payload),
    .io_out_2_0_bits_flow_ingress_node(switch_io_out_2_0_bits_flow_ingress_node),
    .io_out_1_0_valid(switch_io_out_1_0_valid),
    .io_out_1_0_bits_head(switch_io_out_1_0_bits_head),
    .io_out_1_0_bits_tail(switch_io_out_1_0_bits_tail),
    .io_out_1_0_bits_payload(switch_io_out_1_0_bits_payload),
    .io_out_1_0_bits_flow_ingress_node(switch_io_out_1_0_bits_flow_ingress_node),
    .io_out_1_0_bits_flow_egress_node(switch_io_out_1_0_bits_flow_egress_node),
    .io_out_1_0_bits_virt_channel_id(switch_io_out_1_0_bits_virt_channel_id),
    .io_out_0_0_valid(switch_io_out_0_0_valid),
    .io_out_0_0_bits_head(switch_io_out_0_0_bits_head),
    .io_out_0_0_bits_tail(switch_io_out_0_0_bits_tail),
    .io_out_0_0_bits_payload(switch_io_out_0_0_bits_payload),
    .io_out_0_0_bits_flow_ingress_node(switch_io_out_0_0_bits_flow_ingress_node),
    .io_out_0_0_bits_flow_egress_node(switch_io_out_0_0_bits_flow_egress_node),
    .io_out_0_0_bits_virt_channel_id(switch_io_out_0_0_bits_virt_channel_id),
    .io_sel_2_0_2_0(switch_io_sel_2_0_2_0),
    .io_sel_2_0_1_0(switch_io_sel_2_0_1_0),
    .io_sel_2_0_0_0(switch_io_sel_2_0_0_0),
    .io_sel_1_0_2_0(switch_io_sel_1_0_2_0),
    .io_sel_1_0_1_0(switch_io_sel_1_0_1_0),
    .io_sel_1_0_0_0(switch_io_sel_1_0_0_0),
    .io_sel_0_0_2_0(switch_io_sel_0_0_2_0),
    .io_sel_0_0_1_0(switch_io_sel_0_0_1_0),
    .io_sel_0_0_0_0(switch_io_sel_0_0_0_0)
  );
  SwitchAllocator switch_allocator ( // @[Router.scala 130:34]
    .clock(switch_allocator_clock),
    .reset(switch_allocator_reset),
    .io_req_2_0_ready(switch_allocator_io_req_2_0_ready),
    .io_req_2_0_valid(switch_allocator_io_req_2_0_valid),
    .io_req_2_0_bits_vc_sel_2_0(switch_allocator_io_req_2_0_bits_vc_sel_2_0),
    .io_req_2_0_bits_vc_sel_1_0(switch_allocator_io_req_2_0_bits_vc_sel_1_0),
    .io_req_2_0_bits_vc_sel_1_1(switch_allocator_io_req_2_0_bits_vc_sel_1_1),
    .io_req_2_0_bits_vc_sel_1_2(switch_allocator_io_req_2_0_bits_vc_sel_1_2),
    .io_req_2_0_bits_vc_sel_1_3(switch_allocator_io_req_2_0_bits_vc_sel_1_3),
    .io_req_2_0_bits_vc_sel_0_0(switch_allocator_io_req_2_0_bits_vc_sel_0_0),
    .io_req_2_0_bits_vc_sel_0_1(switch_allocator_io_req_2_0_bits_vc_sel_0_1),
    .io_req_2_0_bits_vc_sel_0_2(switch_allocator_io_req_2_0_bits_vc_sel_0_2),
    .io_req_2_0_bits_vc_sel_0_3(switch_allocator_io_req_2_0_bits_vc_sel_0_3),
    .io_req_2_0_bits_tail(switch_allocator_io_req_2_0_bits_tail),
    .io_req_1_0_ready(switch_allocator_io_req_1_0_ready),
    .io_req_1_0_valid(switch_allocator_io_req_1_0_valid),
    .io_req_1_0_bits_vc_sel_2_0(switch_allocator_io_req_1_0_bits_vc_sel_2_0),
    .io_req_1_0_bits_vc_sel_1_0(switch_allocator_io_req_1_0_bits_vc_sel_1_0),
    .io_req_1_0_bits_vc_sel_1_1(switch_allocator_io_req_1_0_bits_vc_sel_1_1),
    .io_req_1_0_bits_vc_sel_1_2(switch_allocator_io_req_1_0_bits_vc_sel_1_2),
    .io_req_1_0_bits_vc_sel_1_3(switch_allocator_io_req_1_0_bits_vc_sel_1_3),
    .io_req_1_0_bits_vc_sel_0_0(switch_allocator_io_req_1_0_bits_vc_sel_0_0),
    .io_req_1_0_bits_vc_sel_0_1(switch_allocator_io_req_1_0_bits_vc_sel_0_1),
    .io_req_1_0_bits_vc_sel_0_2(switch_allocator_io_req_1_0_bits_vc_sel_0_2),
    .io_req_1_0_bits_vc_sel_0_3(switch_allocator_io_req_1_0_bits_vc_sel_0_3),
    .io_req_1_0_bits_tail(switch_allocator_io_req_1_0_bits_tail),
    .io_req_0_0_ready(switch_allocator_io_req_0_0_ready),
    .io_req_0_0_valid(switch_allocator_io_req_0_0_valid),
    .io_req_0_0_bits_vc_sel_2_0(switch_allocator_io_req_0_0_bits_vc_sel_2_0),
    .io_req_0_0_bits_vc_sel_1_0(switch_allocator_io_req_0_0_bits_vc_sel_1_0),
    .io_req_0_0_bits_vc_sel_1_1(switch_allocator_io_req_0_0_bits_vc_sel_1_1),
    .io_req_0_0_bits_vc_sel_1_2(switch_allocator_io_req_0_0_bits_vc_sel_1_2),
    .io_req_0_0_bits_vc_sel_1_3(switch_allocator_io_req_0_0_bits_vc_sel_1_3),
    .io_req_0_0_bits_vc_sel_0_0(switch_allocator_io_req_0_0_bits_vc_sel_0_0),
    .io_req_0_0_bits_vc_sel_0_1(switch_allocator_io_req_0_0_bits_vc_sel_0_1),
    .io_req_0_0_bits_vc_sel_0_2(switch_allocator_io_req_0_0_bits_vc_sel_0_2),
    .io_req_0_0_bits_vc_sel_0_3(switch_allocator_io_req_0_0_bits_vc_sel_0_3),
    .io_req_0_0_bits_tail(switch_allocator_io_req_0_0_bits_tail),
    .io_credit_alloc_2_0_alloc(switch_allocator_io_credit_alloc_2_0_alloc),
    .io_credit_alloc_2_0_tail(switch_allocator_io_credit_alloc_2_0_tail),
    .io_credit_alloc_1_0_alloc(switch_allocator_io_credit_alloc_1_0_alloc),
    .io_credit_alloc_1_1_alloc(switch_allocator_io_credit_alloc_1_1_alloc),
    .io_credit_alloc_1_2_alloc(switch_allocator_io_credit_alloc_1_2_alloc),
    .io_credit_alloc_1_3_alloc(switch_allocator_io_credit_alloc_1_3_alloc),
    .io_credit_alloc_0_0_alloc(switch_allocator_io_credit_alloc_0_0_alloc),
    .io_credit_alloc_0_1_alloc(switch_allocator_io_credit_alloc_0_1_alloc),
    .io_credit_alloc_0_2_alloc(switch_allocator_io_credit_alloc_0_2_alloc),
    .io_credit_alloc_0_3_alloc(switch_allocator_io_credit_alloc_0_3_alloc),
    .io_switch_sel_2_0_2_0(switch_allocator_io_switch_sel_2_0_2_0),
    .io_switch_sel_2_0_1_0(switch_allocator_io_switch_sel_2_0_1_0),
    .io_switch_sel_2_0_0_0(switch_allocator_io_switch_sel_2_0_0_0),
    .io_switch_sel_1_0_2_0(switch_allocator_io_switch_sel_1_0_2_0),
    .io_switch_sel_1_0_1_0(switch_allocator_io_switch_sel_1_0_1_0),
    .io_switch_sel_1_0_0_0(switch_allocator_io_switch_sel_1_0_0_0),
    .io_switch_sel_0_0_2_0(switch_allocator_io_switch_sel_0_0_2_0),
    .io_switch_sel_0_0_1_0(switch_allocator_io_switch_sel_0_0_1_0),
    .io_switch_sel_0_0_0_0(switch_allocator_io_switch_sel_0_0_0_0)
  );
  RotatingSingleVCAllocator vc_allocator ( // @[Router.scala 131:30]
    .clock(vc_allocator_clock),
    .reset(vc_allocator_reset),
    .io_req_2_ready(vc_allocator_io_req_2_ready),
    .io_req_2_valid(vc_allocator_io_req_2_valid),
    .io_req_2_bits_vc_sel_2_0(vc_allocator_io_req_2_bits_vc_sel_2_0),
    .io_req_2_bits_vc_sel_1_0(vc_allocator_io_req_2_bits_vc_sel_1_0),
    .io_req_2_bits_vc_sel_1_1(vc_allocator_io_req_2_bits_vc_sel_1_1),
    .io_req_2_bits_vc_sel_1_2(vc_allocator_io_req_2_bits_vc_sel_1_2),
    .io_req_2_bits_vc_sel_1_3(vc_allocator_io_req_2_bits_vc_sel_1_3),
    .io_req_2_bits_vc_sel_0_0(vc_allocator_io_req_2_bits_vc_sel_0_0),
    .io_req_2_bits_vc_sel_0_1(vc_allocator_io_req_2_bits_vc_sel_0_1),
    .io_req_2_bits_vc_sel_0_2(vc_allocator_io_req_2_bits_vc_sel_0_2),
    .io_req_2_bits_vc_sel_0_3(vc_allocator_io_req_2_bits_vc_sel_0_3),
    .io_req_1_ready(vc_allocator_io_req_1_ready),
    .io_req_1_valid(vc_allocator_io_req_1_valid),
    .io_req_1_bits_vc_sel_2_0(vc_allocator_io_req_1_bits_vc_sel_2_0),
    .io_req_1_bits_vc_sel_1_0(vc_allocator_io_req_1_bits_vc_sel_1_0),
    .io_req_1_bits_vc_sel_1_1(vc_allocator_io_req_1_bits_vc_sel_1_1),
    .io_req_1_bits_vc_sel_1_2(vc_allocator_io_req_1_bits_vc_sel_1_2),
    .io_req_1_bits_vc_sel_1_3(vc_allocator_io_req_1_bits_vc_sel_1_3),
    .io_req_1_bits_vc_sel_0_0(vc_allocator_io_req_1_bits_vc_sel_0_0),
    .io_req_1_bits_vc_sel_0_1(vc_allocator_io_req_1_bits_vc_sel_0_1),
    .io_req_1_bits_vc_sel_0_2(vc_allocator_io_req_1_bits_vc_sel_0_2),
    .io_req_1_bits_vc_sel_0_3(vc_allocator_io_req_1_bits_vc_sel_0_3),
    .io_req_0_ready(vc_allocator_io_req_0_ready),
    .io_req_0_valid(vc_allocator_io_req_0_valid),
    .io_req_0_bits_vc_sel_2_0(vc_allocator_io_req_0_bits_vc_sel_2_0),
    .io_req_0_bits_vc_sel_1_0(vc_allocator_io_req_0_bits_vc_sel_1_0),
    .io_req_0_bits_vc_sel_1_1(vc_allocator_io_req_0_bits_vc_sel_1_1),
    .io_req_0_bits_vc_sel_1_2(vc_allocator_io_req_0_bits_vc_sel_1_2),
    .io_req_0_bits_vc_sel_1_3(vc_allocator_io_req_0_bits_vc_sel_1_3),
    .io_req_0_bits_vc_sel_0_0(vc_allocator_io_req_0_bits_vc_sel_0_0),
    .io_req_0_bits_vc_sel_0_1(vc_allocator_io_req_0_bits_vc_sel_0_1),
    .io_req_0_bits_vc_sel_0_2(vc_allocator_io_req_0_bits_vc_sel_0_2),
    .io_req_0_bits_vc_sel_0_3(vc_allocator_io_req_0_bits_vc_sel_0_3),
    .io_resp_2_vc_sel_2_0(vc_allocator_io_resp_2_vc_sel_2_0),
    .io_resp_2_vc_sel_1_0(vc_allocator_io_resp_2_vc_sel_1_0),
    .io_resp_2_vc_sel_1_1(vc_allocator_io_resp_2_vc_sel_1_1),
    .io_resp_2_vc_sel_1_2(vc_allocator_io_resp_2_vc_sel_1_2),
    .io_resp_2_vc_sel_1_3(vc_allocator_io_resp_2_vc_sel_1_3),
    .io_resp_2_vc_sel_0_0(vc_allocator_io_resp_2_vc_sel_0_0),
    .io_resp_2_vc_sel_0_1(vc_allocator_io_resp_2_vc_sel_0_1),
    .io_resp_2_vc_sel_0_2(vc_allocator_io_resp_2_vc_sel_0_2),
    .io_resp_2_vc_sel_0_3(vc_allocator_io_resp_2_vc_sel_0_3),
    .io_resp_1_vc_sel_2_0(vc_allocator_io_resp_1_vc_sel_2_0),
    .io_resp_1_vc_sel_1_0(vc_allocator_io_resp_1_vc_sel_1_0),
    .io_resp_1_vc_sel_1_1(vc_allocator_io_resp_1_vc_sel_1_1),
    .io_resp_1_vc_sel_1_2(vc_allocator_io_resp_1_vc_sel_1_2),
    .io_resp_1_vc_sel_1_3(vc_allocator_io_resp_1_vc_sel_1_3),
    .io_resp_1_vc_sel_0_0(vc_allocator_io_resp_1_vc_sel_0_0),
    .io_resp_1_vc_sel_0_1(vc_allocator_io_resp_1_vc_sel_0_1),
    .io_resp_1_vc_sel_0_2(vc_allocator_io_resp_1_vc_sel_0_2),
    .io_resp_1_vc_sel_0_3(vc_allocator_io_resp_1_vc_sel_0_3),
    .io_resp_0_vc_sel_2_0(vc_allocator_io_resp_0_vc_sel_2_0),
    .io_resp_0_vc_sel_1_0(vc_allocator_io_resp_0_vc_sel_1_0),
    .io_resp_0_vc_sel_1_1(vc_allocator_io_resp_0_vc_sel_1_1),
    .io_resp_0_vc_sel_1_2(vc_allocator_io_resp_0_vc_sel_1_2),
    .io_resp_0_vc_sel_1_3(vc_allocator_io_resp_0_vc_sel_1_3),
    .io_resp_0_vc_sel_0_0(vc_allocator_io_resp_0_vc_sel_0_0),
    .io_resp_0_vc_sel_0_1(vc_allocator_io_resp_0_vc_sel_0_1),
    .io_resp_0_vc_sel_0_2(vc_allocator_io_resp_0_vc_sel_0_2),
    .io_resp_0_vc_sel_0_3(vc_allocator_io_resp_0_vc_sel_0_3),
    .io_channel_status_2_0_occupied(vc_allocator_io_channel_status_2_0_occupied),
    .io_channel_status_1_0_occupied(vc_allocator_io_channel_status_1_0_occupied),
    .io_channel_status_1_1_occupied(vc_allocator_io_channel_status_1_1_occupied),
    .io_channel_status_1_2_occupied(vc_allocator_io_channel_status_1_2_occupied),
    .io_channel_status_1_3_occupied(vc_allocator_io_channel_status_1_3_occupied),
    .io_channel_status_0_0_occupied(vc_allocator_io_channel_status_0_0_occupied),
    .io_channel_status_0_1_occupied(vc_allocator_io_channel_status_0_1_occupied),
    .io_channel_status_0_2_occupied(vc_allocator_io_channel_status_0_2_occupied),
    .io_channel_status_0_3_occupied(vc_allocator_io_channel_status_0_3_occupied),
    .io_out_allocs_2_0_alloc(vc_allocator_io_out_allocs_2_0_alloc),
    .io_out_allocs_1_0_alloc(vc_allocator_io_out_allocs_1_0_alloc),
    .io_out_allocs_1_1_alloc(vc_allocator_io_out_allocs_1_1_alloc),
    .io_out_allocs_1_2_alloc(vc_allocator_io_out_allocs_1_2_alloc),
    .io_out_allocs_1_3_alloc(vc_allocator_io_out_allocs_1_3_alloc),
    .io_out_allocs_0_0_alloc(vc_allocator_io_out_allocs_0_0_alloc),
    .io_out_allocs_0_1_alloc(vc_allocator_io_out_allocs_0_1_alloc),
    .io_out_allocs_0_2_alloc(vc_allocator_io_out_allocs_0_2_alloc),
    .io_out_allocs_0_3_alloc(vc_allocator_io_out_allocs_0_3_alloc)
  );
  RouteComputer route_computer ( // @[Router.scala 134:32]
    .io_req_2_bits_flow_ingress_node(route_computer_io_req_2_bits_flow_ingress_node),
    .io_req_2_bits_flow_egress_node(route_computer_io_req_2_bits_flow_egress_node),
    .io_req_1_bits_src_virt_id(route_computer_io_req_1_bits_src_virt_id),
    .io_req_1_bits_flow_ingress_node(route_computer_io_req_1_bits_flow_ingress_node),
    .io_req_1_bits_flow_egress_node(route_computer_io_req_1_bits_flow_egress_node),
    .io_req_0_bits_src_virt_id(route_computer_io_req_0_bits_src_virt_id),
    .io_req_0_bits_flow_ingress_node(route_computer_io_req_0_bits_flow_ingress_node),
    .io_req_0_bits_flow_egress_node(route_computer_io_req_0_bits_flow_egress_node),
    .io_resp_2_vc_sel_1_0(route_computer_io_resp_2_vc_sel_1_0),
    .io_resp_2_vc_sel_1_1(route_computer_io_resp_2_vc_sel_1_1),
    .io_resp_2_vc_sel_1_2(route_computer_io_resp_2_vc_sel_1_2),
    .io_resp_2_vc_sel_1_3(route_computer_io_resp_2_vc_sel_1_3),
    .io_resp_2_vc_sel_0_0(route_computer_io_resp_2_vc_sel_0_0),
    .io_resp_2_vc_sel_0_1(route_computer_io_resp_2_vc_sel_0_1),
    .io_resp_2_vc_sel_0_2(route_computer_io_resp_2_vc_sel_0_2),
    .io_resp_2_vc_sel_0_3(route_computer_io_resp_2_vc_sel_0_3),
    .io_resp_1_vc_sel_1_0(route_computer_io_resp_1_vc_sel_1_0),
    .io_resp_1_vc_sel_1_1(route_computer_io_resp_1_vc_sel_1_1),
    .io_resp_1_vc_sel_1_2(route_computer_io_resp_1_vc_sel_1_2),
    .io_resp_1_vc_sel_0_0(route_computer_io_resp_1_vc_sel_0_0),
    .io_resp_1_vc_sel_0_1(route_computer_io_resp_1_vc_sel_0_1),
    .io_resp_1_vc_sel_0_2(route_computer_io_resp_1_vc_sel_0_2),
    .io_resp_1_vc_sel_0_3(route_computer_io_resp_1_vc_sel_0_3),
    .io_resp_0_vc_sel_1_0(route_computer_io_resp_0_vc_sel_1_0),
    .io_resp_0_vc_sel_1_1(route_computer_io_resp_0_vc_sel_1_1),
    .io_resp_0_vc_sel_1_2(route_computer_io_resp_0_vc_sel_1_2),
    .io_resp_0_vc_sel_0_0(route_computer_io_resp_0_vc_sel_0_0),
    .io_resp_0_vc_sel_0_1(route_computer_io_resp_0_vc_sel_0_1),
    .io_resp_0_vc_sel_0_2(route_computer_io_resp_0_vc_sel_0_2),
    .io_resp_0_vc_sel_0_3(route_computer_io_resp_0_vc_sel_0_3)
  );
  plusarg_reader #(.FORMAT("noc_util_sample_rate=%d"), .DEFAULT(0), .WIDTH(20)) plusarg_reader ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_out)
  );
  assign auto_debug_out_va_stall_0 = input_unit_0_from_1_io_debug_va_stall; // @[Nodes.scala 1212:84 Router.scala 190:92]
  assign auto_debug_out_va_stall_1 = input_unit_1_from_3_io_debug_va_stall; // @[Nodes.scala 1212:84 Router.scala 190:92]
  assign auto_debug_out_sa_stall_0 = input_unit_0_from_1_io_debug_sa_stall; // @[Nodes.scala 1212:84 Router.scala 191:92]
  assign auto_debug_out_sa_stall_1 = input_unit_1_from_3_io_debug_sa_stall; // @[Nodes.scala 1212:84 Router.scala 191:92]
  assign auto_egress_nodes_out_flit_valid = egress_unit_2_to_0_io_out_valid; // @[Nodes.scala 1212:84 Router.scala 144:65]
  assign auto_egress_nodes_out_flit_bits_head = egress_unit_2_to_0_io_out_bits_head; // @[Nodes.scala 1212:84 Router.scala 144:65]
  assign auto_egress_nodes_out_flit_bits_tail = egress_unit_2_to_0_io_out_bits_tail; // @[Nodes.scala 1212:84 Router.scala 144:65]
  assign auto_egress_nodes_out_flit_bits_payload = egress_unit_2_to_0_io_out_bits_payload; // @[Nodes.scala 1212:84 Router.scala 144:65]
  assign auto_egress_nodes_out_flit_bits_ingress_id = egress_unit_2_to_0_io_out_bits_ingress_id; // @[Nodes.scala 1212:84 Router.scala 144:65]
  assign auto_ingress_nodes_in_flit_ready = ingress_unit_2_from_0_io_in_ready; // @[Nodes.scala 1215:84 Router.scala 142:68]
  assign auto_source_nodes_out_1_flit_0_valid = output_unit_1_to_3_io_out_flit_0_valid; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_1_flit_0_bits_head = output_unit_1_to_3_io_out_flit_0_bits_head; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_1_flit_0_bits_tail = output_unit_1_to_3_io_out_flit_0_bits_tail; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_1_flit_0_bits_payload = output_unit_1_to_3_io_out_flit_0_bits_payload; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_1_flit_0_bits_flow_ingress_node = output_unit_1_to_3_io_out_flit_0_bits_flow_ingress_node
    ; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_1_flit_0_bits_flow_egress_node = output_unit_1_to_3_io_out_flit_0_bits_flow_egress_node; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_1_flit_0_bits_virt_channel_id = output_unit_1_to_3_io_out_flit_0_bits_virt_channel_id; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_0_flit_0_valid = output_unit_0_to_1_io_out_flit_0_valid; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_0_flit_0_bits_head = output_unit_0_to_1_io_out_flit_0_bits_head; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_0_flit_0_bits_tail = output_unit_0_to_1_io_out_flit_0_bits_tail; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_0_flit_0_bits_payload = output_unit_0_to_1_io_out_flit_0_bits_payload; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_0_flit_0_bits_flow_ingress_node = output_unit_0_to_1_io_out_flit_0_bits_flow_ingress_node
    ; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_0_flit_0_bits_flow_egress_node = output_unit_0_to_1_io_out_flit_0_bits_flow_egress_node; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_0_flit_0_bits_virt_channel_id = output_unit_0_to_1_io_out_flit_0_bits_virt_channel_id; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_dest_nodes_in_1_credit_return = input_unit_1_from_3_io_in_credit_return; // @[Nodes.scala 1215:84 Router.scala 141:68]
  assign auto_dest_nodes_in_1_vc_free = input_unit_1_from_3_io_in_vc_free; // @[Nodes.scala 1215:84 Router.scala 141:68]
  assign auto_dest_nodes_in_0_credit_return = input_unit_0_from_1_io_in_credit_return; // @[Nodes.scala 1215:84 Router.scala 141:68]
  assign auto_dest_nodes_in_0_vc_free = input_unit_0_from_1_io_in_vc_free; // @[Nodes.scala 1215:84 Router.scala 141:68]
  assign monitor_clock = clock;
  assign monitor_reset = reset;
  assign monitor_io_in_flit_0_valid = auto_dest_nodes_in_0_flit_0_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_io_in_flit_0_bits_head = auto_dest_nodes_in_0_flit_0_bits_head; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_io_in_flit_0_bits_tail = auto_dest_nodes_in_0_flit_0_bits_tail; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_io_in_flit_0_bits_flow_ingress_node = auto_dest_nodes_in_0_flit_0_bits_flow_ingress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_io_in_flit_0_bits_flow_egress_node = auto_dest_nodes_in_0_flit_0_bits_flow_egress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_io_in_flit_0_bits_virt_channel_id = auto_dest_nodes_in_0_flit_0_bits_virt_channel_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_1_clock = clock;
  assign monitor_1_reset = reset;
  assign monitor_1_io_in_flit_0_valid = auto_dest_nodes_in_1_flit_0_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_1_io_in_flit_0_bits_head = auto_dest_nodes_in_1_flit_0_bits_head; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_1_io_in_flit_0_bits_tail = auto_dest_nodes_in_1_flit_0_bits_tail; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_1_io_in_flit_0_bits_flow_ingress_node = auto_dest_nodes_in_1_flit_0_bits_flow_ingress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_1_io_in_flit_0_bits_flow_egress_node = auto_dest_nodes_in_1_flit_0_bits_flow_egress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_1_io_in_flit_0_bits_virt_channel_id = auto_dest_nodes_in_1_flit_0_bits_virt_channel_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_1_clock = clock;
  assign input_unit_0_from_1_reset = reset;
  assign input_unit_0_from_1_io_router_resp_vc_sel_1_0 = route_computer_io_resp_0_vc_sel_1_0; // @[Router.scala 148:38]
  assign input_unit_0_from_1_io_router_resp_vc_sel_1_1 = route_computer_io_resp_0_vc_sel_1_1; // @[Router.scala 148:38]
  assign input_unit_0_from_1_io_router_resp_vc_sel_1_2 = route_computer_io_resp_0_vc_sel_1_2; // @[Router.scala 148:38]
  assign input_unit_0_from_1_io_router_resp_vc_sel_0_0 = route_computer_io_resp_0_vc_sel_0_0; // @[Router.scala 148:38]
  assign input_unit_0_from_1_io_router_resp_vc_sel_0_1 = route_computer_io_resp_0_vc_sel_0_1; // @[Router.scala 148:38]
  assign input_unit_0_from_1_io_router_resp_vc_sel_0_2 = route_computer_io_resp_0_vc_sel_0_2; // @[Router.scala 148:38]
  assign input_unit_0_from_1_io_router_resp_vc_sel_0_3 = route_computer_io_resp_0_vc_sel_0_3; // @[Router.scala 148:38]
  assign input_unit_0_from_1_io_vcalloc_req_ready = vc_allocator_io_req_0_ready; // @[Router.scala 151:23]
  assign input_unit_0_from_1_io_vcalloc_resp_vc_sel_2_0 = vc_allocator_io_resp_0_vc_sel_2_0; // @[Router.scala 153:39]
  assign input_unit_0_from_1_io_vcalloc_resp_vc_sel_1_0 = vc_allocator_io_resp_0_vc_sel_1_0; // @[Router.scala 153:39]
  assign input_unit_0_from_1_io_vcalloc_resp_vc_sel_1_1 = vc_allocator_io_resp_0_vc_sel_1_1; // @[Router.scala 153:39]
  assign input_unit_0_from_1_io_vcalloc_resp_vc_sel_1_2 = vc_allocator_io_resp_0_vc_sel_1_2; // @[Router.scala 153:39]
  assign input_unit_0_from_1_io_vcalloc_resp_vc_sel_0_0 = vc_allocator_io_resp_0_vc_sel_0_0; // @[Router.scala 153:39]
  assign input_unit_0_from_1_io_vcalloc_resp_vc_sel_0_1 = vc_allocator_io_resp_0_vc_sel_0_1; // @[Router.scala 153:39]
  assign input_unit_0_from_1_io_vcalloc_resp_vc_sel_0_2 = vc_allocator_io_resp_0_vc_sel_0_2; // @[Router.scala 153:39]
  assign input_unit_0_from_1_io_vcalloc_resp_vc_sel_0_3 = vc_allocator_io_resp_0_vc_sel_0_3; // @[Router.scala 153:39]
  assign input_unit_0_from_1_io_out_credit_available_2_0 = egress_unit_2_to_0_io_credit_available_0; // @[Router.scala 162:42]
  assign input_unit_0_from_1_io_out_credit_available_1_0 = output_unit_1_to_3_io_credit_available_0; // @[Router.scala 162:42]
  assign input_unit_0_from_1_io_out_credit_available_1_1 = output_unit_1_to_3_io_credit_available_1; // @[Router.scala 162:42]
  assign input_unit_0_from_1_io_out_credit_available_1_2 = output_unit_1_to_3_io_credit_available_2; // @[Router.scala 162:42]
  assign input_unit_0_from_1_io_out_credit_available_1_3 = output_unit_1_to_3_io_credit_available_3; // @[Router.scala 162:42]
  assign input_unit_0_from_1_io_out_credit_available_0_0 = output_unit_0_to_1_io_credit_available_0; // @[Router.scala 162:42]
  assign input_unit_0_from_1_io_out_credit_available_0_1 = output_unit_0_to_1_io_credit_available_1; // @[Router.scala 162:42]
  assign input_unit_0_from_1_io_out_credit_available_0_2 = output_unit_0_to_1_io_credit_available_2; // @[Router.scala 162:42]
  assign input_unit_0_from_1_io_out_credit_available_0_3 = output_unit_0_to_1_io_credit_available_3; // @[Router.scala 162:42]
  assign input_unit_0_from_1_io_salloc_req_0_ready = switch_allocator_io_req_0_0_ready; // @[Router.scala 165:23]
  assign input_unit_0_from_1_io_in_flit_0_valid = auto_dest_nodes_in_0_flit_0_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_1_io_in_flit_0_bits_head = auto_dest_nodes_in_0_flit_0_bits_head; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_1_io_in_flit_0_bits_tail = auto_dest_nodes_in_0_flit_0_bits_tail; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_1_io_in_flit_0_bits_payload = auto_dest_nodes_in_0_flit_0_bits_payload; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_1_io_in_flit_0_bits_flow_ingress_node = auto_dest_nodes_in_0_flit_0_bits_flow_ingress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_1_io_in_flit_0_bits_flow_egress_node = auto_dest_nodes_in_0_flit_0_bits_flow_egress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_1_io_in_flit_0_bits_virt_channel_id = auto_dest_nodes_in_0_flit_0_bits_virt_channel_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_1_from_3_clock = clock;
  assign input_unit_1_from_3_reset = reset;
  assign input_unit_1_from_3_io_router_resp_vc_sel_1_0 = route_computer_io_resp_1_vc_sel_1_0; // @[Router.scala 148:38]
  assign input_unit_1_from_3_io_router_resp_vc_sel_1_1 = route_computer_io_resp_1_vc_sel_1_1; // @[Router.scala 148:38]
  assign input_unit_1_from_3_io_router_resp_vc_sel_1_2 = route_computer_io_resp_1_vc_sel_1_2; // @[Router.scala 148:38]
  assign input_unit_1_from_3_io_router_resp_vc_sel_0_0 = route_computer_io_resp_1_vc_sel_0_0; // @[Router.scala 148:38]
  assign input_unit_1_from_3_io_router_resp_vc_sel_0_1 = route_computer_io_resp_1_vc_sel_0_1; // @[Router.scala 148:38]
  assign input_unit_1_from_3_io_router_resp_vc_sel_0_2 = route_computer_io_resp_1_vc_sel_0_2; // @[Router.scala 148:38]
  assign input_unit_1_from_3_io_router_resp_vc_sel_0_3 = route_computer_io_resp_1_vc_sel_0_3; // @[Router.scala 148:38]
  assign input_unit_1_from_3_io_vcalloc_req_ready = vc_allocator_io_req_1_ready; // @[Router.scala 151:23]
  assign input_unit_1_from_3_io_vcalloc_resp_vc_sel_2_0 = vc_allocator_io_resp_1_vc_sel_2_0; // @[Router.scala 153:39]
  assign input_unit_1_from_3_io_vcalloc_resp_vc_sel_1_0 = vc_allocator_io_resp_1_vc_sel_1_0; // @[Router.scala 153:39]
  assign input_unit_1_from_3_io_vcalloc_resp_vc_sel_1_1 = vc_allocator_io_resp_1_vc_sel_1_1; // @[Router.scala 153:39]
  assign input_unit_1_from_3_io_vcalloc_resp_vc_sel_1_2 = vc_allocator_io_resp_1_vc_sel_1_2; // @[Router.scala 153:39]
  assign input_unit_1_from_3_io_vcalloc_resp_vc_sel_0_0 = vc_allocator_io_resp_1_vc_sel_0_0; // @[Router.scala 153:39]
  assign input_unit_1_from_3_io_vcalloc_resp_vc_sel_0_1 = vc_allocator_io_resp_1_vc_sel_0_1; // @[Router.scala 153:39]
  assign input_unit_1_from_3_io_vcalloc_resp_vc_sel_0_2 = vc_allocator_io_resp_1_vc_sel_0_2; // @[Router.scala 153:39]
  assign input_unit_1_from_3_io_vcalloc_resp_vc_sel_0_3 = vc_allocator_io_resp_1_vc_sel_0_3; // @[Router.scala 153:39]
  assign input_unit_1_from_3_io_out_credit_available_2_0 = egress_unit_2_to_0_io_credit_available_0; // @[Router.scala 162:42]
  assign input_unit_1_from_3_io_out_credit_available_1_0 = output_unit_1_to_3_io_credit_available_0; // @[Router.scala 162:42]
  assign input_unit_1_from_3_io_out_credit_available_1_1 = output_unit_1_to_3_io_credit_available_1; // @[Router.scala 162:42]
  assign input_unit_1_from_3_io_out_credit_available_1_2 = output_unit_1_to_3_io_credit_available_2; // @[Router.scala 162:42]
  assign input_unit_1_from_3_io_out_credit_available_1_3 = output_unit_1_to_3_io_credit_available_3; // @[Router.scala 162:42]
  assign input_unit_1_from_3_io_out_credit_available_0_0 = output_unit_0_to_1_io_credit_available_0; // @[Router.scala 162:42]
  assign input_unit_1_from_3_io_out_credit_available_0_1 = output_unit_0_to_1_io_credit_available_1; // @[Router.scala 162:42]
  assign input_unit_1_from_3_io_out_credit_available_0_2 = output_unit_0_to_1_io_credit_available_2; // @[Router.scala 162:42]
  assign input_unit_1_from_3_io_out_credit_available_0_3 = output_unit_0_to_1_io_credit_available_3; // @[Router.scala 162:42]
  assign input_unit_1_from_3_io_salloc_req_0_ready = switch_allocator_io_req_1_0_ready; // @[Router.scala 165:23]
  assign input_unit_1_from_3_io_in_flit_0_valid = auto_dest_nodes_in_1_flit_0_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_1_from_3_io_in_flit_0_bits_head = auto_dest_nodes_in_1_flit_0_bits_head; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_1_from_3_io_in_flit_0_bits_tail = auto_dest_nodes_in_1_flit_0_bits_tail; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_1_from_3_io_in_flit_0_bits_payload = auto_dest_nodes_in_1_flit_0_bits_payload; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_1_from_3_io_in_flit_0_bits_flow_ingress_node = auto_dest_nodes_in_1_flit_0_bits_flow_ingress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_1_from_3_io_in_flit_0_bits_flow_egress_node = auto_dest_nodes_in_1_flit_0_bits_flow_egress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_1_from_3_io_in_flit_0_bits_virt_channel_id = auto_dest_nodes_in_1_flit_0_bits_virt_channel_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign ingress_unit_2_from_0_clock = clock;
  assign ingress_unit_2_from_0_reset = reset;
  assign ingress_unit_2_from_0_io_router_resp_vc_sel_1_0 = route_computer_io_resp_2_vc_sel_1_0; // @[Router.scala 148:38]
  assign ingress_unit_2_from_0_io_router_resp_vc_sel_1_1 = route_computer_io_resp_2_vc_sel_1_1; // @[Router.scala 148:38]
  assign ingress_unit_2_from_0_io_router_resp_vc_sel_1_2 = route_computer_io_resp_2_vc_sel_1_2; // @[Router.scala 148:38]
  assign ingress_unit_2_from_0_io_router_resp_vc_sel_1_3 = route_computer_io_resp_2_vc_sel_1_3; // @[Router.scala 148:38]
  assign ingress_unit_2_from_0_io_router_resp_vc_sel_0_0 = route_computer_io_resp_2_vc_sel_0_0; // @[Router.scala 148:38]
  assign ingress_unit_2_from_0_io_router_resp_vc_sel_0_1 = route_computer_io_resp_2_vc_sel_0_1; // @[Router.scala 148:38]
  assign ingress_unit_2_from_0_io_router_resp_vc_sel_0_2 = route_computer_io_resp_2_vc_sel_0_2; // @[Router.scala 148:38]
  assign ingress_unit_2_from_0_io_router_resp_vc_sel_0_3 = route_computer_io_resp_2_vc_sel_0_3; // @[Router.scala 148:38]
  assign ingress_unit_2_from_0_io_vcalloc_req_ready = vc_allocator_io_req_2_ready; // @[Router.scala 151:23]
  assign ingress_unit_2_from_0_io_vcalloc_resp_vc_sel_2_0 = vc_allocator_io_resp_2_vc_sel_2_0; // @[Router.scala 153:39]
  assign ingress_unit_2_from_0_io_vcalloc_resp_vc_sel_1_0 = vc_allocator_io_resp_2_vc_sel_1_0; // @[Router.scala 153:39]
  assign ingress_unit_2_from_0_io_vcalloc_resp_vc_sel_1_1 = vc_allocator_io_resp_2_vc_sel_1_1; // @[Router.scala 153:39]
  assign ingress_unit_2_from_0_io_vcalloc_resp_vc_sel_1_2 = vc_allocator_io_resp_2_vc_sel_1_2; // @[Router.scala 153:39]
  assign ingress_unit_2_from_0_io_vcalloc_resp_vc_sel_1_3 = vc_allocator_io_resp_2_vc_sel_1_3; // @[Router.scala 153:39]
  assign ingress_unit_2_from_0_io_vcalloc_resp_vc_sel_0_0 = vc_allocator_io_resp_2_vc_sel_0_0; // @[Router.scala 153:39]
  assign ingress_unit_2_from_0_io_vcalloc_resp_vc_sel_0_1 = vc_allocator_io_resp_2_vc_sel_0_1; // @[Router.scala 153:39]
  assign ingress_unit_2_from_0_io_vcalloc_resp_vc_sel_0_2 = vc_allocator_io_resp_2_vc_sel_0_2; // @[Router.scala 153:39]
  assign ingress_unit_2_from_0_io_vcalloc_resp_vc_sel_0_3 = vc_allocator_io_resp_2_vc_sel_0_3; // @[Router.scala 153:39]
  assign ingress_unit_2_from_0_io_out_credit_available_2_0 = egress_unit_2_to_0_io_credit_available_0; // @[Router.scala 162:42]
  assign ingress_unit_2_from_0_io_out_credit_available_1_0 = output_unit_1_to_3_io_credit_available_0; // @[Router.scala 162:42]
  assign ingress_unit_2_from_0_io_out_credit_available_1_1 = output_unit_1_to_3_io_credit_available_1; // @[Router.scala 162:42]
  assign ingress_unit_2_from_0_io_out_credit_available_1_2 = output_unit_1_to_3_io_credit_available_2; // @[Router.scala 162:42]
  assign ingress_unit_2_from_0_io_out_credit_available_1_3 = output_unit_1_to_3_io_credit_available_3; // @[Router.scala 162:42]
  assign ingress_unit_2_from_0_io_out_credit_available_0_0 = output_unit_0_to_1_io_credit_available_0; // @[Router.scala 162:42]
  assign ingress_unit_2_from_0_io_out_credit_available_0_1 = output_unit_0_to_1_io_credit_available_1; // @[Router.scala 162:42]
  assign ingress_unit_2_from_0_io_out_credit_available_0_2 = output_unit_0_to_1_io_credit_available_2; // @[Router.scala 162:42]
  assign ingress_unit_2_from_0_io_out_credit_available_0_3 = output_unit_0_to_1_io_credit_available_3; // @[Router.scala 162:42]
  assign ingress_unit_2_from_0_io_salloc_req_0_ready = switch_allocator_io_req_2_0_ready; // @[Router.scala 165:23]
  assign ingress_unit_2_from_0_io_in_valid = auto_ingress_nodes_in_flit_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign ingress_unit_2_from_0_io_in_bits_head = auto_ingress_nodes_in_flit_bits_head; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign ingress_unit_2_from_0_io_in_bits_tail = auto_ingress_nodes_in_flit_bits_tail; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign ingress_unit_2_from_0_io_in_bits_payload = auto_ingress_nodes_in_flit_bits_payload; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign ingress_unit_2_from_0_io_in_bits_egress_id = auto_ingress_nodes_in_flit_bits_egress_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign output_unit_0_to_1_clock = clock;
  assign output_unit_0_to_1_reset = reset;
  assign output_unit_0_to_1_io_in_0_valid = switch_io_out_0_0_valid; // @[Router.scala 172:29]
  assign output_unit_0_to_1_io_in_0_bits_head = switch_io_out_0_0_bits_head; // @[Router.scala 172:29]
  assign output_unit_0_to_1_io_in_0_bits_tail = switch_io_out_0_0_bits_tail; // @[Router.scala 172:29]
  assign output_unit_0_to_1_io_in_0_bits_payload = switch_io_out_0_0_bits_payload; // @[Router.scala 172:29]
  assign output_unit_0_to_1_io_in_0_bits_flow_ingress_node = switch_io_out_0_0_bits_flow_ingress_node; // @[Router.scala 172:29]
  assign output_unit_0_to_1_io_in_0_bits_flow_egress_node = switch_io_out_0_0_bits_flow_egress_node; // @[Router.scala 172:29]
  assign output_unit_0_to_1_io_in_0_bits_virt_channel_id = switch_io_out_0_0_bits_virt_channel_id; // @[Router.scala 172:29]
  assign output_unit_0_to_1_io_allocs_0_alloc = vc_allocator_io_out_allocs_0_0_alloc; // @[Router.scala 157:33]
  assign output_unit_0_to_1_io_allocs_1_alloc = vc_allocator_io_out_allocs_0_1_alloc; // @[Router.scala 157:33]
  assign output_unit_0_to_1_io_allocs_2_alloc = vc_allocator_io_out_allocs_0_2_alloc; // @[Router.scala 157:33]
  assign output_unit_0_to_1_io_allocs_3_alloc = vc_allocator_io_out_allocs_0_3_alloc; // @[Router.scala 157:33]
  assign output_unit_0_to_1_io_credit_alloc_0_alloc = switch_allocator_io_credit_alloc_0_0_alloc; // @[Router.scala 167:39]
  assign output_unit_0_to_1_io_credit_alloc_1_alloc = switch_allocator_io_credit_alloc_0_1_alloc; // @[Router.scala 167:39]
  assign output_unit_0_to_1_io_credit_alloc_2_alloc = switch_allocator_io_credit_alloc_0_2_alloc; // @[Router.scala 167:39]
  assign output_unit_0_to_1_io_credit_alloc_3_alloc = switch_allocator_io_credit_alloc_0_3_alloc; // @[Router.scala 167:39]
  assign output_unit_0_to_1_io_out_credit_return = auto_source_nodes_out_0_credit_return; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign output_unit_0_to_1_io_out_vc_free = auto_source_nodes_out_0_vc_free; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign output_unit_1_to_3_clock = clock;
  assign output_unit_1_to_3_reset = reset;
  assign output_unit_1_to_3_io_in_0_valid = switch_io_out_1_0_valid; // @[Router.scala 172:29]
  assign output_unit_1_to_3_io_in_0_bits_head = switch_io_out_1_0_bits_head; // @[Router.scala 172:29]
  assign output_unit_1_to_3_io_in_0_bits_tail = switch_io_out_1_0_bits_tail; // @[Router.scala 172:29]
  assign output_unit_1_to_3_io_in_0_bits_payload = switch_io_out_1_0_bits_payload; // @[Router.scala 172:29]
  assign output_unit_1_to_3_io_in_0_bits_flow_ingress_node = switch_io_out_1_0_bits_flow_ingress_node; // @[Router.scala 172:29]
  assign output_unit_1_to_3_io_in_0_bits_flow_egress_node = switch_io_out_1_0_bits_flow_egress_node; // @[Router.scala 172:29]
  assign output_unit_1_to_3_io_in_0_bits_virt_channel_id = switch_io_out_1_0_bits_virt_channel_id; // @[Router.scala 172:29]
  assign output_unit_1_to_3_io_allocs_0_alloc = vc_allocator_io_out_allocs_1_0_alloc; // @[Router.scala 157:33]
  assign output_unit_1_to_3_io_allocs_1_alloc = vc_allocator_io_out_allocs_1_1_alloc; // @[Router.scala 157:33]
  assign output_unit_1_to_3_io_allocs_2_alloc = vc_allocator_io_out_allocs_1_2_alloc; // @[Router.scala 157:33]
  assign output_unit_1_to_3_io_allocs_3_alloc = vc_allocator_io_out_allocs_1_3_alloc; // @[Router.scala 157:33]
  assign output_unit_1_to_3_io_credit_alloc_0_alloc = switch_allocator_io_credit_alloc_1_0_alloc; // @[Router.scala 167:39]
  assign output_unit_1_to_3_io_credit_alloc_1_alloc = switch_allocator_io_credit_alloc_1_1_alloc; // @[Router.scala 167:39]
  assign output_unit_1_to_3_io_credit_alloc_2_alloc = switch_allocator_io_credit_alloc_1_2_alloc; // @[Router.scala 167:39]
  assign output_unit_1_to_3_io_credit_alloc_3_alloc = switch_allocator_io_credit_alloc_1_3_alloc; // @[Router.scala 167:39]
  assign output_unit_1_to_3_io_out_credit_return = auto_source_nodes_out_1_credit_return; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign output_unit_1_to_3_io_out_vc_free = auto_source_nodes_out_1_vc_free; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign egress_unit_2_to_0_clock = clock;
  assign egress_unit_2_to_0_reset = reset;
  assign egress_unit_2_to_0_io_in_0_valid = switch_io_out_2_0_valid; // @[Router.scala 172:29]
  assign egress_unit_2_to_0_io_in_0_bits_head = switch_io_out_2_0_bits_head; // @[Router.scala 172:29]
  assign egress_unit_2_to_0_io_in_0_bits_tail = switch_io_out_2_0_bits_tail; // @[Router.scala 172:29]
  assign egress_unit_2_to_0_io_in_0_bits_payload = switch_io_out_2_0_bits_payload; // @[Router.scala 172:29]
  assign egress_unit_2_to_0_io_in_0_bits_flow_ingress_node = switch_io_out_2_0_bits_flow_ingress_node; // @[Router.scala 172:29]
  assign egress_unit_2_to_0_io_allocs_0_alloc = vc_allocator_io_out_allocs_2_0_alloc; // @[Router.scala 157:33]
  assign egress_unit_2_to_0_io_credit_alloc_0_alloc = switch_allocator_io_credit_alloc_2_0_alloc; // @[Router.scala 167:39]
  assign egress_unit_2_to_0_io_credit_alloc_0_tail = switch_allocator_io_credit_alloc_2_0_tail; // @[Router.scala 167:39]
  assign switch_clock = clock;
  assign switch_reset = reset;
  assign switch_io_in_2_0_valid = ingress_unit_2_from_0_io_out_0_valid; // @[Router.scala 170:23]
  assign switch_io_in_2_0_bits_flit_head = ingress_unit_2_from_0_io_out_0_bits_flit_head; // @[Router.scala 170:23]
  assign switch_io_in_2_0_bits_flit_tail = ingress_unit_2_from_0_io_out_0_bits_flit_tail; // @[Router.scala 170:23]
  assign switch_io_in_2_0_bits_flit_payload = ingress_unit_2_from_0_io_out_0_bits_flit_payload; // @[Router.scala 170:23]
  assign switch_io_in_2_0_bits_flit_flow_ingress_node = ingress_unit_2_from_0_io_out_0_bits_flit_flow_ingress_node; // @[Router.scala 170:23]
  assign switch_io_in_2_0_bits_flit_flow_egress_node = ingress_unit_2_from_0_io_out_0_bits_flit_flow_egress_node; // @[Router.scala 170:23]
  assign switch_io_in_2_0_bits_out_virt_channel = ingress_unit_2_from_0_io_out_0_bits_out_virt_channel; // @[Router.scala 170:23]
  assign switch_io_in_1_0_valid = input_unit_1_from_3_io_out_0_valid; // @[Router.scala 170:23]
  assign switch_io_in_1_0_bits_flit_head = input_unit_1_from_3_io_out_0_bits_flit_head; // @[Router.scala 170:23]
  assign switch_io_in_1_0_bits_flit_tail = input_unit_1_from_3_io_out_0_bits_flit_tail; // @[Router.scala 170:23]
  assign switch_io_in_1_0_bits_flit_payload = input_unit_1_from_3_io_out_0_bits_flit_payload; // @[Router.scala 170:23]
  assign switch_io_in_1_0_bits_flit_flow_ingress_node = input_unit_1_from_3_io_out_0_bits_flit_flow_ingress_node; // @[Router.scala 170:23]
  assign switch_io_in_1_0_bits_flit_flow_egress_node = input_unit_1_from_3_io_out_0_bits_flit_flow_egress_node; // @[Router.scala 170:23]
  assign switch_io_in_1_0_bits_out_virt_channel = input_unit_1_from_3_io_out_0_bits_out_virt_channel; // @[Router.scala 170:23]
  assign switch_io_in_0_0_valid = input_unit_0_from_1_io_out_0_valid; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_head = input_unit_0_from_1_io_out_0_bits_flit_head; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_tail = input_unit_0_from_1_io_out_0_bits_flit_tail; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_payload = input_unit_0_from_1_io_out_0_bits_flit_payload; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_flow_ingress_node = input_unit_0_from_1_io_out_0_bits_flit_flow_ingress_node; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_flow_egress_node = input_unit_0_from_1_io_out_0_bits_flit_flow_egress_node; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_out_virt_channel = input_unit_0_from_1_io_out_0_bits_out_virt_channel; // @[Router.scala 170:23]
  assign switch_io_sel_2_0_2_0 = switch_io_sel_REG_2_0_2_0; // @[Router.scala 173:19]
  assign switch_io_sel_2_0_1_0 = switch_io_sel_REG_2_0_1_0; // @[Router.scala 173:19]
  assign switch_io_sel_2_0_0_0 = switch_io_sel_REG_2_0_0_0; // @[Router.scala 173:19]
  assign switch_io_sel_1_0_2_0 = switch_io_sel_REG_1_0_2_0; // @[Router.scala 173:19]
  assign switch_io_sel_1_0_1_0 = switch_io_sel_REG_1_0_1_0; // @[Router.scala 173:19]
  assign switch_io_sel_1_0_0_0 = switch_io_sel_REG_1_0_0_0; // @[Router.scala 173:19]
  assign switch_io_sel_0_0_2_0 = switch_io_sel_REG_0_0_2_0; // @[Router.scala 173:19]
  assign switch_io_sel_0_0_1_0 = switch_io_sel_REG_0_0_1_0; // @[Router.scala 173:19]
  assign switch_io_sel_0_0_0_0 = switch_io_sel_REG_0_0_0_0; // @[Router.scala 173:19]
  assign switch_allocator_clock = clock;
  assign switch_allocator_reset = reset;
  assign switch_allocator_io_req_2_0_valid = ingress_unit_2_from_0_io_salloc_req_0_valid; // @[Router.scala 165:23]
  assign switch_allocator_io_req_2_0_bits_vc_sel_2_0 = ingress_unit_2_from_0_io_salloc_req_0_bits_vc_sel_2_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_2_0_bits_vc_sel_1_0 = ingress_unit_2_from_0_io_salloc_req_0_bits_vc_sel_1_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_2_0_bits_vc_sel_1_1 = ingress_unit_2_from_0_io_salloc_req_0_bits_vc_sel_1_1; // @[Router.scala 165:23]
  assign switch_allocator_io_req_2_0_bits_vc_sel_1_2 = ingress_unit_2_from_0_io_salloc_req_0_bits_vc_sel_1_2; // @[Router.scala 165:23]
  assign switch_allocator_io_req_2_0_bits_vc_sel_1_3 = ingress_unit_2_from_0_io_salloc_req_0_bits_vc_sel_1_3; // @[Router.scala 165:23]
  assign switch_allocator_io_req_2_0_bits_vc_sel_0_0 = ingress_unit_2_from_0_io_salloc_req_0_bits_vc_sel_0_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_2_0_bits_vc_sel_0_1 = ingress_unit_2_from_0_io_salloc_req_0_bits_vc_sel_0_1; // @[Router.scala 165:23]
  assign switch_allocator_io_req_2_0_bits_vc_sel_0_2 = ingress_unit_2_from_0_io_salloc_req_0_bits_vc_sel_0_2; // @[Router.scala 165:23]
  assign switch_allocator_io_req_2_0_bits_vc_sel_0_3 = ingress_unit_2_from_0_io_salloc_req_0_bits_vc_sel_0_3; // @[Router.scala 165:23]
  assign switch_allocator_io_req_2_0_bits_tail = ingress_unit_2_from_0_io_salloc_req_0_bits_tail; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_valid = input_unit_1_from_3_io_salloc_req_0_valid; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_vc_sel_2_0 = input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_2_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_vc_sel_1_0 = input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_1_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_vc_sel_1_1 = input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_1_1; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_vc_sel_1_2 = input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_1_2; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_vc_sel_1_3 = input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_1_3; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_vc_sel_0_0 = input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_0_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_vc_sel_0_1 = input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_0_1; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_vc_sel_0_2 = input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_0_2; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_vc_sel_0_3 = input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_0_3; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_tail = input_unit_1_from_3_io_salloc_req_0_bits_tail; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_valid = input_unit_0_from_1_io_salloc_req_0_valid; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_2_0 = input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_2_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_1_0 = input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_1_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_1_1 = input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_1_1; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_1_2 = input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_1_2; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_1_3 = input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_1_3; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_0_0 = input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_0_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_0_1 = input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_0_1; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_0_2 = input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_0_2; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_0_3 = input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_0_3; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_tail = input_unit_0_from_1_io_salloc_req_0_bits_tail; // @[Router.scala 165:23]
  assign vc_allocator_clock = clock;
  assign vc_allocator_reset = reset;
  assign vc_allocator_io_req_2_valid = ingress_unit_2_from_0_io_vcalloc_req_valid; // @[Router.scala 151:23]
  assign vc_allocator_io_req_2_bits_vc_sel_2_0 = ingress_unit_2_from_0_io_vcalloc_req_bits_vc_sel_2_0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_2_bits_vc_sel_1_0 = ingress_unit_2_from_0_io_vcalloc_req_bits_vc_sel_1_0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_2_bits_vc_sel_1_1 = ingress_unit_2_from_0_io_vcalloc_req_bits_vc_sel_1_1; // @[Router.scala 151:23]
  assign vc_allocator_io_req_2_bits_vc_sel_1_2 = ingress_unit_2_from_0_io_vcalloc_req_bits_vc_sel_1_2; // @[Router.scala 151:23]
  assign vc_allocator_io_req_2_bits_vc_sel_1_3 = ingress_unit_2_from_0_io_vcalloc_req_bits_vc_sel_1_3; // @[Router.scala 151:23]
  assign vc_allocator_io_req_2_bits_vc_sel_0_0 = ingress_unit_2_from_0_io_vcalloc_req_bits_vc_sel_0_0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_2_bits_vc_sel_0_1 = ingress_unit_2_from_0_io_vcalloc_req_bits_vc_sel_0_1; // @[Router.scala 151:23]
  assign vc_allocator_io_req_2_bits_vc_sel_0_2 = ingress_unit_2_from_0_io_vcalloc_req_bits_vc_sel_0_2; // @[Router.scala 151:23]
  assign vc_allocator_io_req_2_bits_vc_sel_0_3 = ingress_unit_2_from_0_io_vcalloc_req_bits_vc_sel_0_3; // @[Router.scala 151:23]
  assign vc_allocator_io_req_1_valid = input_unit_1_from_3_io_vcalloc_req_valid; // @[Router.scala 151:23]
  assign vc_allocator_io_req_1_bits_vc_sel_2_0 = input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_2_0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_1_bits_vc_sel_1_0 = input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_1_0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_1_bits_vc_sel_1_1 = input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_1_1; // @[Router.scala 151:23]
  assign vc_allocator_io_req_1_bits_vc_sel_1_2 = input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_1_2; // @[Router.scala 151:23]
  assign vc_allocator_io_req_1_bits_vc_sel_1_3 = 1'h0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_1_bits_vc_sel_0_0 = input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_0_0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_1_bits_vc_sel_0_1 = input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_0_1; // @[Router.scala 151:23]
  assign vc_allocator_io_req_1_bits_vc_sel_0_2 = input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_0_2; // @[Router.scala 151:23]
  assign vc_allocator_io_req_1_bits_vc_sel_0_3 = input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_0_3; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_valid = input_unit_0_from_1_io_vcalloc_req_valid; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_2_0 = input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_2_0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_1_0 = input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_1_0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_1_1 = input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_1_1; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_1_2 = input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_1_2; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_1_3 = 1'h0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_0_0 = input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_0_0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_0_1 = input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_0_1; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_0_2 = input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_0_2; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_0_3 = input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_0_3; // @[Router.scala 151:23]
  assign vc_allocator_io_channel_status_2_0_occupied = egress_unit_2_to_0_io_channel_status_0_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_1_0_occupied = output_unit_1_to_3_io_channel_status_0_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_1_1_occupied = output_unit_1_to_3_io_channel_status_1_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_1_2_occupied = output_unit_1_to_3_io_channel_status_2_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_1_3_occupied = output_unit_1_to_3_io_channel_status_3_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_0_0_occupied = output_unit_0_to_1_io_channel_status_0_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_0_1_occupied = output_unit_0_to_1_io_channel_status_1_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_0_2_occupied = output_unit_0_to_1_io_channel_status_2_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_0_3_occupied = output_unit_0_to_1_io_channel_status_3_occupied; // @[Router.scala 159:23]
  assign route_computer_io_req_2_bits_flow_ingress_node = ingress_unit_2_from_0_io_router_req_bits_flow_ingress_node; // @[Router.scala 146:23]
  assign route_computer_io_req_2_bits_flow_egress_node = ingress_unit_2_from_0_io_router_req_bits_flow_egress_node; // @[Router.scala 146:23]
  assign route_computer_io_req_1_bits_src_virt_id = input_unit_1_from_3_io_router_req_bits_src_virt_id; // @[Router.scala 146:23]
  assign route_computer_io_req_1_bits_flow_ingress_node = input_unit_1_from_3_io_router_req_bits_flow_ingress_node; // @[Router.scala 146:23]
  assign route_computer_io_req_1_bits_flow_egress_node = input_unit_1_from_3_io_router_req_bits_flow_egress_node; // @[Router.scala 146:23]
  assign route_computer_io_req_0_bits_src_virt_id = input_unit_0_from_1_io_router_req_bits_src_virt_id; // @[Router.scala 146:23]
  assign route_computer_io_req_0_bits_flow_ingress_node = input_unit_0_from_1_io_router_req_bits_flow_ingress_node; // @[Router.scala 146:23]
  assign route_computer_io_req_0_bits_flow_egress_node = input_unit_0_from_1_io_router_req_bits_flow_egress_node; // @[Router.scala 146:23]
  always @(posedge clock) begin
    switch_io_sel_REG_2_0_2_0 <= switch_allocator_io_switch_sel_2_0_2_0; // @[Router.scala 176:14]
    switch_io_sel_REG_2_0_1_0 <= switch_allocator_io_switch_sel_2_0_1_0; // @[Router.scala 176:14]
    switch_io_sel_REG_2_0_0_0 <= switch_allocator_io_switch_sel_2_0_0_0; // @[Router.scala 176:14]
    switch_io_sel_REG_1_0_2_0 <= switch_allocator_io_switch_sel_1_0_2_0; // @[Router.scala 176:14]
    switch_io_sel_REG_1_0_1_0 <= switch_allocator_io_switch_sel_1_0_1_0; // @[Router.scala 176:14]
    switch_io_sel_REG_1_0_0_0 <= switch_allocator_io_switch_sel_1_0_0_0; // @[Router.scala 176:14]
    switch_io_sel_REG_0_0_2_0 <= switch_allocator_io_switch_sel_0_0_2_0; // @[Router.scala 176:14]
    switch_io_sel_REG_0_0_1_0 <= switch_allocator_io_switch_sel_0_0_1_0; // @[Router.scala 176:14]
    switch_io_sel_REG_0_0_0_0 <= switch_allocator_io_switch_sel_0_0_0_0; // @[Router.scala 176:14]
    if (reset) begin // @[Router.scala 193:28]
      debug_tsc <= 64'h0; // @[Router.scala 193:28]
    end else begin
      debug_tsc <= _debug_tsc_T_1; // @[Router.scala 194:15]
    end
    if (reset) begin // @[Router.scala 195:31]
      debug_sample <= 64'h0; // @[Router.scala 195:31]
    end else if (debug_sample == _GEN_6) begin // @[Router.scala 198:47]
      debug_sample <= 64'h0; // @[Router.scala 198:62]
    end else begin
      debug_sample <= _debug_sample_T_1; // @[Router.scala 196:18]
    end
    if (reset) begin // @[Router.scala 201:29]
      util_ctr <= 64'h0; // @[Router.scala 201:29]
    end else begin
      util_ctr <= _util_ctr_T_1; // @[Router.scala 203:16]
    end
    if (reset) begin // @[Router.scala 202:26]
      fired <= 1'h0; // @[Router.scala 202:26]
    end else if (plusarg_reader_out != 20'h0 & _T_2 & fired) begin // @[Router.scala 205:81]
      fired <= auto_dest_nodes_in_0_flit_0_valid; // @[Router.scala 208:15]
    end else begin
      fired <= fired | auto_dest_nodes_in_0_flit_0_valid; // @[Router.scala 204:13]
    end
    if (reset) begin // @[Router.scala 201:29]
      util_ctr_1 <= 64'h0; // @[Router.scala 201:29]
    end else begin
      util_ctr_1 <= _util_ctr_T_3; // @[Router.scala 203:16]
    end
    if (reset) begin // @[Router.scala 202:26]
      fired_1 <= 1'h0; // @[Router.scala 202:26]
    end else if (plusarg_reader_out != 20'h0 & _T_2 & fired_1) begin // @[Router.scala 205:81]
      fired_1 <= auto_dest_nodes_in_1_flit_0_valid; // @[Router.scala 208:15]
    end else begin
      fired_1 <= fired_1 | auto_dest_nodes_in_1_flit_0_valid; // @[Router.scala 204:13]
    end
    if (reset) begin // @[Router.scala 201:29]
      util_ctr_2 <= 64'h0; // @[Router.scala 201:29]
    end else begin
      util_ctr_2 <= _util_ctr_T_5; // @[Router.scala 203:16]
    end
    if (reset) begin // @[Router.scala 202:26]
      fired_2 <= 1'h0; // @[Router.scala 202:26]
    end else if (plusarg_reader_out != 20'h0 & _T_2 & fired_2) begin // @[Router.scala 205:81]
      fired_2 <= _T_19; // @[Router.scala 208:15]
    end else begin
      fired_2 <= fired_2 | _T_19; // @[Router.scala 204:13]
    end
    if (reset) begin // @[Router.scala 201:29]
      util_ctr_3 <= 64'h0; // @[Router.scala 201:29]
    end else begin
      util_ctr_3 <= _util_ctr_T_7; // @[Router.scala 203:16]
    end
    if (reset) begin // @[Router.scala 202:26]
      fired_3 <= 1'h0; // @[Router.scala 202:26]
    end else if (plusarg_reader_out != 20'h0 & _T_2 & fired_3) begin // @[Router.scala 205:81]
      fired_3 <= x1_2_flit_valid; // @[Router.scala 208:15]
    end else begin
      fired_3 <= fired_3 | x1_2_flit_valid; // @[Router.scala 204:13]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8 & ~reset) begin
          $fwrite(32'h80000002,"nocsample %d 1 0 %d\n",debug_tsc,util_ctr); // @[Router.scala 207:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_16 & ~reset) begin
          $fwrite(32'h80000002,"nocsample %d 3 0 %d\n",debug_tsc,util_ctr_1); // @[Router.scala 207:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_25 & ~reset) begin
          $fwrite(32'h80000002,"nocsample %d i0 0 %d\n",debug_tsc,util_ctr_2); // @[Router.scala 207:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_34 & ~reset) begin
          $fwrite(32'h80000002,"nocsample %d 0 e0 %d\n",debug_tsc,util_ctr_3); // @[Router.scala 207:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  switch_io_sel_REG_2_0_2_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  switch_io_sel_REG_2_0_1_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  switch_io_sel_REG_2_0_0_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  switch_io_sel_REG_1_0_2_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  switch_io_sel_REG_1_0_1_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  switch_io_sel_REG_1_0_0_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  switch_io_sel_REG_0_0_2_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  switch_io_sel_REG_0_0_1_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  switch_io_sel_REG_0_0_0_0 = _RAND_8[0:0];
  _RAND_9 = {2{`RANDOM}};
  debug_tsc = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  debug_sample = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  util_ctr = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  fired = _RAND_12[0:0];
  _RAND_13 = {2{`RANDOM}};
  util_ctr_1 = _RAND_13[63:0];
  _RAND_14 = {1{`RANDOM}};
  fired_1 = _RAND_14[0:0];
  _RAND_15 = {2{`RANDOM}};
  util_ctr_2 = _RAND_15[63:0];
  _RAND_16 = {1{`RANDOM}};
  fired_2 = _RAND_16[0:0];
  _RAND_17 = {2{`RANDOM}};
  util_ctr_3 = _RAND_17[63:0];
  _RAND_18 = {1{`RANDOM}};
  fired_3 = _RAND_18[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ClockSinkDomain(
  output [1:0]  auto_routers_debug_out_va_stall_0,
  output [1:0]  auto_routers_debug_out_va_stall_1,
  output [1:0]  auto_routers_debug_out_sa_stall_0,
  output [1:0]  auto_routers_debug_out_sa_stall_1,
  output        auto_routers_egress_nodes_out_flit_valid,
  output        auto_routers_egress_nodes_out_flit_bits_head,
  output        auto_routers_egress_nodes_out_flit_bits_tail,
  output [63:0] auto_routers_egress_nodes_out_flit_bits_payload,
  output [1:0]  auto_routers_egress_nodes_out_flit_bits_ingress_id,
  output        auto_routers_ingress_nodes_in_flit_ready,
  input         auto_routers_ingress_nodes_in_flit_valid,
  input         auto_routers_ingress_nodes_in_flit_bits_head,
  input         auto_routers_ingress_nodes_in_flit_bits_tail,
  input  [63:0] auto_routers_ingress_nodes_in_flit_bits_payload,
  input  [1:0]  auto_routers_ingress_nodes_in_flit_bits_egress_id,
  output        auto_routers_source_nodes_out_1_flit_0_valid,
  output        auto_routers_source_nodes_out_1_flit_0_bits_head,
  output        auto_routers_source_nodes_out_1_flit_0_bits_tail,
  output [63:0] auto_routers_source_nodes_out_1_flit_0_bits_payload,
  output [1:0]  auto_routers_source_nodes_out_1_flit_0_bits_flow_ingress_node,
  output [1:0]  auto_routers_source_nodes_out_1_flit_0_bits_flow_egress_node,
  output [1:0]  auto_routers_source_nodes_out_1_flit_0_bits_virt_channel_id,
  input  [3:0]  auto_routers_source_nodes_out_1_credit_return,
  input  [3:0]  auto_routers_source_nodes_out_1_vc_free,
  output        auto_routers_source_nodes_out_0_flit_0_valid,
  output        auto_routers_source_nodes_out_0_flit_0_bits_head,
  output        auto_routers_source_nodes_out_0_flit_0_bits_tail,
  output [63:0] auto_routers_source_nodes_out_0_flit_0_bits_payload,
  output [1:0]  auto_routers_source_nodes_out_0_flit_0_bits_flow_ingress_node,
  output [1:0]  auto_routers_source_nodes_out_0_flit_0_bits_flow_egress_node,
  output [1:0]  auto_routers_source_nodes_out_0_flit_0_bits_virt_channel_id,
  input  [3:0]  auto_routers_source_nodes_out_0_credit_return,
  input  [3:0]  auto_routers_source_nodes_out_0_vc_free,
  input         auto_routers_dest_nodes_in_1_flit_0_valid,
  input         auto_routers_dest_nodes_in_1_flit_0_bits_head,
  input         auto_routers_dest_nodes_in_1_flit_0_bits_tail,
  input  [63:0] auto_routers_dest_nodes_in_1_flit_0_bits_payload,
  input  [1:0]  auto_routers_dest_nodes_in_1_flit_0_bits_flow_ingress_node,
  input  [1:0]  auto_routers_dest_nodes_in_1_flit_0_bits_flow_egress_node,
  input  [1:0]  auto_routers_dest_nodes_in_1_flit_0_bits_virt_channel_id,
  output [3:0]  auto_routers_dest_nodes_in_1_credit_return,
  output [3:0]  auto_routers_dest_nodes_in_1_vc_free,
  input         auto_routers_dest_nodes_in_0_flit_0_valid,
  input         auto_routers_dest_nodes_in_0_flit_0_bits_head,
  input         auto_routers_dest_nodes_in_0_flit_0_bits_tail,
  input  [63:0] auto_routers_dest_nodes_in_0_flit_0_bits_payload,
  input  [1:0]  auto_routers_dest_nodes_in_0_flit_0_bits_flow_ingress_node,
  input  [1:0]  auto_routers_dest_nodes_in_0_flit_0_bits_flow_egress_node,
  input  [1:0]  auto_routers_dest_nodes_in_0_flit_0_bits_virt_channel_id,
  output [3:0]  auto_routers_dest_nodes_in_0_credit_return,
  output [3:0]  auto_routers_dest_nodes_in_0_vc_free,
  input         auto_clock_in_clock,
  input         auto_clock_in_reset
);
  wire  routers_clock; // @[NoC.scala 64:22]
  wire  routers_reset; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_debug_out_va_stall_0; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_debug_out_va_stall_1; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_debug_out_sa_stall_0; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_debug_out_sa_stall_1; // @[NoC.scala 64:22]
  wire  routers_auto_egress_nodes_out_flit_valid; // @[NoC.scala 64:22]
  wire  routers_auto_egress_nodes_out_flit_bits_head; // @[NoC.scala 64:22]
  wire  routers_auto_egress_nodes_out_flit_bits_tail; // @[NoC.scala 64:22]
  wire [63:0] routers_auto_egress_nodes_out_flit_bits_payload; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_egress_nodes_out_flit_bits_ingress_id; // @[NoC.scala 64:22]
  wire  routers_auto_ingress_nodes_in_flit_ready; // @[NoC.scala 64:22]
  wire  routers_auto_ingress_nodes_in_flit_valid; // @[NoC.scala 64:22]
  wire  routers_auto_ingress_nodes_in_flit_bits_head; // @[NoC.scala 64:22]
  wire  routers_auto_ingress_nodes_in_flit_bits_tail; // @[NoC.scala 64:22]
  wire [63:0] routers_auto_ingress_nodes_in_flit_bits_payload; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_ingress_nodes_in_flit_bits_egress_id; // @[NoC.scala 64:22]
  wire  routers_auto_source_nodes_out_1_flit_0_valid; // @[NoC.scala 64:22]
  wire  routers_auto_source_nodes_out_1_flit_0_bits_head; // @[NoC.scala 64:22]
  wire  routers_auto_source_nodes_out_1_flit_0_bits_tail; // @[NoC.scala 64:22]
  wire [63:0] routers_auto_source_nodes_out_1_flit_0_bits_payload; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_source_nodes_out_1_flit_0_bits_flow_ingress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_source_nodes_out_1_flit_0_bits_flow_egress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_source_nodes_out_1_flit_0_bits_virt_channel_id; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_source_nodes_out_1_credit_return; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_source_nodes_out_1_vc_free; // @[NoC.scala 64:22]
  wire  routers_auto_source_nodes_out_0_flit_0_valid; // @[NoC.scala 64:22]
  wire  routers_auto_source_nodes_out_0_flit_0_bits_head; // @[NoC.scala 64:22]
  wire  routers_auto_source_nodes_out_0_flit_0_bits_tail; // @[NoC.scala 64:22]
  wire [63:0] routers_auto_source_nodes_out_0_flit_0_bits_payload; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_source_nodes_out_0_flit_0_bits_flow_ingress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_source_nodes_out_0_flit_0_bits_flow_egress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_source_nodes_out_0_flit_0_bits_virt_channel_id; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_source_nodes_out_0_credit_return; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_source_nodes_out_0_vc_free; // @[NoC.scala 64:22]
  wire  routers_auto_dest_nodes_in_1_flit_0_valid; // @[NoC.scala 64:22]
  wire  routers_auto_dest_nodes_in_1_flit_0_bits_head; // @[NoC.scala 64:22]
  wire  routers_auto_dest_nodes_in_1_flit_0_bits_tail; // @[NoC.scala 64:22]
  wire [63:0] routers_auto_dest_nodes_in_1_flit_0_bits_payload; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_dest_nodes_in_1_flit_0_bits_flow_ingress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_dest_nodes_in_1_flit_0_bits_flow_egress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_dest_nodes_in_1_flit_0_bits_virt_channel_id; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_dest_nodes_in_1_credit_return; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_dest_nodes_in_1_vc_free; // @[NoC.scala 64:22]
  wire  routers_auto_dest_nodes_in_0_flit_0_valid; // @[NoC.scala 64:22]
  wire  routers_auto_dest_nodes_in_0_flit_0_bits_head; // @[NoC.scala 64:22]
  wire  routers_auto_dest_nodes_in_0_flit_0_bits_tail; // @[NoC.scala 64:22]
  wire [63:0] routers_auto_dest_nodes_in_0_flit_0_bits_payload; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_dest_nodes_in_0_flit_0_bits_flow_ingress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_dest_nodes_in_0_flit_0_bits_flow_egress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_dest_nodes_in_0_flit_0_bits_virt_channel_id; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_dest_nodes_in_0_credit_return; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_dest_nodes_in_0_vc_free; // @[NoC.scala 64:22]
  Router routers ( // @[NoC.scala 64:22]
    .clock(routers_clock),
    .reset(routers_reset),
    .auto_debug_out_va_stall_0(routers_auto_debug_out_va_stall_0),
    .auto_debug_out_va_stall_1(routers_auto_debug_out_va_stall_1),
    .auto_debug_out_sa_stall_0(routers_auto_debug_out_sa_stall_0),
    .auto_debug_out_sa_stall_1(routers_auto_debug_out_sa_stall_1),
    .auto_egress_nodes_out_flit_valid(routers_auto_egress_nodes_out_flit_valid),
    .auto_egress_nodes_out_flit_bits_head(routers_auto_egress_nodes_out_flit_bits_head),
    .auto_egress_nodes_out_flit_bits_tail(routers_auto_egress_nodes_out_flit_bits_tail),
    .auto_egress_nodes_out_flit_bits_payload(routers_auto_egress_nodes_out_flit_bits_payload),
    .auto_egress_nodes_out_flit_bits_ingress_id(routers_auto_egress_nodes_out_flit_bits_ingress_id),
    .auto_ingress_nodes_in_flit_ready(routers_auto_ingress_nodes_in_flit_ready),
    .auto_ingress_nodes_in_flit_valid(routers_auto_ingress_nodes_in_flit_valid),
    .auto_ingress_nodes_in_flit_bits_head(routers_auto_ingress_nodes_in_flit_bits_head),
    .auto_ingress_nodes_in_flit_bits_tail(routers_auto_ingress_nodes_in_flit_bits_tail),
    .auto_ingress_nodes_in_flit_bits_payload(routers_auto_ingress_nodes_in_flit_bits_payload),
    .auto_ingress_nodes_in_flit_bits_egress_id(routers_auto_ingress_nodes_in_flit_bits_egress_id),
    .auto_source_nodes_out_1_flit_0_valid(routers_auto_source_nodes_out_1_flit_0_valid),
    .auto_source_nodes_out_1_flit_0_bits_head(routers_auto_source_nodes_out_1_flit_0_bits_head),
    .auto_source_nodes_out_1_flit_0_bits_tail(routers_auto_source_nodes_out_1_flit_0_bits_tail),
    .auto_source_nodes_out_1_flit_0_bits_payload(routers_auto_source_nodes_out_1_flit_0_bits_payload),
    .auto_source_nodes_out_1_flit_0_bits_flow_ingress_node(routers_auto_source_nodes_out_1_flit_0_bits_flow_ingress_node
      ),
    .auto_source_nodes_out_1_flit_0_bits_flow_egress_node(routers_auto_source_nodes_out_1_flit_0_bits_flow_egress_node),
    .auto_source_nodes_out_1_flit_0_bits_virt_channel_id(routers_auto_source_nodes_out_1_flit_0_bits_virt_channel_id),
    .auto_source_nodes_out_1_credit_return(routers_auto_source_nodes_out_1_credit_return),
    .auto_source_nodes_out_1_vc_free(routers_auto_source_nodes_out_1_vc_free),
    .auto_source_nodes_out_0_flit_0_valid(routers_auto_source_nodes_out_0_flit_0_valid),
    .auto_source_nodes_out_0_flit_0_bits_head(routers_auto_source_nodes_out_0_flit_0_bits_head),
    .auto_source_nodes_out_0_flit_0_bits_tail(routers_auto_source_nodes_out_0_flit_0_bits_tail),
    .auto_source_nodes_out_0_flit_0_bits_payload(routers_auto_source_nodes_out_0_flit_0_bits_payload),
    .auto_source_nodes_out_0_flit_0_bits_flow_ingress_node(routers_auto_source_nodes_out_0_flit_0_bits_flow_ingress_node
      ),
    .auto_source_nodes_out_0_flit_0_bits_flow_egress_node(routers_auto_source_nodes_out_0_flit_0_bits_flow_egress_node),
    .auto_source_nodes_out_0_flit_0_bits_virt_channel_id(routers_auto_source_nodes_out_0_flit_0_bits_virt_channel_id),
    .auto_source_nodes_out_0_credit_return(routers_auto_source_nodes_out_0_credit_return),
    .auto_source_nodes_out_0_vc_free(routers_auto_source_nodes_out_0_vc_free),
    .auto_dest_nodes_in_1_flit_0_valid(routers_auto_dest_nodes_in_1_flit_0_valid),
    .auto_dest_nodes_in_1_flit_0_bits_head(routers_auto_dest_nodes_in_1_flit_0_bits_head),
    .auto_dest_nodes_in_1_flit_0_bits_tail(routers_auto_dest_nodes_in_1_flit_0_bits_tail),
    .auto_dest_nodes_in_1_flit_0_bits_payload(routers_auto_dest_nodes_in_1_flit_0_bits_payload),
    .auto_dest_nodes_in_1_flit_0_bits_flow_ingress_node(routers_auto_dest_nodes_in_1_flit_0_bits_flow_ingress_node),
    .auto_dest_nodes_in_1_flit_0_bits_flow_egress_node(routers_auto_dest_nodes_in_1_flit_0_bits_flow_egress_node),
    .auto_dest_nodes_in_1_flit_0_bits_virt_channel_id(routers_auto_dest_nodes_in_1_flit_0_bits_virt_channel_id),
    .auto_dest_nodes_in_1_credit_return(routers_auto_dest_nodes_in_1_credit_return),
    .auto_dest_nodes_in_1_vc_free(routers_auto_dest_nodes_in_1_vc_free),
    .auto_dest_nodes_in_0_flit_0_valid(routers_auto_dest_nodes_in_0_flit_0_valid),
    .auto_dest_nodes_in_0_flit_0_bits_head(routers_auto_dest_nodes_in_0_flit_0_bits_head),
    .auto_dest_nodes_in_0_flit_0_bits_tail(routers_auto_dest_nodes_in_0_flit_0_bits_tail),
    .auto_dest_nodes_in_0_flit_0_bits_payload(routers_auto_dest_nodes_in_0_flit_0_bits_payload),
    .auto_dest_nodes_in_0_flit_0_bits_flow_ingress_node(routers_auto_dest_nodes_in_0_flit_0_bits_flow_ingress_node),
    .auto_dest_nodes_in_0_flit_0_bits_flow_egress_node(routers_auto_dest_nodes_in_0_flit_0_bits_flow_egress_node),
    .auto_dest_nodes_in_0_flit_0_bits_virt_channel_id(routers_auto_dest_nodes_in_0_flit_0_bits_virt_channel_id),
    .auto_dest_nodes_in_0_credit_return(routers_auto_dest_nodes_in_0_credit_return),
    .auto_dest_nodes_in_0_vc_free(routers_auto_dest_nodes_in_0_vc_free)
  );
  assign auto_routers_debug_out_va_stall_0 = routers_auto_debug_out_va_stall_0; // @[LazyModule.scala 368:12]
  assign auto_routers_debug_out_va_stall_1 = routers_auto_debug_out_va_stall_1; // @[LazyModule.scala 368:12]
  assign auto_routers_debug_out_sa_stall_0 = routers_auto_debug_out_sa_stall_0; // @[LazyModule.scala 368:12]
  assign auto_routers_debug_out_sa_stall_1 = routers_auto_debug_out_sa_stall_1; // @[LazyModule.scala 368:12]
  assign auto_routers_egress_nodes_out_flit_valid = routers_auto_egress_nodes_out_flit_valid; // @[LazyModule.scala 368:12]
  assign auto_routers_egress_nodes_out_flit_bits_head = routers_auto_egress_nodes_out_flit_bits_head; // @[LazyModule.scala 368:12]
  assign auto_routers_egress_nodes_out_flit_bits_tail = routers_auto_egress_nodes_out_flit_bits_tail; // @[LazyModule.scala 368:12]
  assign auto_routers_egress_nodes_out_flit_bits_payload = routers_auto_egress_nodes_out_flit_bits_payload; // @[LazyModule.scala 368:12]
  assign auto_routers_egress_nodes_out_flit_bits_ingress_id = routers_auto_egress_nodes_out_flit_bits_ingress_id; // @[LazyModule.scala 368:12]
  assign auto_routers_ingress_nodes_in_flit_ready = routers_auto_ingress_nodes_in_flit_ready; // @[LazyModule.scala 366:16]
  assign auto_routers_source_nodes_out_1_flit_0_valid = routers_auto_source_nodes_out_1_flit_0_valid; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_1_flit_0_bits_head = routers_auto_source_nodes_out_1_flit_0_bits_head; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_1_flit_0_bits_tail = routers_auto_source_nodes_out_1_flit_0_bits_tail; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_1_flit_0_bits_payload = routers_auto_source_nodes_out_1_flit_0_bits_payload; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_1_flit_0_bits_flow_ingress_node =
    routers_auto_source_nodes_out_1_flit_0_bits_flow_ingress_node; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_1_flit_0_bits_flow_egress_node =
    routers_auto_source_nodes_out_1_flit_0_bits_flow_egress_node; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_1_flit_0_bits_virt_channel_id =
    routers_auto_source_nodes_out_1_flit_0_bits_virt_channel_id; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_0_flit_0_valid = routers_auto_source_nodes_out_0_flit_0_valid; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_0_flit_0_bits_head = routers_auto_source_nodes_out_0_flit_0_bits_head; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_0_flit_0_bits_tail = routers_auto_source_nodes_out_0_flit_0_bits_tail; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_0_flit_0_bits_payload = routers_auto_source_nodes_out_0_flit_0_bits_payload; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_0_flit_0_bits_flow_ingress_node =
    routers_auto_source_nodes_out_0_flit_0_bits_flow_ingress_node; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_0_flit_0_bits_flow_egress_node =
    routers_auto_source_nodes_out_0_flit_0_bits_flow_egress_node; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_0_flit_0_bits_virt_channel_id =
    routers_auto_source_nodes_out_0_flit_0_bits_virt_channel_id; // @[LazyModule.scala 368:12]
  assign auto_routers_dest_nodes_in_1_credit_return = routers_auto_dest_nodes_in_1_credit_return; // @[LazyModule.scala 366:16]
  assign auto_routers_dest_nodes_in_1_vc_free = routers_auto_dest_nodes_in_1_vc_free; // @[LazyModule.scala 366:16]
  assign auto_routers_dest_nodes_in_0_credit_return = routers_auto_dest_nodes_in_0_credit_return; // @[LazyModule.scala 366:16]
  assign auto_routers_dest_nodes_in_0_vc_free = routers_auto_dest_nodes_in_0_vc_free; // @[LazyModule.scala 366:16]
  assign routers_clock = auto_clock_in_clock; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign routers_reset = auto_clock_in_reset; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign routers_auto_ingress_nodes_in_flit_valid = auto_routers_ingress_nodes_in_flit_valid; // @[LazyModule.scala 366:16]
  assign routers_auto_ingress_nodes_in_flit_bits_head = auto_routers_ingress_nodes_in_flit_bits_head; // @[LazyModule.scala 366:16]
  assign routers_auto_ingress_nodes_in_flit_bits_tail = auto_routers_ingress_nodes_in_flit_bits_tail; // @[LazyModule.scala 366:16]
  assign routers_auto_ingress_nodes_in_flit_bits_payload = auto_routers_ingress_nodes_in_flit_bits_payload; // @[LazyModule.scala 366:16]
  assign routers_auto_ingress_nodes_in_flit_bits_egress_id = auto_routers_ingress_nodes_in_flit_bits_egress_id; // @[LazyModule.scala 366:16]
  assign routers_auto_source_nodes_out_1_credit_return = auto_routers_source_nodes_out_1_credit_return; // @[LazyModule.scala 368:12]
  assign routers_auto_source_nodes_out_1_vc_free = auto_routers_source_nodes_out_1_vc_free; // @[LazyModule.scala 368:12]
  assign routers_auto_source_nodes_out_0_credit_return = auto_routers_source_nodes_out_0_credit_return; // @[LazyModule.scala 368:12]
  assign routers_auto_source_nodes_out_0_vc_free = auto_routers_source_nodes_out_0_vc_free; // @[LazyModule.scala 368:12]
  assign routers_auto_dest_nodes_in_1_flit_0_valid = auto_routers_dest_nodes_in_1_flit_0_valid; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_1_flit_0_bits_head = auto_routers_dest_nodes_in_1_flit_0_bits_head; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_1_flit_0_bits_tail = auto_routers_dest_nodes_in_1_flit_0_bits_tail; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_1_flit_0_bits_payload = auto_routers_dest_nodes_in_1_flit_0_bits_payload; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_1_flit_0_bits_flow_ingress_node =
    auto_routers_dest_nodes_in_1_flit_0_bits_flow_ingress_node; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_1_flit_0_bits_flow_egress_node =
    auto_routers_dest_nodes_in_1_flit_0_bits_flow_egress_node; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_1_flit_0_bits_virt_channel_id =
    auto_routers_dest_nodes_in_1_flit_0_bits_virt_channel_id; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_0_flit_0_valid = auto_routers_dest_nodes_in_0_flit_0_valid; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_0_flit_0_bits_head = auto_routers_dest_nodes_in_0_flit_0_bits_head; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_0_flit_0_bits_tail = auto_routers_dest_nodes_in_0_flit_0_bits_tail; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_0_flit_0_bits_payload = auto_routers_dest_nodes_in_0_flit_0_bits_payload; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_0_flit_0_bits_flow_ingress_node =
    auto_routers_dest_nodes_in_0_flit_0_bits_flow_ingress_node; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_0_flit_0_bits_flow_egress_node =
    auto_routers_dest_nodes_in_0_flit_0_bits_flow_egress_node; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_0_flit_0_bits_virt_channel_id =
    auto_routers_dest_nodes_in_0_flit_0_bits_virt_channel_id; // @[LazyModule.scala 366:16]
endmodule
module NoCMonitor_2(
  input        clock,
  input        reset,
  input        io_in_flit_0_valid,
  input        io_in_flit_0_bits_head,
  input        io_in_flit_0_bits_tail,
  input  [1:0] io_in_flit_0_bits_flow_ingress_node,
  input  [1:0] io_in_flit_0_bits_flow_egress_node,
  input  [1:0] io_in_flit_0_bits_virt_channel_id
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg  in_flight_0; // @[Monitor.scala 16:26]
  reg  in_flight_1; // @[Monitor.scala 16:26]
  reg  in_flight_2; // @[Monitor.scala 16:26]
  reg  in_flight_3; // @[Monitor.scala 16:26]
  wire  _GEN_0 = 2'h0 == io_in_flit_0_bits_virt_channel_id | in_flight_0; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_1 = 2'h1 == io_in_flit_0_bits_virt_channel_id | in_flight_1; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_2 = 2'h2 == io_in_flit_0_bits_virt_channel_id | in_flight_2; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_3 = 2'h3 == io_in_flit_0_bits_virt_channel_id | in_flight_3; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_5 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? in_flight_1 : in_flight_0; // @[Monitor.scala 22:{17,17}]
  wire  _GEN_6 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? in_flight_2 : _GEN_5; // @[Monitor.scala 22:{17,17}]
  wire  _GEN_7 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? in_flight_3 : _GEN_6; // @[Monitor.scala 22:{17,17}]
  wire  _T_2 = ~reset; // @[Monitor.scala 22:16]
  wire  _GEN_8 = io_in_flit_0_bits_head ? _GEN_0 : in_flight_0; // @[Monitor.scala 16:26 20:29]
  wire  _GEN_9 = io_in_flit_0_bits_head ? _GEN_1 : in_flight_1; // @[Monitor.scala 16:26 20:29]
  wire  _GEN_10 = io_in_flit_0_bits_head ? _GEN_2 : in_flight_2; // @[Monitor.scala 16:26 20:29]
  wire  _GEN_11 = io_in_flit_0_bits_head ? _GEN_3 : in_flight_3; // @[Monitor.scala 16:26 20:29]
  wire  _T_4 = io_in_flit_0_valid & io_in_flit_0_bits_head; // @[Monitor.scala 29:22]
  wire  _T_7 = io_in_flit_0_bits_flow_egress_node == 2'h1; // @[Types.scala 54:21]
  wire  _T_8 = io_in_flit_0_bits_flow_ingress_node == 2'h3 & _T_7; // @[Types.scala 53:39]
  wire  _T_20 = io_in_flit_0_bits_flow_ingress_node == 2'h0 & _T_7; // @[Types.scala 53:39]
  wire  _T_26 = io_in_flit_0_bits_flow_egress_node == 2'h2; // @[Types.scala 54:21]
  wire  _T_27 = io_in_flit_0_bits_flow_ingress_node == 2'h0 & _T_26; // @[Types.scala 53:39]
  wire  _T_40 = _T_20 | _T_27 | _T_8; // @[package.scala 73:59]
  wire  _GEN_29 = _T_4 & ~reset; // @[Monitor.scala 22:16]
  always @(posedge clock) begin
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_0 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h0 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_0 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_0 <= _GEN_8;
        end
      end else begin
        in_flight_0 <= _GEN_8;
      end
    end
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_1 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h1 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_1 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_1 <= _GEN_9;
        end
      end else begin
        in_flight_1 <= _GEN_9;
      end
    end
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_2 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h2 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_2 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_2 <= _GEN_10;
        end
      end else begin
        in_flight_2 <= _GEN_10;
      end
    end
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_3 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h3 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_3 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_3 <= _GEN_11;
        end
      end else begin
        in_flight_3 <= _GEN_11;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4 & ~reset & ~(~_GEN_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed: Flit head/tail sequencing is broken\n    at Monitor.scala:22 assert (!in_flight(flit.bits.virt_channel_id), \"Flit head/tail sequencing is broken\")\n"
            ); // @[Monitor.scala 22:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h0 | _T_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h1 | _T_40)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h2 | _T_40)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h3 | _T_40)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  in_flight_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  in_flight_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  in_flight_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  in_flight_3 = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (_T_4 & ~reset) begin
      assert(~_GEN_7); // @[Monitor.scala 22:16]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h0 | _T_8); // @[Monitor.scala 32:17]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h1 | _T_40); // @[Monitor.scala 32:17]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h2 | _T_40); // @[Monitor.scala 32:17]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h3 | _T_40); // @[Monitor.scala 32:17]
    end
  end
endmodule
module NoCMonitor_3(
  input        clock,
  input        reset,
  input        io_in_flit_0_valid,
  input        io_in_flit_0_bits_head,
  input        io_in_flit_0_bits_tail,
  input  [1:0] io_in_flit_0_bits_flow_ingress_node,
  input  [1:0] io_in_flit_0_bits_flow_egress_node,
  input  [1:0] io_in_flit_0_bits_virt_channel_id
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg  in_flight_0; // @[Monitor.scala 16:26]
  reg  in_flight_1; // @[Monitor.scala 16:26]
  reg  in_flight_2; // @[Monitor.scala 16:26]
  reg  in_flight_3; // @[Monitor.scala 16:26]
  wire  _GEN_0 = 2'h0 == io_in_flit_0_bits_virt_channel_id | in_flight_0; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_1 = 2'h1 == io_in_flit_0_bits_virt_channel_id | in_flight_1; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_2 = 2'h2 == io_in_flit_0_bits_virt_channel_id | in_flight_2; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_3 = 2'h3 == io_in_flit_0_bits_virt_channel_id | in_flight_3; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_5 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? in_flight_1 : in_flight_0; // @[Monitor.scala 22:{17,17}]
  wire  _GEN_6 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? in_flight_2 : _GEN_5; // @[Monitor.scala 22:{17,17}]
  wire  _GEN_7 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? in_flight_3 : _GEN_6; // @[Monitor.scala 22:{17,17}]
  wire  _T_2 = ~reset; // @[Monitor.scala 22:16]
  wire  _GEN_8 = io_in_flit_0_bits_head ? _GEN_0 : in_flight_0; // @[Monitor.scala 16:26 20:29]
  wire  _GEN_9 = io_in_flit_0_bits_head ? _GEN_1 : in_flight_1; // @[Monitor.scala 16:26 20:29]
  wire  _GEN_10 = io_in_flit_0_bits_head ? _GEN_2 : in_flight_2; // @[Monitor.scala 16:26 20:29]
  wire  _GEN_11 = io_in_flit_0_bits_head ? _GEN_3 : in_flight_3; // @[Monitor.scala 16:26 20:29]
  wire  _T_4 = io_in_flit_0_valid & io_in_flit_0_bits_head; // @[Monitor.scala 29:22]
  wire  _T_7 = io_in_flit_0_bits_flow_egress_node == 2'h1; // @[Types.scala 54:21]
  wire  _T_8 = io_in_flit_0_bits_flow_ingress_node == 2'h3 & _T_7; // @[Types.scala 53:39]
  wire  _T_19 = io_in_flit_0_bits_flow_egress_node == 2'h0; // @[Types.scala 54:21]
  wire  _T_20 = io_in_flit_0_bits_flow_ingress_node == 2'h2 & _T_19; // @[Types.scala 53:39]
  wire  _T_27 = io_in_flit_0_bits_flow_ingress_node == 2'h2 & _T_7; // @[Types.scala 53:39]
  wire  _T_40 = _T_20 | _T_27 | _T_8; // @[package.scala 73:59]
  wire  _GEN_29 = _T_4 & ~reset; // @[Monitor.scala 22:16]
  always @(posedge clock) begin
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_0 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h0 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_0 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_0 <= _GEN_8;
        end
      end else begin
        in_flight_0 <= _GEN_8;
      end
    end
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_1 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h1 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_1 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_1 <= _GEN_9;
        end
      end else begin
        in_flight_1 <= _GEN_9;
      end
    end
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_2 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h2 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_2 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_2 <= _GEN_10;
        end
      end else begin
        in_flight_2 <= _GEN_10;
      end
    end
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_3 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h3 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_3 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_3 <= _GEN_11;
        end
      end else begin
        in_flight_3 <= _GEN_11;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4 & ~reset & ~(~_GEN_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed: Flit head/tail sequencing is broken\n    at Monitor.scala:22 assert (!in_flight(flit.bits.virt_channel_id), \"Flit head/tail sequencing is broken\")\n"
            ); // @[Monitor.scala 22:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h0 | _T_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h1 | _T_40)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h2 | _T_40)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h3 | _T_40)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  in_flight_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  in_flight_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  in_flight_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  in_flight_3 = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (_T_4 & ~reset) begin
      assert(~_GEN_7); // @[Monitor.scala 22:16]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h0 | _T_8); // @[Monitor.scala 32:17]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h1 | _T_40); // @[Monitor.scala 32:17]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h2 | _T_40); // @[Monitor.scala 32:17]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h3 | _T_40); // @[Monitor.scala 32:17]
    end
  end
endmodule
module InputUnit_2(
  input         clock,
  input         reset,
  output        io_router_req_valid,
  output [1:0]  io_router_req_bits_src_virt_id,
  output [1:0]  io_router_req_bits_flow_ingress_node,
  output [1:0]  io_router_req_bits_flow_egress_node,
  input         io_router_resp_vc_sel_1_0,
  input         io_router_resp_vc_sel_1_1,
  input         io_router_resp_vc_sel_1_2,
  input         io_router_resp_vc_sel_1_3,
  input         io_router_resp_vc_sel_0_0,
  input         io_router_resp_vc_sel_0_1,
  input         io_router_resp_vc_sel_0_2,
  input         io_router_resp_vc_sel_0_3,
  input         io_vcalloc_req_ready,
  output        io_vcalloc_req_valid,
  output        io_vcalloc_req_bits_vc_sel_2_0,
  output        io_vcalloc_req_bits_vc_sel_1_0,
  output        io_vcalloc_req_bits_vc_sel_1_1,
  output        io_vcalloc_req_bits_vc_sel_1_2,
  output        io_vcalloc_req_bits_vc_sel_1_3,
  output        io_vcalloc_req_bits_vc_sel_0_0,
  output        io_vcalloc_req_bits_vc_sel_0_1,
  output        io_vcalloc_req_bits_vc_sel_0_2,
  output        io_vcalloc_req_bits_vc_sel_0_3,
  input         io_vcalloc_resp_vc_sel_2_0,
  input         io_vcalloc_resp_vc_sel_1_0,
  input         io_vcalloc_resp_vc_sel_1_1,
  input         io_vcalloc_resp_vc_sel_1_2,
  input         io_vcalloc_resp_vc_sel_1_3,
  input         io_vcalloc_resp_vc_sel_0_0,
  input         io_vcalloc_resp_vc_sel_0_1,
  input         io_vcalloc_resp_vc_sel_0_2,
  input         io_vcalloc_resp_vc_sel_0_3,
  input         io_out_credit_available_2_0,
  input         io_out_credit_available_1_0,
  input         io_out_credit_available_1_1,
  input         io_out_credit_available_1_2,
  input         io_out_credit_available_1_3,
  input         io_out_credit_available_0_0,
  input         io_out_credit_available_0_1,
  input         io_out_credit_available_0_2,
  input         io_out_credit_available_0_3,
  input         io_salloc_req_0_ready,
  output        io_salloc_req_0_valid,
  output        io_salloc_req_0_bits_vc_sel_2_0,
  output        io_salloc_req_0_bits_vc_sel_1_0,
  output        io_salloc_req_0_bits_vc_sel_1_1,
  output        io_salloc_req_0_bits_vc_sel_1_2,
  output        io_salloc_req_0_bits_vc_sel_1_3,
  output        io_salloc_req_0_bits_vc_sel_0_0,
  output        io_salloc_req_0_bits_vc_sel_0_1,
  output        io_salloc_req_0_bits_vc_sel_0_2,
  output        io_salloc_req_0_bits_vc_sel_0_3,
  output        io_salloc_req_0_bits_tail,
  output        io_out_0_valid,
  output        io_out_0_bits_flit_head,
  output        io_out_0_bits_flit_tail,
  output [63:0] io_out_0_bits_flit_payload,
  output [1:0]  io_out_0_bits_flit_flow_ingress_node,
  output [1:0]  io_out_0_bits_flit_flow_egress_node,
  output [1:0]  io_out_0_bits_out_virt_channel,
  output [1:0]  io_debug_va_stall,
  output [1:0]  io_debug_sa_stall,
  input         io_in_flit_0_valid,
  input         io_in_flit_0_bits_head,
  input         io_in_flit_0_bits_tail,
  input  [63:0] io_in_flit_0_bits_payload,
  input  [1:0]  io_in_flit_0_bits_flow_ingress_node,
  input  [1:0]  io_in_flit_0_bits_flow_egress_node,
  input  [1:0]  io_in_flit_0_bits_virt_channel_id,
  output [3:0]  io_in_credit_return,
  output [3:0]  io_in_vc_free
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
`endif // RANDOMIZE_REG_INIT
  wire  input_buffer_clock; // @[InputUnit.scala 180:28]
  wire  input_buffer_reset; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_enq_0_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_enq_0_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_enq_0_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_enq_0_bits_payload; // @[InputUnit.scala 180:28]
  wire [1:0] input_buffer_io_enq_0_bits_virt_channel_id; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_0_ready; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_0_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_0_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_0_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_deq_0_bits_payload; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_ready; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_deq_1_bits_payload; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_ready; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_deq_2_bits_payload; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_3_ready; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_3_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_3_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_3_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_deq_3_bits_payload; // @[InputUnit.scala 180:28]
  wire  route_arbiter_io_in_0_valid; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_0_bits_flow_ingress_node; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_0_bits_flow_egress_node; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_1_ready; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_1_valid; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_1_bits_flow_ingress_node; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_1_bits_flow_egress_node; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_2_ready; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_2_valid; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_2_bits_flow_ingress_node; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_2_bits_flow_egress_node; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_3_ready; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_3_valid; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_3_bits_flow_ingress_node; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_3_bits_flow_egress_node; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_out_valid; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_out_bits_src_virt_id; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_out_bits_flow_ingress_node; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_out_bits_flow_egress_node; // @[InputUnit.scala 186:29]
  wire  salloc_arb_clock; // @[InputUnit.scala 279:26]
  wire  salloc_arb_reset; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_bits_vc_sel_2_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_bits_vc_sel_1_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_bits_tail; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_vc_sel_2_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_vc_sel_1_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_vc_sel_1_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_vc_sel_0_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_tail; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_2_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_1_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_1_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_1_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_0_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_0_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_tail; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_2_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_1_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_1_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_1_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_1_3; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_0_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_0_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_0_3; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_tail; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_2_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_1_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_1_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_1_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_1_3; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_0_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_0_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_0_3; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_tail; // @[InputUnit.scala 279:26]
  wire [3:0] salloc_arb_io_chosen_oh_0; // @[InputUnit.scala 279:26]
  reg [2:0] states_0_g; // @[InputUnit.scala 191:19]
  reg  states_0_vc_sel_2_0; // @[InputUnit.scala 191:19]
  reg  states_0_vc_sel_1_0; // @[InputUnit.scala 191:19]
  reg  states_0_vc_sel_0_0; // @[InputUnit.scala 191:19]
  reg [1:0] states_0_flow_ingress_node; // @[InputUnit.scala 191:19]
  reg [1:0] states_0_flow_egress_node; // @[InputUnit.scala 191:19]
  reg [2:0] states_1_g; // @[InputUnit.scala 191:19]
  reg  states_1_vc_sel_2_0; // @[InputUnit.scala 191:19]
  reg  states_1_vc_sel_1_0; // @[InputUnit.scala 191:19]
  reg  states_1_vc_sel_1_1; // @[InputUnit.scala 191:19]
  reg  states_1_vc_sel_0_1; // @[InputUnit.scala 191:19]
  reg [1:0] states_1_flow_ingress_node; // @[InputUnit.scala 191:19]
  reg [1:0] states_1_flow_egress_node; // @[InputUnit.scala 191:19]
  reg [2:0] states_2_g; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_2_0; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_1_0; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_1_1; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_1_2; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_0_1; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_0_2; // @[InputUnit.scala 191:19]
  reg [1:0] states_2_flow_ingress_node; // @[InputUnit.scala 191:19]
  reg [1:0] states_2_flow_egress_node; // @[InputUnit.scala 191:19]
  reg [2:0] states_3_g; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_2_0; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_1_0; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_1_1; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_1_2; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_1_3; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_0_1; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_0_2; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_0_3; // @[InputUnit.scala 191:19]
  reg [1:0] states_3_flow_ingress_node; // @[InputUnit.scala 191:19]
  reg [1:0] states_3_flow_egress_node; // @[InputUnit.scala 191:19]
  wire  _T = io_in_flit_0_valid & io_in_flit_0_bits_head; // @[InputUnit.scala 194:32]
  wire  _T_3 = ~reset; // @[InputUnit.scala 196:13]
  wire [2:0] _GEN_1 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? states_1_g : states_0_g; // @[InputUnit.scala 197:{27,27}]
  wire [2:0] _GEN_2 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? states_2_g : _GEN_1; // @[InputUnit.scala 197:{27,27}]
  wire [2:0] _GEN_3 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? states_3_g : _GEN_2; // @[InputUnit.scala 197:{27,27}]
  wire  at_dest = io_in_flit_0_bits_flow_egress_node == 2'h1; // @[InputUnit.scala 198:57]
  wire [2:0] _states_g_T = at_dest ? 3'h2 : 3'h1; // @[InputUnit.scala 199:26]
  wire [2:0] _GEN_4 = 2'h0 == io_in_flit_0_bits_virt_channel_id ? _states_g_T : states_0_g; // @[InputUnit.scala 191:19 199:{20,20}]
  wire [2:0] _GEN_5 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? _states_g_T : states_1_g; // @[InputUnit.scala 191:19 199:{20,20}]
  wire [2:0] _GEN_6 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? _states_g_T : states_2_g; // @[InputUnit.scala 191:19 199:{20,20}]
  wire [2:0] _GEN_7 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? _states_g_T : states_3_g; // @[InputUnit.scala 191:19 199:{20,20}]
  wire  _GEN_8 = 2'h0 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_0_vc_sel_0_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_13 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_1_vc_sel_0_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_14 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_0_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_15 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_0_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_18 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_0_2; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_19 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_0_2; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_23 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_0_3; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_24 = 2'h0 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_0_vc_sel_1_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_25 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_1_vc_sel_1_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_26 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_1_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_27 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_1_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_29 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_1_vc_sel_1_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_30 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_1_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_31 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_1_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_34 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_1_2; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_35 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_1_2; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_39 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_1_3; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_40 = 2'h0 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_0_vc_sel_2_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_41 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_1_vc_sel_2_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_42 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_2_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_43 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_2_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_44 = 2'h0 == io_in_flit_0_bits_virt_channel_id | _GEN_40; // @[InputUnit.scala 203:{44,44}]
  wire  _GEN_45 = 2'h1 == io_in_flit_0_bits_virt_channel_id | _GEN_41; // @[InputUnit.scala 203:{44,44}]
  wire  _GEN_46 = 2'h2 == io_in_flit_0_bits_virt_channel_id | _GEN_42; // @[InputUnit.scala 203:{44,44}]
  wire  _GEN_47 = 2'h3 == io_in_flit_0_bits_virt_channel_id | _GEN_43; // @[InputUnit.scala 203:{44,44}]
  wire [2:0] _GEN_72 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_4 : states_0_g; // @[InputUnit.scala 191:19 194:60]
  wire [2:0] _GEN_73 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_5 : states_1_g; // @[InputUnit.scala 191:19 194:60]
  wire [2:0] _GEN_74 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_6 : states_2_g; // @[InputUnit.scala 191:19 194:60]
  wire [2:0] _GEN_75 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_7 : states_3_g; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_76 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_8 : states_0_vc_sel_0_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_81 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_13 : states_1_vc_sel_0_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_82 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_14 : states_2_vc_sel_0_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_83 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_15 : states_3_vc_sel_0_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_86 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_18 : states_2_vc_sel_0_2; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_87 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_19 : states_3_vc_sel_0_2; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_91 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_23 : states_3_vc_sel_0_3; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_92 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_24 : states_0_vc_sel_1_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_93 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_25 : states_1_vc_sel_1_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_94 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_26 : states_2_vc_sel_1_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_95 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_27 : states_3_vc_sel_1_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_97 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_29 : states_1_vc_sel_1_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_98 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_30 : states_2_vc_sel_1_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_99 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_31 : states_3_vc_sel_1_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_102 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_34 : states_2_vc_sel_1_2; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_103 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_35 : states_3_vc_sel_1_2; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_107 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_39 : states_3_vc_sel_1_3; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_108 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_44 : states_0_vc_sel_2_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_109 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_45 : states_1_vc_sel_2_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_110 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_46 : states_2_vc_sel_2_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_111 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_47 : states_3_vc_sel_2_0; // @[InputUnit.scala 191:19 194:60]
  wire  _T_10 = route_arbiter_io_in_0_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_132 = _T_10 ? 3'h2 : _GEN_72; // @[InputUnit.scala 215:{23,29}]
  wire  _T_11 = route_arbiter_io_in_1_ready & route_arbiter_io_in_1_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_133 = _T_11 ? 3'h2 : _GEN_73; // @[InputUnit.scala 215:{23,29}]
  wire  _T_12 = route_arbiter_io_in_2_ready & route_arbiter_io_in_2_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_134 = _T_12 ? 3'h2 : _GEN_74; // @[InputUnit.scala 215:{23,29}]
  wire  _T_13 = route_arbiter_io_in_3_ready & route_arbiter_io_in_3_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_135 = _T_13 ? 3'h2 : _GEN_75; // @[InputUnit.scala 215:{23,29}]
  wire [2:0] _GEN_137 = 2'h1 == io_router_req_bits_src_virt_id ? states_1_g : states_0_g; // @[InputUnit.scala 224:{25,25}]
  wire [2:0] _GEN_138 = 2'h2 == io_router_req_bits_src_virt_id ? states_2_g : _GEN_137; // @[InputUnit.scala 224:{25,25}]
  wire [2:0] _GEN_139 = 2'h3 == io_router_req_bits_src_virt_id ? states_3_g : _GEN_138; // @[InputUnit.scala 224:{25,25}]
  wire [2:0] _GEN_140 = 2'h0 == io_router_req_bits_src_virt_id ? 3'h2 : _GEN_132; // @[InputUnit.scala 225:{18,18}]
  wire [2:0] _GEN_141 = 2'h1 == io_router_req_bits_src_virt_id ? 3'h2 : _GEN_133; // @[InputUnit.scala 225:{18,18}]
  wire [2:0] _GEN_142 = 2'h2 == io_router_req_bits_src_virt_id ? 3'h2 : _GEN_134; // @[InputUnit.scala 225:{18,18}]
  wire [2:0] _GEN_143 = 2'h3 == io_router_req_bits_src_virt_id ? 3'h2 : _GEN_135; // @[InputUnit.scala 225:{18,18}]
  wire  _GEN_144 = 2'h0 == io_router_req_bits_src_virt_id ? 1'h0 : _GEN_108; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_145 = 2'h0 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_0 : _GEN_92; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_149 = 2'h0 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_0 : _GEN_76; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_153 = 2'h1 == io_router_req_bits_src_virt_id ? 1'h0 : _GEN_109; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_154 = 2'h1 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_0 : _GEN_93; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_155 = 2'h1 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_1 : _GEN_97; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_159 = 2'h1 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_1 : _GEN_81; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_162 = 2'h2 == io_router_req_bits_src_virt_id ? 1'h0 : _GEN_110; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_163 = 2'h2 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_0 : _GEN_94; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_164 = 2'h2 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_1 : _GEN_98; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_165 = 2'h2 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_2 : _GEN_102; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_168 = 2'h2 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_1 : _GEN_82; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_169 = 2'h2 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_2 : _GEN_86; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_171 = 2'h3 == io_router_req_bits_src_virt_id ? 1'h0 : _GEN_111; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_172 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_0 : _GEN_95; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_173 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_1 : _GEN_99; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_174 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_2 : _GEN_103; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_175 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_3 : _GEN_107; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_177 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_1 : _GEN_83; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_178 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_2 : _GEN_87; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_179 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_3 : _GEN_91; // @[InputUnit.scala 227:25 228:26]
  wire [2:0] _GEN_180 = io_router_req_valid ? _GEN_140 : _GEN_132; // @[InputUnit.scala 222:31]
  wire [2:0] _GEN_181 = io_router_req_valid ? _GEN_141 : _GEN_133; // @[InputUnit.scala 222:31]
  wire [2:0] _GEN_182 = io_router_req_valid ? _GEN_142 : _GEN_134; // @[InputUnit.scala 222:31]
  wire [2:0] _GEN_183 = io_router_req_valid ? _GEN_143 : _GEN_135; // @[InputUnit.scala 222:31]
  wire  _GEN_184 = io_router_req_valid ? _GEN_144 : _GEN_108; // @[InputUnit.scala 222:31]
  wire  _GEN_185 = io_router_req_valid ? _GEN_145 : _GEN_92; // @[InputUnit.scala 222:31]
  wire  _GEN_189 = io_router_req_valid ? _GEN_149 : _GEN_76; // @[InputUnit.scala 222:31]
  wire  _GEN_193 = io_router_req_valid ? _GEN_153 : _GEN_109; // @[InputUnit.scala 222:31]
  wire  _GEN_194 = io_router_req_valid ? _GEN_154 : _GEN_93; // @[InputUnit.scala 222:31]
  wire  _GEN_195 = io_router_req_valid ? _GEN_155 : _GEN_97; // @[InputUnit.scala 222:31]
  wire  _GEN_199 = io_router_req_valid ? _GEN_159 : _GEN_81; // @[InputUnit.scala 222:31]
  wire  _GEN_202 = io_router_req_valid ? _GEN_162 : _GEN_110; // @[InputUnit.scala 222:31]
  wire  _GEN_203 = io_router_req_valid ? _GEN_163 : _GEN_94; // @[InputUnit.scala 222:31]
  wire  _GEN_204 = io_router_req_valid ? _GEN_164 : _GEN_98; // @[InputUnit.scala 222:31]
  wire  _GEN_205 = io_router_req_valid ? _GEN_165 : _GEN_102; // @[InputUnit.scala 222:31]
  wire  _GEN_208 = io_router_req_valid ? _GEN_168 : _GEN_82; // @[InputUnit.scala 222:31]
  wire  _GEN_209 = io_router_req_valid ? _GEN_169 : _GEN_86; // @[InputUnit.scala 222:31]
  wire  _GEN_211 = io_router_req_valid ? _GEN_171 : _GEN_111; // @[InputUnit.scala 222:31]
  wire  _GEN_212 = io_router_req_valid ? _GEN_172 : _GEN_95; // @[InputUnit.scala 222:31]
  wire  _GEN_213 = io_router_req_valid ? _GEN_173 : _GEN_99; // @[InputUnit.scala 222:31]
  wire  _GEN_214 = io_router_req_valid ? _GEN_174 : _GEN_103; // @[InputUnit.scala 222:31]
  wire  _GEN_215 = io_router_req_valid ? _GEN_175 : _GEN_107; // @[InputUnit.scala 222:31]
  wire  _GEN_217 = io_router_req_valid ? _GEN_177 : _GEN_83; // @[InputUnit.scala 222:31]
  wire  _GEN_218 = io_router_req_valid ? _GEN_178 : _GEN_87; // @[InputUnit.scala 222:31]
  wire  _GEN_219 = io_router_req_valid ? _GEN_179 : _GEN_91; // @[InputUnit.scala 222:31]
  reg [3:0] mask; // @[InputUnit.scala 233:21]
  wire  vcalloc_vals_1 = states_1_g == 3'h2; // @[InputUnit.scala 249:32]
  wire  vcalloc_vals_0 = states_0_g == 3'h2; // @[InputUnit.scala 249:32]
  wire  vcalloc_vals_3 = states_3_g == 3'h2; // @[InputUnit.scala 249:32]
  wire  vcalloc_vals_2 = states_2_g == 3'h2; // @[InputUnit.scala 249:32]
  wire [3:0] _vcalloc_filter_T = {vcalloc_vals_3,vcalloc_vals_2,vcalloc_vals_1,vcalloc_vals_0}; // @[InputUnit.scala 236:59]
  wire [3:0] _vcalloc_filter_T_2 = ~mask; // @[InputUnit.scala 236:89]
  wire [3:0] _vcalloc_filter_T_3 = _vcalloc_filter_T & _vcalloc_filter_T_2; // @[InputUnit.scala 236:87]
  wire [7:0] _vcalloc_filter_T_4 = {vcalloc_vals_3,vcalloc_vals_2,vcalloc_vals_1,vcalloc_vals_0,_vcalloc_filter_T_3}; // @[Cat.scala 33:92]
  wire [7:0] _vcalloc_filter_T_13 = _vcalloc_filter_T_4[7] ? 8'h80 : 8'h0; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_14 = _vcalloc_filter_T_4[6] ? 8'h40 : _vcalloc_filter_T_13; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_15 = _vcalloc_filter_T_4[5] ? 8'h20 : _vcalloc_filter_T_14; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_16 = _vcalloc_filter_T_4[4] ? 8'h10 : _vcalloc_filter_T_15; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_17 = _vcalloc_filter_T_4[3] ? 8'h8 : _vcalloc_filter_T_16; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_18 = _vcalloc_filter_T_4[2] ? 8'h4 : _vcalloc_filter_T_17; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_19 = _vcalloc_filter_T_4[1] ? 8'h2 : _vcalloc_filter_T_18; // @[Mux.scala 47:70]
  wire [7:0] vcalloc_filter = _vcalloc_filter_T_4[0] ? 8'h1 : _vcalloc_filter_T_19; // @[Mux.scala 47:70]
  wire [3:0] vcalloc_sel = vcalloc_filter[3:0] | vcalloc_filter[7:4]; // @[InputUnit.scala 237:58]
  wire [3:0] _mask_T = 4'h1 << io_router_req_bits_src_virt_id; // @[InputUnit.scala 240:18]
  wire [3:0] _mask_T_2 = _mask_T - 4'h1; // @[InputUnit.scala 240:53]
  wire  _T_26 = vcalloc_vals_0 | vcalloc_vals_1 | vcalloc_vals_2 | vcalloc_vals_3; // @[package.scala 73:59]
  wire [1:0] _mask_T_12 = vcalloc_sel[1] ? 2'h3 : 2'h0; // @[Mux.scala 27:73]
  wire [2:0] _mask_T_13 = vcalloc_sel[2] ? 3'h7 : 3'h0; // @[Mux.scala 27:73]
  wire [3:0] _mask_T_14 = vcalloc_sel[3] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [1:0] _GEN_60 = {{1'd0}, vcalloc_sel[0]}; // @[Mux.scala 27:73]
  wire [1:0] _mask_T_15 = _GEN_60 | _mask_T_12; // @[Mux.scala 27:73]
  wire [2:0] _GEN_61 = {{1'd0}, _mask_T_15}; // @[Mux.scala 27:73]
  wire [2:0] _mask_T_16 = _GEN_61 | _mask_T_13; // @[Mux.scala 27:73]
  wire [3:0] _GEN_62 = {{1'd0}, _mask_T_16}; // @[Mux.scala 27:73]
  wire [3:0] _mask_T_17 = _GEN_62 | _mask_T_14; // @[Mux.scala 27:73]
  wire [2:0] _GEN_222 = vcalloc_vals_0 & vcalloc_sel[0] & io_vcalloc_req_ready ? 3'h3 : _GEN_180; // @[InputUnit.scala 253:{76,82}]
  wire [2:0] _GEN_223 = vcalloc_vals_1 & vcalloc_sel[1] & io_vcalloc_req_ready ? 3'h3 : _GEN_181; // @[InputUnit.scala 253:{76,82}]
  wire [2:0] _GEN_224 = vcalloc_vals_2 & vcalloc_sel[2] & io_vcalloc_req_ready ? 3'h3 : _GEN_182; // @[InputUnit.scala 253:{76,82}]
  wire [2:0] _GEN_225 = vcalloc_vals_3 & vcalloc_sel[3] & io_vcalloc_req_ready ? 3'h3 : _GEN_183; // @[InputUnit.scala 253:{76,82}]
  wire [1:0] _io_debug_va_stall_T = vcalloc_vals_0 + vcalloc_vals_1; // @[Bitwise.scala 51:90]
  wire [1:0] _io_debug_va_stall_T_2 = vcalloc_vals_2 + vcalloc_vals_3; // @[Bitwise.scala 51:90]
  wire [2:0] _io_debug_va_stall_T_4 = _io_debug_va_stall_T + _io_debug_va_stall_T_2; // @[Bitwise.scala 51:90]
  wire [2:0] _GEN_63 = {{2'd0}, io_vcalloc_req_ready}; // @[InputUnit.scala 266:47]
  wire [2:0] _io_debug_va_stall_T_7 = _io_debug_va_stall_T_4 - _GEN_63; // @[InputUnit.scala 266:47]
  wire  _T_39 = io_vcalloc_req_ready & io_vcalloc_req_valid; // @[Decoupled.scala 51:35]
  wire [8:0] _credit_available_T = {states_0_vc_sel_2_0,1'h0,1'h0,1'h0,states_0_vc_sel_1_0,2'h0,1'h0,states_0_vc_sel_0_0
    }; // @[InputUnit.scala 287:40]
  wire [8:0] _credit_available_T_1 = {io_out_credit_available_2_0,io_out_credit_available_1_3,
    io_out_credit_available_1_2,io_out_credit_available_1_1,io_out_credit_available_1_0,io_out_credit_available_0_3,
    io_out_credit_available_0_2,io_out_credit_available_0_1,io_out_credit_available_0_0}; // @[InputUnit.scala 287:73]
  wire [8:0] _credit_available_T_2 = _credit_available_T & _credit_available_T_1; // @[InputUnit.scala 287:47]
  wire  credit_available = _credit_available_T_2 != 9'h0; // @[InputUnit.scala 287:81]
  wire  _T_60 = salloc_arb_io_in_0_ready & salloc_arb_io_in_0_valid; // @[Decoupled.scala 51:35]
  wire [8:0] _credit_available_T_3 = {states_1_vc_sel_2_0,1'h0,1'h0,states_1_vc_sel_1_1,states_1_vc_sel_1_0,2'h0,
    states_1_vc_sel_0_1,1'h0}; // @[InputUnit.scala 287:40]
  wire [8:0] _credit_available_T_5 = _credit_available_T_3 & _credit_available_T_1; // @[InputUnit.scala 287:47]
  wire  credit_available_1 = _credit_available_T_5 != 9'h0; // @[InputUnit.scala 287:81]
  wire  _T_62 = salloc_arb_io_in_1_ready & salloc_arb_io_in_1_valid; // @[Decoupled.scala 51:35]
  wire [8:0] _credit_available_T_6 = {states_2_vc_sel_2_0,1'h0,states_2_vc_sel_1_2,states_2_vc_sel_1_1,
    states_2_vc_sel_1_0,1'h0,states_2_vc_sel_0_2,states_2_vc_sel_0_1,1'h0}; // @[InputUnit.scala 287:40]
  wire [8:0] _credit_available_T_8 = _credit_available_T_6 & _credit_available_T_1; // @[InputUnit.scala 287:47]
  wire  credit_available_2 = _credit_available_T_8 != 9'h0; // @[InputUnit.scala 287:81]
  wire  _T_64 = salloc_arb_io_in_2_ready & salloc_arb_io_in_2_valid; // @[Decoupled.scala 51:35]
  wire [8:0] _credit_available_T_9 = {states_3_vc_sel_2_0,states_3_vc_sel_1_3,states_3_vc_sel_1_2,states_3_vc_sel_1_1,
    states_3_vc_sel_1_0,states_3_vc_sel_0_3,states_3_vc_sel_0_2,states_3_vc_sel_0_1,1'h0}; // @[InputUnit.scala 287:40]
  wire [8:0] _credit_available_T_11 = _credit_available_T_9 & _credit_available_T_1; // @[InputUnit.scala 287:47]
  wire  credit_available_3 = _credit_available_T_11 != 9'h0; // @[InputUnit.scala 287:81]
  wire  _T_66 = salloc_arb_io_in_3_ready & salloc_arb_io_in_3_valid; // @[Decoupled.scala 51:35]
  wire  _io_debug_sa_stall_T_1 = salloc_arb_io_in_0_valid & ~salloc_arb_io_in_0_ready; // @[InputUnit.scala 301:67]
  wire  _io_debug_sa_stall_T_3 = salloc_arb_io_in_1_valid & ~salloc_arb_io_in_1_ready; // @[InputUnit.scala 301:67]
  wire  _io_debug_sa_stall_T_5 = salloc_arb_io_in_2_valid & ~salloc_arb_io_in_2_ready; // @[InputUnit.scala 301:67]
  wire  _io_debug_sa_stall_T_7 = salloc_arb_io_in_3_valid & ~salloc_arb_io_in_3_ready; // @[InputUnit.scala 301:67]
  wire [1:0] _io_debug_sa_stall_T_8 = _io_debug_sa_stall_T_1 + _io_debug_sa_stall_T_3; // @[Bitwise.scala 51:90]
  wire [1:0] _io_debug_sa_stall_T_10 = _io_debug_sa_stall_T_5 + _io_debug_sa_stall_T_7; // @[Bitwise.scala 51:90]
  wire [2:0] _io_debug_sa_stall_T_12 = _io_debug_sa_stall_T_8 + _io_debug_sa_stall_T_10; // @[Bitwise.scala 51:90]
  reg  salloc_outs_0_valid; // @[InputUnit.scala 318:8]
  reg [1:0] salloc_outs_0_out_vid; // @[InputUnit.scala 318:8]
  reg  salloc_outs_0_flit_head; // @[InputUnit.scala 318:8]
  reg  salloc_outs_0_flit_tail; // @[InputUnit.scala 318:8]
  reg [63:0] salloc_outs_0_flit_payload; // @[InputUnit.scala 318:8]
  reg [1:0] salloc_outs_0_flit_flow_ingress_node; // @[InputUnit.scala 318:8]
  reg [1:0] salloc_outs_0_flit_flow_egress_node; // @[InputUnit.scala 318:8]
  wire  _io_in_credit_return_T = salloc_arb_io_out_0_ready & salloc_arb_io_out_0_valid; // @[Decoupled.scala 51:35]
  wire  _io_in_vc_free_T_11 = salloc_arb_io_chosen_oh_0[0] & input_buffer_io_deq_0_bits_tail | salloc_arb_io_chosen_oh_0
    [1] & input_buffer_io_deq_1_bits_tail | salloc_arb_io_chosen_oh_0[2] & input_buffer_io_deq_2_bits_tail |
    salloc_arb_io_chosen_oh_0[3] & input_buffer_io_deq_3_bits_tail; // @[Mux.scala 27:73]
  wire  vc_sel_0_0 = salloc_arb_io_chosen_oh_0[0] & states_0_vc_sel_0_0; // @[Mux.scala 27:73]
  wire  vc_sel_0_1 = salloc_arb_io_chosen_oh_0[1] & states_1_vc_sel_0_1 | salloc_arb_io_chosen_oh_0[2] &
    states_2_vc_sel_0_1 | salloc_arb_io_chosen_oh_0[3] & states_3_vc_sel_0_1; // @[Mux.scala 27:73]
  wire  vc_sel_0_2 = salloc_arb_io_chosen_oh_0[2] & states_2_vc_sel_0_2 | salloc_arb_io_chosen_oh_0[3] &
    states_3_vc_sel_0_2; // @[Mux.scala 27:73]
  wire  vc_sel_0_3 = salloc_arb_io_chosen_oh_0[3] & states_3_vc_sel_0_3; // @[Mux.scala 27:73]
  wire  vc_sel_1_0 = salloc_arb_io_chosen_oh_0[0] & states_0_vc_sel_1_0 | salloc_arb_io_chosen_oh_0[1] &
    states_1_vc_sel_1_0 | salloc_arb_io_chosen_oh_0[2] & states_2_vc_sel_1_0 | salloc_arb_io_chosen_oh_0[3] &
    states_3_vc_sel_1_0; // @[Mux.scala 27:73]
  wire  vc_sel_1_1 = salloc_arb_io_chosen_oh_0[1] & states_1_vc_sel_1_1 | salloc_arb_io_chosen_oh_0[2] &
    states_2_vc_sel_1_1 | salloc_arb_io_chosen_oh_0[3] & states_3_vc_sel_1_1; // @[Mux.scala 27:73]
  wire  vc_sel_1_2 = salloc_arb_io_chosen_oh_0[2] & states_2_vc_sel_1_2 | salloc_arb_io_chosen_oh_0[3] &
    states_3_vc_sel_1_2; // @[Mux.scala 27:73]
  wire  vc_sel_1_3 = salloc_arb_io_chosen_oh_0[3] & states_3_vc_sel_1_3; // @[Mux.scala 27:73]
  wire  channel_oh_0 = vc_sel_0_0 | vc_sel_0_1 | vc_sel_0_2 | vc_sel_0_3; // @[InputUnit.scala 334:43]
  wire  channel_oh_1 = vc_sel_1_0 | vc_sel_1_1 | vc_sel_1_2 | vc_sel_1_3; // @[InputUnit.scala 334:43]
  wire [3:0] _virt_channel_T = {vc_sel_0_3,vc_sel_0_2,vc_sel_0_1,vc_sel_0_0}; // @[OneHot.scala 22:45]
  wire [1:0] virt_channel_hi_1 = _virt_channel_T[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] virt_channel_lo_1 = _virt_channel_T[1:0]; // @[OneHot.scala 31:18]
  wire  _virt_channel_T_1 = |virt_channel_hi_1; // @[OneHot.scala 32:14]
  wire [1:0] _virt_channel_T_2 = virt_channel_hi_1 | virt_channel_lo_1; // @[OneHot.scala 32:28]
  wire [1:0] _virt_channel_T_4 = {_virt_channel_T_1,_virt_channel_T_2[1]}; // @[Cat.scala 33:92]
  wire [3:0] _virt_channel_T_5 = {vc_sel_1_3,vc_sel_1_2,vc_sel_1_1,vc_sel_1_0}; // @[OneHot.scala 22:45]
  wire [1:0] virt_channel_hi_3 = _virt_channel_T_5[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] virt_channel_lo_3 = _virt_channel_T_5[1:0]; // @[OneHot.scala 31:18]
  wire  _virt_channel_T_6 = |virt_channel_hi_3; // @[OneHot.scala 32:14]
  wire [1:0] _virt_channel_T_7 = virt_channel_hi_3 | virt_channel_lo_3; // @[OneHot.scala 32:28]
  wire [1:0] _virt_channel_T_9 = {_virt_channel_T_6,_virt_channel_T_7[1]}; // @[Cat.scala 33:92]
  wire [1:0] _virt_channel_T_10 = channel_oh_0 ? _virt_channel_T_4 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _virt_channel_T_11 = channel_oh_1 ? _virt_channel_T_9 : 2'h0; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_4 = salloc_arb_io_chosen_oh_0[0] ? input_buffer_io_deq_0_bits_payload : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_5 = salloc_arb_io_chosen_oh_0[1] ? input_buffer_io_deq_1_bits_payload : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_6 = salloc_arb_io_chosen_oh_0[2] ? input_buffer_io_deq_2_bits_payload : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_7 = salloc_arb_io_chosen_oh_0[3] ? input_buffer_io_deq_3_bits_payload : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_8 = _salloc_outs_0_flit_payload_T_4 | _salloc_outs_0_flit_payload_T_5; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_9 = _salloc_outs_0_flit_payload_T_8 | _salloc_outs_0_flit_payload_T_6; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_11 = salloc_arb_io_chosen_oh_0[0] ? states_0_flow_egress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_12 = salloc_arb_io_chosen_oh_0[1] ? states_1_flow_egress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_13 = salloc_arb_io_chosen_oh_0[2] ? states_2_flow_egress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_14 = salloc_arb_io_chosen_oh_0[3] ? states_3_flow_egress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_15 = _salloc_outs_0_flit_flow_T_11 | _salloc_outs_0_flit_flow_T_12; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_16 = _salloc_outs_0_flit_flow_T_15 | _salloc_outs_0_flit_flow_T_13; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_25 = salloc_arb_io_chosen_oh_0[0] ? states_0_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_26 = salloc_arb_io_chosen_oh_0[1] ? states_1_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_27 = salloc_arb_io_chosen_oh_0[2] ? states_2_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_28 = salloc_arb_io_chosen_oh_0[3] ? states_3_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_29 = _salloc_outs_0_flit_flow_T_25 | _salloc_outs_0_flit_flow_T_26; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_30 = _salloc_outs_0_flit_flow_T_29 | _salloc_outs_0_flit_flow_T_27; // @[Mux.scala 27:73]
  InputBuffer input_buffer ( // @[InputUnit.scala 180:28]
    .clock(input_buffer_clock),
    .reset(input_buffer_reset),
    .io_enq_0_valid(input_buffer_io_enq_0_valid),
    .io_enq_0_bits_head(input_buffer_io_enq_0_bits_head),
    .io_enq_0_bits_tail(input_buffer_io_enq_0_bits_tail),
    .io_enq_0_bits_payload(input_buffer_io_enq_0_bits_payload),
    .io_enq_0_bits_virt_channel_id(input_buffer_io_enq_0_bits_virt_channel_id),
    .io_deq_0_ready(input_buffer_io_deq_0_ready),
    .io_deq_0_valid(input_buffer_io_deq_0_valid),
    .io_deq_0_bits_head(input_buffer_io_deq_0_bits_head),
    .io_deq_0_bits_tail(input_buffer_io_deq_0_bits_tail),
    .io_deq_0_bits_payload(input_buffer_io_deq_0_bits_payload),
    .io_deq_1_ready(input_buffer_io_deq_1_ready),
    .io_deq_1_valid(input_buffer_io_deq_1_valid),
    .io_deq_1_bits_head(input_buffer_io_deq_1_bits_head),
    .io_deq_1_bits_tail(input_buffer_io_deq_1_bits_tail),
    .io_deq_1_bits_payload(input_buffer_io_deq_1_bits_payload),
    .io_deq_2_ready(input_buffer_io_deq_2_ready),
    .io_deq_2_valid(input_buffer_io_deq_2_valid),
    .io_deq_2_bits_head(input_buffer_io_deq_2_bits_head),
    .io_deq_2_bits_tail(input_buffer_io_deq_2_bits_tail),
    .io_deq_2_bits_payload(input_buffer_io_deq_2_bits_payload),
    .io_deq_3_ready(input_buffer_io_deq_3_ready),
    .io_deq_3_valid(input_buffer_io_deq_3_valid),
    .io_deq_3_bits_head(input_buffer_io_deq_3_bits_head),
    .io_deq_3_bits_tail(input_buffer_io_deq_3_bits_tail),
    .io_deq_3_bits_payload(input_buffer_io_deq_3_bits_payload)
  );
  Arbiter route_arbiter ( // @[InputUnit.scala 186:29]
    .io_in_0_valid(route_arbiter_io_in_0_valid),
    .io_in_0_bits_flow_ingress_node(route_arbiter_io_in_0_bits_flow_ingress_node),
    .io_in_0_bits_flow_egress_node(route_arbiter_io_in_0_bits_flow_egress_node),
    .io_in_1_ready(route_arbiter_io_in_1_ready),
    .io_in_1_valid(route_arbiter_io_in_1_valid),
    .io_in_1_bits_flow_ingress_node(route_arbiter_io_in_1_bits_flow_ingress_node),
    .io_in_1_bits_flow_egress_node(route_arbiter_io_in_1_bits_flow_egress_node),
    .io_in_2_ready(route_arbiter_io_in_2_ready),
    .io_in_2_valid(route_arbiter_io_in_2_valid),
    .io_in_2_bits_flow_ingress_node(route_arbiter_io_in_2_bits_flow_ingress_node),
    .io_in_2_bits_flow_egress_node(route_arbiter_io_in_2_bits_flow_egress_node),
    .io_in_3_ready(route_arbiter_io_in_3_ready),
    .io_in_3_valid(route_arbiter_io_in_3_valid),
    .io_in_3_bits_flow_ingress_node(route_arbiter_io_in_3_bits_flow_ingress_node),
    .io_in_3_bits_flow_egress_node(route_arbiter_io_in_3_bits_flow_egress_node),
    .io_out_valid(route_arbiter_io_out_valid),
    .io_out_bits_src_virt_id(route_arbiter_io_out_bits_src_virt_id),
    .io_out_bits_flow_ingress_node(route_arbiter_io_out_bits_flow_ingress_node),
    .io_out_bits_flow_egress_node(route_arbiter_io_out_bits_flow_egress_node)
  );
  SwitchArbiter salloc_arb ( // @[InputUnit.scala 279:26]
    .clock(salloc_arb_clock),
    .reset(salloc_arb_reset),
    .io_in_0_ready(salloc_arb_io_in_0_ready),
    .io_in_0_valid(salloc_arb_io_in_0_valid),
    .io_in_0_bits_vc_sel_2_0(salloc_arb_io_in_0_bits_vc_sel_2_0),
    .io_in_0_bits_vc_sel_1_0(salloc_arb_io_in_0_bits_vc_sel_1_0),
    .io_in_0_bits_vc_sel_0_0(salloc_arb_io_in_0_bits_vc_sel_0_0),
    .io_in_0_bits_tail(salloc_arb_io_in_0_bits_tail),
    .io_in_1_ready(salloc_arb_io_in_1_ready),
    .io_in_1_valid(salloc_arb_io_in_1_valid),
    .io_in_1_bits_vc_sel_2_0(salloc_arb_io_in_1_bits_vc_sel_2_0),
    .io_in_1_bits_vc_sel_1_0(salloc_arb_io_in_1_bits_vc_sel_1_0),
    .io_in_1_bits_vc_sel_1_1(salloc_arb_io_in_1_bits_vc_sel_1_1),
    .io_in_1_bits_vc_sel_0_0(salloc_arb_io_in_1_bits_vc_sel_0_0),
    .io_in_1_bits_vc_sel_0_1(salloc_arb_io_in_1_bits_vc_sel_0_1),
    .io_in_1_bits_tail(salloc_arb_io_in_1_bits_tail),
    .io_in_2_ready(salloc_arb_io_in_2_ready),
    .io_in_2_valid(salloc_arb_io_in_2_valid),
    .io_in_2_bits_vc_sel_2_0(salloc_arb_io_in_2_bits_vc_sel_2_0),
    .io_in_2_bits_vc_sel_1_0(salloc_arb_io_in_2_bits_vc_sel_1_0),
    .io_in_2_bits_vc_sel_1_1(salloc_arb_io_in_2_bits_vc_sel_1_1),
    .io_in_2_bits_vc_sel_1_2(salloc_arb_io_in_2_bits_vc_sel_1_2),
    .io_in_2_bits_vc_sel_0_0(salloc_arb_io_in_2_bits_vc_sel_0_0),
    .io_in_2_bits_vc_sel_0_1(salloc_arb_io_in_2_bits_vc_sel_0_1),
    .io_in_2_bits_vc_sel_0_2(salloc_arb_io_in_2_bits_vc_sel_0_2),
    .io_in_2_bits_tail(salloc_arb_io_in_2_bits_tail),
    .io_in_3_ready(salloc_arb_io_in_3_ready),
    .io_in_3_valid(salloc_arb_io_in_3_valid),
    .io_in_3_bits_vc_sel_2_0(salloc_arb_io_in_3_bits_vc_sel_2_0),
    .io_in_3_bits_vc_sel_1_0(salloc_arb_io_in_3_bits_vc_sel_1_0),
    .io_in_3_bits_vc_sel_1_1(salloc_arb_io_in_3_bits_vc_sel_1_1),
    .io_in_3_bits_vc_sel_1_2(salloc_arb_io_in_3_bits_vc_sel_1_2),
    .io_in_3_bits_vc_sel_1_3(salloc_arb_io_in_3_bits_vc_sel_1_3),
    .io_in_3_bits_vc_sel_0_0(salloc_arb_io_in_3_bits_vc_sel_0_0),
    .io_in_3_bits_vc_sel_0_1(salloc_arb_io_in_3_bits_vc_sel_0_1),
    .io_in_3_bits_vc_sel_0_2(salloc_arb_io_in_3_bits_vc_sel_0_2),
    .io_in_3_bits_vc_sel_0_3(salloc_arb_io_in_3_bits_vc_sel_0_3),
    .io_in_3_bits_tail(salloc_arb_io_in_3_bits_tail),
    .io_out_0_ready(salloc_arb_io_out_0_ready),
    .io_out_0_valid(salloc_arb_io_out_0_valid),
    .io_out_0_bits_vc_sel_2_0(salloc_arb_io_out_0_bits_vc_sel_2_0),
    .io_out_0_bits_vc_sel_1_0(salloc_arb_io_out_0_bits_vc_sel_1_0),
    .io_out_0_bits_vc_sel_1_1(salloc_arb_io_out_0_bits_vc_sel_1_1),
    .io_out_0_bits_vc_sel_1_2(salloc_arb_io_out_0_bits_vc_sel_1_2),
    .io_out_0_bits_vc_sel_1_3(salloc_arb_io_out_0_bits_vc_sel_1_3),
    .io_out_0_bits_vc_sel_0_0(salloc_arb_io_out_0_bits_vc_sel_0_0),
    .io_out_0_bits_vc_sel_0_1(salloc_arb_io_out_0_bits_vc_sel_0_1),
    .io_out_0_bits_vc_sel_0_2(salloc_arb_io_out_0_bits_vc_sel_0_2),
    .io_out_0_bits_vc_sel_0_3(salloc_arb_io_out_0_bits_vc_sel_0_3),
    .io_out_0_bits_tail(salloc_arb_io_out_0_bits_tail),
    .io_chosen_oh_0(salloc_arb_io_chosen_oh_0)
  );
  assign io_router_req_valid = route_arbiter_io_out_valid; // @[InputUnit.scala 189:17]
  assign io_router_req_bits_src_virt_id = route_arbiter_io_out_bits_src_virt_id; // @[InputUnit.scala 189:17]
  assign io_router_req_bits_flow_ingress_node = route_arbiter_io_out_bits_flow_ingress_node; // @[InputUnit.scala 189:17]
  assign io_router_req_bits_flow_egress_node = route_arbiter_io_out_bits_flow_egress_node; // @[InputUnit.scala 189:17]
  assign io_vcalloc_req_valid = vcalloc_vals_0 | vcalloc_vals_1 | vcalloc_vals_2 | vcalloc_vals_3; // @[package.scala 73:59]
  assign io_vcalloc_req_bits_vc_sel_2_0 = vcalloc_sel[0] & states_0_vc_sel_2_0 | vcalloc_sel[1] & states_1_vc_sel_2_0 |
    vcalloc_sel[2] & states_2_vc_sel_2_0 | vcalloc_sel[3] & states_3_vc_sel_2_0; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_1_0 = vcalloc_sel[0] & states_0_vc_sel_1_0 | vcalloc_sel[1] & states_1_vc_sel_1_0 |
    vcalloc_sel[2] & states_2_vc_sel_1_0 | vcalloc_sel[3] & states_3_vc_sel_1_0; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_1_1 = vcalloc_sel[1] & states_1_vc_sel_1_1 | vcalloc_sel[2] & states_2_vc_sel_1_1 |
    vcalloc_sel[3] & states_3_vc_sel_1_1; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_1_2 = vcalloc_sel[2] & states_2_vc_sel_1_2 | vcalloc_sel[3] & states_3_vc_sel_1_2; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_1_3 = vcalloc_sel[3] & states_3_vc_sel_1_3; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_0_0 = vcalloc_sel[0] & states_0_vc_sel_0_0; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_0_1 = vcalloc_sel[1] & states_1_vc_sel_0_1 | vcalloc_sel[2] & states_2_vc_sel_0_1 |
    vcalloc_sel[3] & states_3_vc_sel_0_1; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_0_2 = vcalloc_sel[2] & states_2_vc_sel_0_2 | vcalloc_sel[3] & states_3_vc_sel_0_2; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_0_3 = vcalloc_sel[3] & states_3_vc_sel_0_3; // @[Mux.scala 27:73]
  assign io_salloc_req_0_valid = salloc_arb_io_out_0_valid; // @[InputUnit.scala 302:17 303:19 305:35]
  assign io_salloc_req_0_bits_vc_sel_2_0 = salloc_arb_io_out_0_bits_vc_sel_2_0; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_1_0 = salloc_arb_io_out_0_bits_vc_sel_1_0; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_1_1 = salloc_arb_io_out_0_bits_vc_sel_1_1; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_1_2 = salloc_arb_io_out_0_bits_vc_sel_1_2; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_1_3 = salloc_arb_io_out_0_bits_vc_sel_1_3; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_0_0 = salloc_arb_io_out_0_bits_vc_sel_0_0; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_0_1 = salloc_arb_io_out_0_bits_vc_sel_0_1; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_0_2 = salloc_arb_io_out_0_bits_vc_sel_0_2; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_0_3 = salloc_arb_io_out_0_bits_vc_sel_0_3; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_tail = salloc_arb_io_out_0_bits_tail; // @[InputUnit.scala 302:17]
  assign io_out_0_valid = salloc_outs_0_valid; // @[InputUnit.scala 349:21]
  assign io_out_0_bits_flit_head = salloc_outs_0_flit_head; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_flit_tail = salloc_outs_0_flit_tail; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_flit_payload = salloc_outs_0_flit_payload; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_flit_flow_ingress_node = salloc_outs_0_flit_flow_ingress_node; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_flit_flow_egress_node = salloc_outs_0_flit_flow_egress_node; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_out_virt_channel = salloc_outs_0_out_vid; // @[InputUnit.scala 351:37]
  assign io_debug_va_stall = _io_debug_va_stall_T_7[1:0]; // @[InputUnit.scala 266:21]
  assign io_debug_sa_stall = _io_debug_sa_stall_T_12[1:0]; // @[InputUnit.scala 301:21]
  assign io_in_credit_return = _io_in_credit_return_T ? salloc_arb_io_chosen_oh_0 : 4'h0; // @[InputUnit.scala 322:8]
  assign io_in_vc_free = _io_in_credit_return_T & _io_in_vc_free_T_11 ? salloc_arb_io_chosen_oh_0 : 4'h0; // @[InputUnit.scala 325:8]
  assign input_buffer_clock = clock;
  assign input_buffer_reset = reset;
  assign input_buffer_io_enq_0_valid = io_in_flit_0_valid; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_head = io_in_flit_0_bits_head; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_tail = io_in_flit_0_bits_tail; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_payload = io_in_flit_0_bits_payload; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_virt_channel_id = io_in_flit_0_bits_virt_channel_id; // @[InputUnit.scala 182:28]
  assign input_buffer_io_deq_0_ready = salloc_arb_io_in_0_ready; // @[InputUnit.scala 295:36]
  assign input_buffer_io_deq_1_ready = salloc_arb_io_in_1_ready; // @[InputUnit.scala 295:36]
  assign input_buffer_io_deq_2_ready = salloc_arb_io_in_2_ready; // @[InputUnit.scala 295:36]
  assign input_buffer_io_deq_3_ready = salloc_arb_io_in_3_ready; // @[InputUnit.scala 295:36]
  assign route_arbiter_io_in_0_valid = states_0_g == 3'h1; // @[InputUnit.scala 212:22]
  assign route_arbiter_io_in_0_bits_flow_ingress_node = states_0_flow_ingress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_0_bits_flow_egress_node = states_0_flow_egress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_1_valid = states_1_g == 3'h1; // @[InputUnit.scala 212:22]
  assign route_arbiter_io_in_1_bits_flow_ingress_node = states_1_flow_ingress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_1_bits_flow_egress_node = states_1_flow_egress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_2_valid = states_2_g == 3'h1; // @[InputUnit.scala 212:22]
  assign route_arbiter_io_in_2_bits_flow_ingress_node = states_2_flow_ingress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_2_bits_flow_egress_node = states_2_flow_egress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_3_valid = states_3_g == 3'h1; // @[InputUnit.scala 212:22]
  assign route_arbiter_io_in_3_bits_flow_ingress_node = states_3_flow_ingress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_3_bits_flow_egress_node = states_3_flow_egress_node; // @[InputUnit.scala 213:19]
  assign salloc_arb_clock = clock;
  assign salloc_arb_reset = reset;
  assign salloc_arb_io_in_0_valid = states_0_g == 3'h3 & credit_available & input_buffer_io_deq_0_valid; // @[InputUnit.scala 288:50]
  assign salloc_arb_io_in_0_bits_vc_sel_2_0 = states_0_vc_sel_2_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_0_bits_vc_sel_1_0 = states_0_vc_sel_1_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_0_bits_vc_sel_0_0 = states_0_vc_sel_0_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_0_bits_tail = input_buffer_io_deq_0_bits_tail; // @[InputUnit.scala 291:19]
  assign salloc_arb_io_in_1_valid = states_1_g == 3'h3 & credit_available_1 & input_buffer_io_deq_1_valid; // @[InputUnit.scala 288:50]
  assign salloc_arb_io_in_1_bits_vc_sel_2_0 = states_1_vc_sel_2_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_1_bits_vc_sel_1_0 = states_1_vc_sel_1_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_1_bits_vc_sel_1_1 = states_1_vc_sel_1_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_1_bits_vc_sel_0_0 = 1'h0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_1_bits_vc_sel_0_1 = states_1_vc_sel_0_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_1_bits_tail = input_buffer_io_deq_1_bits_tail; // @[InputUnit.scala 291:19]
  assign salloc_arb_io_in_2_valid = states_2_g == 3'h3 & credit_available_2 & input_buffer_io_deq_2_valid; // @[InputUnit.scala 288:50]
  assign salloc_arb_io_in_2_bits_vc_sel_2_0 = states_2_vc_sel_2_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_1_0 = states_2_vc_sel_1_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_1_1 = states_2_vc_sel_1_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_1_2 = states_2_vc_sel_1_2; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_0_0 = 1'h0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_0_1 = states_2_vc_sel_0_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_0_2 = states_2_vc_sel_0_2; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_tail = input_buffer_io_deq_2_bits_tail; // @[InputUnit.scala 291:19]
  assign salloc_arb_io_in_3_valid = states_3_g == 3'h3 & credit_available_3 & input_buffer_io_deq_3_valid; // @[InputUnit.scala 288:50]
  assign salloc_arb_io_in_3_bits_vc_sel_2_0 = states_3_vc_sel_2_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_1_0 = states_3_vc_sel_1_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_1_1 = states_3_vc_sel_1_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_1_2 = states_3_vc_sel_1_2; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_1_3 = states_3_vc_sel_1_3; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_0_0 = 1'h0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_0_1 = states_3_vc_sel_0_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_0_2 = states_3_vc_sel_0_2; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_0_3 = states_3_vc_sel_0_3; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_tail = input_buffer_io_deq_3_bits_tail; // @[InputUnit.scala 291:19]
  assign salloc_arb_io_out_0_ready = io_salloc_req_0_ready; // @[InputUnit.scala 302:17 303:19 304:39]
  always @(posedge clock) begin
    if (reset) begin // @[InputUnit.scala 377:23]
      states_0_g <= 3'h0; // @[InputUnit.scala 378:24]
    end else if (_T_60 & input_buffer_io_deq_0_bits_tail) begin // @[InputUnit.scala 292:35]
      states_0_g <= 3'h0; // @[InputUnit.scala 293:13]
    end else if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[0]) begin // @[InputUnit.scala 270:29]
        states_0_g <= 3'h3; // @[InputUnit.scala 272:21]
      end else begin
        states_0_g <= _GEN_222;
      end
    end else begin
      states_0_g <= _GEN_222;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[0]) begin // @[InputUnit.scala 270:29]
        states_0_vc_sel_2_0 <= io_vcalloc_resp_vc_sel_2_0; // @[InputUnit.scala 271:26]
      end else begin
        states_0_vc_sel_2_0 <= _GEN_184;
      end
    end else begin
      states_0_vc_sel_2_0 <= _GEN_184;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[0]) begin // @[InputUnit.scala 270:29]
        states_0_vc_sel_1_0 <= io_vcalloc_resp_vc_sel_1_0; // @[InputUnit.scala 271:26]
      end else begin
        states_0_vc_sel_1_0 <= _GEN_185;
      end
    end else begin
      states_0_vc_sel_1_0 <= _GEN_185;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[0]) begin // @[InputUnit.scala 270:29]
        states_0_vc_sel_0_0 <= io_vcalloc_resp_vc_sel_0_0; // @[InputUnit.scala 271:26]
      end else begin
        states_0_vc_sel_0_0 <= _GEN_189;
      end
    end else begin
      states_0_vc_sel_0_0 <= _GEN_189;
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h0 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_0_flow_ingress_node <= io_in_flit_0_bits_flow_ingress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h0 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_0_flow_egress_node <= io_in_flit_0_bits_flow_egress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (reset) begin // @[InputUnit.scala 377:23]
      states_1_g <= 3'h0; // @[InputUnit.scala 378:24]
    end else if (_T_62 & input_buffer_io_deq_1_bits_tail) begin // @[InputUnit.scala 292:35]
      states_1_g <= 3'h0; // @[InputUnit.scala 293:13]
    end else if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_g <= 3'h3; // @[InputUnit.scala 272:21]
      end else begin
        states_1_g <= _GEN_223;
      end
    end else begin
      states_1_g <= _GEN_223;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_vc_sel_2_0 <= io_vcalloc_resp_vc_sel_2_0; // @[InputUnit.scala 271:26]
      end else begin
        states_1_vc_sel_2_0 <= _GEN_193;
      end
    end else begin
      states_1_vc_sel_2_0 <= _GEN_193;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_vc_sel_1_0 <= io_vcalloc_resp_vc_sel_1_0; // @[InputUnit.scala 271:26]
      end else begin
        states_1_vc_sel_1_0 <= _GEN_194;
      end
    end else begin
      states_1_vc_sel_1_0 <= _GEN_194;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_vc_sel_1_1 <= io_vcalloc_resp_vc_sel_1_1; // @[InputUnit.scala 271:26]
      end else begin
        states_1_vc_sel_1_1 <= _GEN_195;
      end
    end else begin
      states_1_vc_sel_1_1 <= _GEN_195;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_vc_sel_0_1 <= io_vcalloc_resp_vc_sel_0_1; // @[InputUnit.scala 271:26]
      end else begin
        states_1_vc_sel_0_1 <= _GEN_199;
      end
    end else begin
      states_1_vc_sel_0_1 <= _GEN_199;
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h1 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_1_flow_ingress_node <= io_in_flit_0_bits_flow_ingress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h1 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_1_flow_egress_node <= io_in_flit_0_bits_flow_egress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (reset) begin // @[InputUnit.scala 377:23]
      states_2_g <= 3'h0; // @[InputUnit.scala 378:24]
    end else if (_T_64 & input_buffer_io_deq_2_bits_tail) begin // @[InputUnit.scala 292:35]
      states_2_g <= 3'h0; // @[InputUnit.scala 293:13]
    end else if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_g <= 3'h3; // @[InputUnit.scala 272:21]
      end else begin
        states_2_g <= _GEN_224;
      end
    end else begin
      states_2_g <= _GEN_224;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_2_0 <= io_vcalloc_resp_vc_sel_2_0; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_2_0 <= _GEN_202;
      end
    end else begin
      states_2_vc_sel_2_0 <= _GEN_202;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_1_0 <= io_vcalloc_resp_vc_sel_1_0; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_1_0 <= _GEN_203;
      end
    end else begin
      states_2_vc_sel_1_0 <= _GEN_203;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_1_1 <= io_vcalloc_resp_vc_sel_1_1; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_1_1 <= _GEN_204;
      end
    end else begin
      states_2_vc_sel_1_1 <= _GEN_204;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_1_2 <= io_vcalloc_resp_vc_sel_1_2; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_1_2 <= _GEN_205;
      end
    end else begin
      states_2_vc_sel_1_2 <= _GEN_205;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_0_1 <= io_vcalloc_resp_vc_sel_0_1; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_0_1 <= _GEN_208;
      end
    end else begin
      states_2_vc_sel_0_1 <= _GEN_208;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_0_2 <= io_vcalloc_resp_vc_sel_0_2; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_0_2 <= _GEN_209;
      end
    end else begin
      states_2_vc_sel_0_2 <= _GEN_209;
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h2 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_2_flow_ingress_node <= io_in_flit_0_bits_flow_ingress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h2 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_2_flow_egress_node <= io_in_flit_0_bits_flow_egress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (reset) begin // @[InputUnit.scala 377:23]
      states_3_g <= 3'h0; // @[InputUnit.scala 378:24]
    end else if (_T_66 & input_buffer_io_deq_3_bits_tail) begin // @[InputUnit.scala 292:35]
      states_3_g <= 3'h0; // @[InputUnit.scala 293:13]
    end else if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_g <= 3'h3; // @[InputUnit.scala 272:21]
      end else begin
        states_3_g <= _GEN_225;
      end
    end else begin
      states_3_g <= _GEN_225;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_2_0 <= io_vcalloc_resp_vc_sel_2_0; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_2_0 <= _GEN_211;
      end
    end else begin
      states_3_vc_sel_2_0 <= _GEN_211;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_1_0 <= io_vcalloc_resp_vc_sel_1_0; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_1_0 <= _GEN_212;
      end
    end else begin
      states_3_vc_sel_1_0 <= _GEN_212;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_1_1 <= io_vcalloc_resp_vc_sel_1_1; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_1_1 <= _GEN_213;
      end
    end else begin
      states_3_vc_sel_1_1 <= _GEN_213;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_1_2 <= io_vcalloc_resp_vc_sel_1_2; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_1_2 <= _GEN_214;
      end
    end else begin
      states_3_vc_sel_1_2 <= _GEN_214;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_1_3 <= io_vcalloc_resp_vc_sel_1_3; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_1_3 <= _GEN_215;
      end
    end else begin
      states_3_vc_sel_1_3 <= _GEN_215;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_0_1 <= io_vcalloc_resp_vc_sel_0_1; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_0_1 <= _GEN_217;
      end
    end else begin
      states_3_vc_sel_0_1 <= _GEN_217;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_0_2 <= io_vcalloc_resp_vc_sel_0_2; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_0_2 <= _GEN_218;
      end
    end else begin
      states_3_vc_sel_0_2 <= _GEN_218;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_0_3 <= io_vcalloc_resp_vc_sel_0_3; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_0_3 <= _GEN_219;
      end
    end else begin
      states_3_vc_sel_0_3 <= _GEN_219;
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h3 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_3_flow_ingress_node <= io_in_flit_0_bits_flow_ingress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h3 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_3_flow_egress_node <= io_in_flit_0_bits_flow_egress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (reset) begin // @[InputUnit.scala 233:21]
      mask <= 4'h0; // @[InputUnit.scala 233:21]
    end else if (io_router_req_valid) begin // @[InputUnit.scala 239:31]
      mask <= _mask_T_2; // @[InputUnit.scala 240:10]
    end else if (_T_26) begin // @[InputUnit.scala 241:34]
      mask <= _mask_T_17; // @[InputUnit.scala 242:10]
    end
    salloc_outs_0_valid <= salloc_arb_io_out_0_ready & salloc_arb_io_out_0_valid; // @[Decoupled.scala 51:35]
    salloc_outs_0_out_vid <= _virt_channel_T_10 | _virt_channel_T_11; // @[Mux.scala 27:73]
    salloc_outs_0_flit_head <= salloc_arb_io_chosen_oh_0[0] & input_buffer_io_deq_0_bits_head |
      salloc_arb_io_chosen_oh_0[1] & input_buffer_io_deq_1_bits_head | salloc_arb_io_chosen_oh_0[2] &
      input_buffer_io_deq_2_bits_head | salloc_arb_io_chosen_oh_0[3] & input_buffer_io_deq_3_bits_head; // @[Mux.scala 27:73]
    salloc_outs_0_flit_tail <= salloc_arb_io_chosen_oh_0[0] & input_buffer_io_deq_0_bits_tail |
      salloc_arb_io_chosen_oh_0[1] & input_buffer_io_deq_1_bits_tail | salloc_arb_io_chosen_oh_0[2] &
      input_buffer_io_deq_2_bits_tail | salloc_arb_io_chosen_oh_0[3] & input_buffer_io_deq_3_bits_tail; // @[Mux.scala 27:73]
    salloc_outs_0_flit_payload <= _salloc_outs_0_flit_payload_T_9 | _salloc_outs_0_flit_payload_T_7; // @[Mux.scala 27:73]
    salloc_outs_0_flit_flow_ingress_node <= _salloc_outs_0_flit_flow_T_30 | _salloc_outs_0_flit_flow_T_28; // @[Mux.scala 27:73]
    salloc_outs_0_flit_flow_egress_node <= _salloc_outs_0_flit_flow_T_16 | _salloc_outs_0_flit_flow_T_14; // @[Mux.scala 27:73]
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T & _T_3 & ~(_GEN_3 == 3'h0)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:197 assert(states(id).g === g_i)\n"); // @[InputUnit.scala 197:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_router_req_valid & _T_3 & ~(_GEN_139 == 3'h1)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:224 assert(states(id).g === g_r)\n"); // @[InputUnit.scala 224:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_39 & vcalloc_sel[0] & _T_3 & ~vcalloc_vals_0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:274 assert(states(i).g === g_v)\n"); // @[InputUnit.scala 274:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_39 & vcalloc_sel[1] & _T_3 & ~vcalloc_vals_1) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:274 assert(states(i).g === g_v)\n"); // @[InputUnit.scala 274:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_39 & vcalloc_sel[2] & _T_3 & ~vcalloc_vals_2) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:274 assert(states(i).g === g_v)\n"); // @[InputUnit.scala 274:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_39 & vcalloc_sel[3] & _T_3 & ~vcalloc_vals_3) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:274 assert(states(i).g === g_v)\n"); // @[InputUnit.scala 274:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  states_0_g = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  states_0_vc_sel_2_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  states_0_vc_sel_1_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  states_0_vc_sel_0_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  states_0_flow_ingress_node = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  states_0_flow_egress_node = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  states_1_g = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  states_1_vc_sel_2_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  states_1_vc_sel_1_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  states_1_vc_sel_1_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  states_1_vc_sel_0_1 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  states_1_flow_ingress_node = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  states_1_flow_egress_node = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  states_2_g = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  states_2_vc_sel_2_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  states_2_vc_sel_1_0 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  states_2_vc_sel_1_1 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  states_2_vc_sel_1_2 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  states_2_vc_sel_0_1 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  states_2_vc_sel_0_2 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  states_2_flow_ingress_node = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  states_2_flow_egress_node = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  states_3_g = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  states_3_vc_sel_2_0 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  states_3_vc_sel_1_0 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  states_3_vc_sel_1_1 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  states_3_vc_sel_1_2 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  states_3_vc_sel_1_3 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  states_3_vc_sel_0_1 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  states_3_vc_sel_0_2 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  states_3_vc_sel_0_3 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  states_3_flow_ingress_node = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  states_3_flow_egress_node = _RAND_32[1:0];
  _RAND_33 = {1{`RANDOM}};
  mask = _RAND_33[3:0];
  _RAND_34 = {1{`RANDOM}};
  salloc_outs_0_valid = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  salloc_outs_0_out_vid = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  salloc_outs_0_flit_head = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  salloc_outs_0_flit_tail = _RAND_37[0:0];
  _RAND_38 = {2{`RANDOM}};
  salloc_outs_0_flit_payload = _RAND_38[63:0];
  _RAND_39 = {1{`RANDOM}};
  salloc_outs_0_flit_flow_ingress_node = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  salloc_outs_0_flit_flow_egress_node = _RAND_40[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (_T & ~reset) begin
      assert(1'h1); // @[InputUnit.scala 196:13]
    end
    //
    if (_T & _T_3) begin
      assert(_GEN_3 == 3'h0); // @[InputUnit.scala 197:13]
    end
    //
    if (io_router_req_valid & _T_3) begin
      assert(_GEN_139 == 3'h1); // @[InputUnit.scala 224:11]
    end
    //
    if (_T_39 & vcalloc_sel[0] & _T_3) begin
      assert(vcalloc_vals_0); // @[InputUnit.scala 274:17]
    end
    //
    if (_T_39 & vcalloc_sel[1] & _T_3) begin
      assert(vcalloc_vals_1); // @[InputUnit.scala 274:17]
    end
    //
    if (_T_39 & vcalloc_sel[2] & _T_3) begin
      assert(vcalloc_vals_2); // @[InputUnit.scala 274:17]
    end
    //
    if (_T_39 & vcalloc_sel[3] & _T_3) begin
      assert(vcalloc_vals_3); // @[InputUnit.scala 274:17]
    end
  end
endmodule
module InputUnit_3(
  input         clock,
  input         reset,
  output        io_router_req_valid,
  output [1:0]  io_router_req_bits_src_virt_id,
  output [1:0]  io_router_req_bits_flow_ingress_node,
  output [1:0]  io_router_req_bits_flow_egress_node,
  input         io_router_resp_vc_sel_1_0,
  input         io_router_resp_vc_sel_1_1,
  input         io_router_resp_vc_sel_1_2,
  input         io_router_resp_vc_sel_1_3,
  input         io_router_resp_vc_sel_0_0,
  input         io_router_resp_vc_sel_0_1,
  input         io_router_resp_vc_sel_0_2,
  input         io_router_resp_vc_sel_0_3,
  input         io_vcalloc_req_ready,
  output        io_vcalloc_req_valid,
  output        io_vcalloc_req_bits_vc_sel_2_0,
  output        io_vcalloc_req_bits_vc_sel_1_0,
  output        io_vcalloc_req_bits_vc_sel_1_1,
  output        io_vcalloc_req_bits_vc_sel_1_2,
  output        io_vcalloc_req_bits_vc_sel_1_3,
  output        io_vcalloc_req_bits_vc_sel_0_0,
  output        io_vcalloc_req_bits_vc_sel_0_1,
  output        io_vcalloc_req_bits_vc_sel_0_2,
  output        io_vcalloc_req_bits_vc_sel_0_3,
  input         io_vcalloc_resp_vc_sel_2_0,
  input         io_vcalloc_resp_vc_sel_1_0,
  input         io_vcalloc_resp_vc_sel_1_1,
  input         io_vcalloc_resp_vc_sel_1_2,
  input         io_vcalloc_resp_vc_sel_1_3,
  input         io_vcalloc_resp_vc_sel_0_0,
  input         io_vcalloc_resp_vc_sel_0_1,
  input         io_vcalloc_resp_vc_sel_0_2,
  input         io_vcalloc_resp_vc_sel_0_3,
  input         io_out_credit_available_2_0,
  input         io_out_credit_available_1_0,
  input         io_out_credit_available_1_1,
  input         io_out_credit_available_1_2,
  input         io_out_credit_available_1_3,
  input         io_out_credit_available_0_0,
  input         io_out_credit_available_0_1,
  input         io_out_credit_available_0_2,
  input         io_out_credit_available_0_3,
  input         io_salloc_req_0_ready,
  output        io_salloc_req_0_valid,
  output        io_salloc_req_0_bits_vc_sel_2_0,
  output        io_salloc_req_0_bits_vc_sel_1_0,
  output        io_salloc_req_0_bits_vc_sel_1_1,
  output        io_salloc_req_0_bits_vc_sel_1_2,
  output        io_salloc_req_0_bits_vc_sel_1_3,
  output        io_salloc_req_0_bits_vc_sel_0_0,
  output        io_salloc_req_0_bits_vc_sel_0_1,
  output        io_salloc_req_0_bits_vc_sel_0_2,
  output        io_salloc_req_0_bits_vc_sel_0_3,
  output        io_salloc_req_0_bits_tail,
  output        io_out_0_valid,
  output        io_out_0_bits_flit_head,
  output        io_out_0_bits_flit_tail,
  output [63:0] io_out_0_bits_flit_payload,
  output [1:0]  io_out_0_bits_flit_flow_ingress_node,
  output [1:0]  io_out_0_bits_flit_flow_egress_node,
  output [1:0]  io_out_0_bits_out_virt_channel,
  output [1:0]  io_debug_va_stall,
  output [1:0]  io_debug_sa_stall,
  input         io_in_flit_0_valid,
  input         io_in_flit_0_bits_head,
  input         io_in_flit_0_bits_tail,
  input  [63:0] io_in_flit_0_bits_payload,
  input  [1:0]  io_in_flit_0_bits_flow_ingress_node,
  input  [1:0]  io_in_flit_0_bits_flow_egress_node,
  input  [1:0]  io_in_flit_0_bits_virt_channel_id,
  output [3:0]  io_in_credit_return,
  output [3:0]  io_in_vc_free
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
`endif // RANDOMIZE_REG_INIT
  wire  input_buffer_clock; // @[InputUnit.scala 180:28]
  wire  input_buffer_reset; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_enq_0_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_enq_0_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_enq_0_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_enq_0_bits_payload; // @[InputUnit.scala 180:28]
  wire [1:0] input_buffer_io_enq_0_bits_virt_channel_id; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_0_ready; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_0_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_0_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_0_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_deq_0_bits_payload; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_ready; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_deq_1_bits_payload; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_ready; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_deq_2_bits_payload; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_3_ready; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_3_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_3_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_3_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_deq_3_bits_payload; // @[InputUnit.scala 180:28]
  wire  route_arbiter_io_in_0_valid; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_0_bits_flow_ingress_node; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_0_bits_flow_egress_node; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_1_ready; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_1_valid; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_1_bits_flow_ingress_node; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_1_bits_flow_egress_node; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_2_ready; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_2_valid; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_2_bits_flow_ingress_node; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_2_bits_flow_egress_node; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_3_ready; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_3_valid; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_3_bits_flow_ingress_node; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_3_bits_flow_egress_node; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_out_valid; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_out_bits_src_virt_id; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_out_bits_flow_ingress_node; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_out_bits_flow_egress_node; // @[InputUnit.scala 186:29]
  wire  salloc_arb_clock; // @[InputUnit.scala 279:26]
  wire  salloc_arb_reset; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_bits_vc_sel_2_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_bits_vc_sel_1_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_bits_tail; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_vc_sel_2_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_vc_sel_1_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_vc_sel_1_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_vc_sel_0_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_tail; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_2_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_1_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_1_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_1_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_0_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_0_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_tail; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_2_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_1_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_1_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_1_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_1_3; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_0_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_0_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_0_3; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_tail; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_2_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_1_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_1_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_1_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_1_3; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_0_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_0_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_0_3; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_tail; // @[InputUnit.scala 279:26]
  wire [3:0] salloc_arb_io_chosen_oh_0; // @[InputUnit.scala 279:26]
  reg [2:0] states_0_g; // @[InputUnit.scala 191:19]
  reg  states_0_vc_sel_2_0; // @[InputUnit.scala 191:19]
  reg  states_0_vc_sel_1_0; // @[InputUnit.scala 191:19]
  reg  states_0_vc_sel_0_0; // @[InputUnit.scala 191:19]
  reg [1:0] states_0_flow_ingress_node; // @[InputUnit.scala 191:19]
  reg [1:0] states_0_flow_egress_node; // @[InputUnit.scala 191:19]
  reg [2:0] states_1_g; // @[InputUnit.scala 191:19]
  reg  states_1_vc_sel_2_0; // @[InputUnit.scala 191:19]
  reg  states_1_vc_sel_1_1; // @[InputUnit.scala 191:19]
  reg  states_1_vc_sel_0_0; // @[InputUnit.scala 191:19]
  reg  states_1_vc_sel_0_1; // @[InputUnit.scala 191:19]
  reg [1:0] states_1_flow_ingress_node; // @[InputUnit.scala 191:19]
  reg [1:0] states_1_flow_egress_node; // @[InputUnit.scala 191:19]
  reg [2:0] states_2_g; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_2_0; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_1_1; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_1_2; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_0_0; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_0_1; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_0_2; // @[InputUnit.scala 191:19]
  reg [1:0] states_2_flow_ingress_node; // @[InputUnit.scala 191:19]
  reg [1:0] states_2_flow_egress_node; // @[InputUnit.scala 191:19]
  reg [2:0] states_3_g; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_2_0; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_1_1; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_1_2; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_1_3; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_0_0; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_0_1; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_0_2; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_0_3; // @[InputUnit.scala 191:19]
  reg [1:0] states_3_flow_ingress_node; // @[InputUnit.scala 191:19]
  reg [1:0] states_3_flow_egress_node; // @[InputUnit.scala 191:19]
  wire  _T = io_in_flit_0_valid & io_in_flit_0_bits_head; // @[InputUnit.scala 194:32]
  wire  _T_3 = ~reset; // @[InputUnit.scala 196:13]
  wire [2:0] _GEN_1 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? states_1_g : states_0_g; // @[InputUnit.scala 197:{27,27}]
  wire [2:0] _GEN_2 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? states_2_g : _GEN_1; // @[InputUnit.scala 197:{27,27}]
  wire [2:0] _GEN_3 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? states_3_g : _GEN_2; // @[InputUnit.scala 197:{27,27}]
  wire  at_dest = io_in_flit_0_bits_flow_egress_node == 2'h1; // @[InputUnit.scala 198:57]
  wire [2:0] _states_g_T = at_dest ? 3'h2 : 3'h1; // @[InputUnit.scala 199:26]
  wire [2:0] _GEN_4 = 2'h0 == io_in_flit_0_bits_virt_channel_id ? _states_g_T : states_0_g; // @[InputUnit.scala 191:19 199:{20,20}]
  wire [2:0] _GEN_5 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? _states_g_T : states_1_g; // @[InputUnit.scala 191:19 199:{20,20}]
  wire [2:0] _GEN_6 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? _states_g_T : states_2_g; // @[InputUnit.scala 191:19 199:{20,20}]
  wire [2:0] _GEN_7 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? _states_g_T : states_3_g; // @[InputUnit.scala 191:19 199:{20,20}]
  wire  _GEN_8 = 2'h0 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_0_vc_sel_0_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_9 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_1_vc_sel_0_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_10 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_0_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_11 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_0_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_13 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_1_vc_sel_0_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_14 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_0_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_15 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_0_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_18 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_0_2; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_19 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_0_2; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_23 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_0_3; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_24 = 2'h0 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_0_vc_sel_1_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_29 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_1_vc_sel_1_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_30 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_1_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_31 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_1_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_34 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_1_2; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_35 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_1_2; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_39 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_1_3; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_40 = 2'h0 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_0_vc_sel_2_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_41 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_1_vc_sel_2_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_42 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_2_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_43 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_2_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_44 = 2'h0 == io_in_flit_0_bits_virt_channel_id | _GEN_40; // @[InputUnit.scala 203:{44,44}]
  wire  _GEN_45 = 2'h1 == io_in_flit_0_bits_virt_channel_id | _GEN_41; // @[InputUnit.scala 203:{44,44}]
  wire  _GEN_46 = 2'h2 == io_in_flit_0_bits_virt_channel_id | _GEN_42; // @[InputUnit.scala 203:{44,44}]
  wire  _GEN_47 = 2'h3 == io_in_flit_0_bits_virt_channel_id | _GEN_43; // @[InputUnit.scala 203:{44,44}]
  wire [2:0] _GEN_72 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_4 : states_0_g; // @[InputUnit.scala 191:19 194:60]
  wire [2:0] _GEN_73 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_5 : states_1_g; // @[InputUnit.scala 191:19 194:60]
  wire [2:0] _GEN_74 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_6 : states_2_g; // @[InputUnit.scala 191:19 194:60]
  wire [2:0] _GEN_75 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_7 : states_3_g; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_76 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_8 : states_0_vc_sel_0_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_77 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_9 : states_1_vc_sel_0_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_78 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_10 : states_2_vc_sel_0_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_79 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_11 : states_3_vc_sel_0_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_81 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_13 : states_1_vc_sel_0_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_82 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_14 : states_2_vc_sel_0_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_83 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_15 : states_3_vc_sel_0_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_86 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_18 : states_2_vc_sel_0_2; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_87 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_19 : states_3_vc_sel_0_2; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_91 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_23 : states_3_vc_sel_0_3; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_92 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_24 : states_0_vc_sel_1_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_97 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_29 : states_1_vc_sel_1_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_98 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_30 : states_2_vc_sel_1_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_99 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_31 : states_3_vc_sel_1_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_102 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_34 : states_2_vc_sel_1_2; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_103 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_35 : states_3_vc_sel_1_2; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_107 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_39 : states_3_vc_sel_1_3; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_108 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_44 : states_0_vc_sel_2_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_109 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_45 : states_1_vc_sel_2_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_110 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_46 : states_2_vc_sel_2_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_111 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_47 : states_3_vc_sel_2_0; // @[InputUnit.scala 191:19 194:60]
  wire  _T_10 = route_arbiter_io_in_0_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_132 = _T_10 ? 3'h2 : _GEN_72; // @[InputUnit.scala 215:{23,29}]
  wire  _T_11 = route_arbiter_io_in_1_ready & route_arbiter_io_in_1_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_133 = _T_11 ? 3'h2 : _GEN_73; // @[InputUnit.scala 215:{23,29}]
  wire  _T_12 = route_arbiter_io_in_2_ready & route_arbiter_io_in_2_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_134 = _T_12 ? 3'h2 : _GEN_74; // @[InputUnit.scala 215:{23,29}]
  wire  _T_13 = route_arbiter_io_in_3_ready & route_arbiter_io_in_3_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_135 = _T_13 ? 3'h2 : _GEN_75; // @[InputUnit.scala 215:{23,29}]
  wire [2:0] _GEN_137 = 2'h1 == io_router_req_bits_src_virt_id ? states_1_g : states_0_g; // @[InputUnit.scala 224:{25,25}]
  wire [2:0] _GEN_138 = 2'h2 == io_router_req_bits_src_virt_id ? states_2_g : _GEN_137; // @[InputUnit.scala 224:{25,25}]
  wire [2:0] _GEN_139 = 2'h3 == io_router_req_bits_src_virt_id ? states_3_g : _GEN_138; // @[InputUnit.scala 224:{25,25}]
  wire [2:0] _GEN_140 = 2'h0 == io_router_req_bits_src_virt_id ? 3'h2 : _GEN_132; // @[InputUnit.scala 225:{18,18}]
  wire [2:0] _GEN_141 = 2'h1 == io_router_req_bits_src_virt_id ? 3'h2 : _GEN_133; // @[InputUnit.scala 225:{18,18}]
  wire [2:0] _GEN_142 = 2'h2 == io_router_req_bits_src_virt_id ? 3'h2 : _GEN_134; // @[InputUnit.scala 225:{18,18}]
  wire [2:0] _GEN_143 = 2'h3 == io_router_req_bits_src_virt_id ? 3'h2 : _GEN_135; // @[InputUnit.scala 225:{18,18}]
  wire  _GEN_144 = 2'h0 == io_router_req_bits_src_virt_id ? 1'h0 : _GEN_108; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_145 = 2'h0 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_0 : _GEN_92; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_149 = 2'h0 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_0 : _GEN_76; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_153 = 2'h1 == io_router_req_bits_src_virt_id ? 1'h0 : _GEN_109; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_155 = 2'h1 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_1 : _GEN_97; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_158 = 2'h1 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_0 : _GEN_77; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_159 = 2'h1 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_1 : _GEN_81; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_162 = 2'h2 == io_router_req_bits_src_virt_id ? 1'h0 : _GEN_110; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_164 = 2'h2 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_1 : _GEN_98; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_165 = 2'h2 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_2 : _GEN_102; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_167 = 2'h2 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_0 : _GEN_78; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_168 = 2'h2 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_1 : _GEN_82; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_169 = 2'h2 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_2 : _GEN_86; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_171 = 2'h3 == io_router_req_bits_src_virt_id ? 1'h0 : _GEN_111; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_173 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_1 : _GEN_99; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_174 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_2 : _GEN_103; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_175 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_3 : _GEN_107; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_176 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_0 : _GEN_79; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_177 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_1 : _GEN_83; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_178 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_2 : _GEN_87; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_179 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_3 : _GEN_91; // @[InputUnit.scala 227:25 228:26]
  wire [2:0] _GEN_180 = io_router_req_valid ? _GEN_140 : _GEN_132; // @[InputUnit.scala 222:31]
  wire [2:0] _GEN_181 = io_router_req_valid ? _GEN_141 : _GEN_133; // @[InputUnit.scala 222:31]
  wire [2:0] _GEN_182 = io_router_req_valid ? _GEN_142 : _GEN_134; // @[InputUnit.scala 222:31]
  wire [2:0] _GEN_183 = io_router_req_valid ? _GEN_143 : _GEN_135; // @[InputUnit.scala 222:31]
  wire  _GEN_184 = io_router_req_valid ? _GEN_144 : _GEN_108; // @[InputUnit.scala 222:31]
  wire  _GEN_185 = io_router_req_valid ? _GEN_145 : _GEN_92; // @[InputUnit.scala 222:31]
  wire  _GEN_189 = io_router_req_valid ? _GEN_149 : _GEN_76; // @[InputUnit.scala 222:31]
  wire  _GEN_193 = io_router_req_valid ? _GEN_153 : _GEN_109; // @[InputUnit.scala 222:31]
  wire  _GEN_195 = io_router_req_valid ? _GEN_155 : _GEN_97; // @[InputUnit.scala 222:31]
  wire  _GEN_198 = io_router_req_valid ? _GEN_158 : _GEN_77; // @[InputUnit.scala 222:31]
  wire  _GEN_199 = io_router_req_valid ? _GEN_159 : _GEN_81; // @[InputUnit.scala 222:31]
  wire  _GEN_202 = io_router_req_valid ? _GEN_162 : _GEN_110; // @[InputUnit.scala 222:31]
  wire  _GEN_204 = io_router_req_valid ? _GEN_164 : _GEN_98; // @[InputUnit.scala 222:31]
  wire  _GEN_205 = io_router_req_valid ? _GEN_165 : _GEN_102; // @[InputUnit.scala 222:31]
  wire  _GEN_207 = io_router_req_valid ? _GEN_167 : _GEN_78; // @[InputUnit.scala 222:31]
  wire  _GEN_208 = io_router_req_valid ? _GEN_168 : _GEN_82; // @[InputUnit.scala 222:31]
  wire  _GEN_209 = io_router_req_valid ? _GEN_169 : _GEN_86; // @[InputUnit.scala 222:31]
  wire  _GEN_211 = io_router_req_valid ? _GEN_171 : _GEN_111; // @[InputUnit.scala 222:31]
  wire  _GEN_213 = io_router_req_valid ? _GEN_173 : _GEN_99; // @[InputUnit.scala 222:31]
  wire  _GEN_214 = io_router_req_valid ? _GEN_174 : _GEN_103; // @[InputUnit.scala 222:31]
  wire  _GEN_215 = io_router_req_valid ? _GEN_175 : _GEN_107; // @[InputUnit.scala 222:31]
  wire  _GEN_216 = io_router_req_valid ? _GEN_176 : _GEN_79; // @[InputUnit.scala 222:31]
  wire  _GEN_217 = io_router_req_valid ? _GEN_177 : _GEN_83; // @[InputUnit.scala 222:31]
  wire  _GEN_218 = io_router_req_valid ? _GEN_178 : _GEN_87; // @[InputUnit.scala 222:31]
  wire  _GEN_219 = io_router_req_valid ? _GEN_179 : _GEN_91; // @[InputUnit.scala 222:31]
  reg [3:0] mask; // @[InputUnit.scala 233:21]
  wire  vcalloc_vals_1 = states_1_g == 3'h2; // @[InputUnit.scala 249:32]
  wire  vcalloc_vals_0 = states_0_g == 3'h2; // @[InputUnit.scala 249:32]
  wire  vcalloc_vals_3 = states_3_g == 3'h2; // @[InputUnit.scala 249:32]
  wire  vcalloc_vals_2 = states_2_g == 3'h2; // @[InputUnit.scala 249:32]
  wire [3:0] _vcalloc_filter_T = {vcalloc_vals_3,vcalloc_vals_2,vcalloc_vals_1,vcalloc_vals_0}; // @[InputUnit.scala 236:59]
  wire [3:0] _vcalloc_filter_T_2 = ~mask; // @[InputUnit.scala 236:89]
  wire [3:0] _vcalloc_filter_T_3 = _vcalloc_filter_T & _vcalloc_filter_T_2; // @[InputUnit.scala 236:87]
  wire [7:0] _vcalloc_filter_T_4 = {vcalloc_vals_3,vcalloc_vals_2,vcalloc_vals_1,vcalloc_vals_0,_vcalloc_filter_T_3}; // @[Cat.scala 33:92]
  wire [7:0] _vcalloc_filter_T_13 = _vcalloc_filter_T_4[7] ? 8'h80 : 8'h0; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_14 = _vcalloc_filter_T_4[6] ? 8'h40 : _vcalloc_filter_T_13; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_15 = _vcalloc_filter_T_4[5] ? 8'h20 : _vcalloc_filter_T_14; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_16 = _vcalloc_filter_T_4[4] ? 8'h10 : _vcalloc_filter_T_15; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_17 = _vcalloc_filter_T_4[3] ? 8'h8 : _vcalloc_filter_T_16; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_18 = _vcalloc_filter_T_4[2] ? 8'h4 : _vcalloc_filter_T_17; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_19 = _vcalloc_filter_T_4[1] ? 8'h2 : _vcalloc_filter_T_18; // @[Mux.scala 47:70]
  wire [7:0] vcalloc_filter = _vcalloc_filter_T_4[0] ? 8'h1 : _vcalloc_filter_T_19; // @[Mux.scala 47:70]
  wire [3:0] vcalloc_sel = vcalloc_filter[3:0] | vcalloc_filter[7:4]; // @[InputUnit.scala 237:58]
  wire [3:0] _mask_T = 4'h1 << io_router_req_bits_src_virt_id; // @[InputUnit.scala 240:18]
  wire [3:0] _mask_T_2 = _mask_T - 4'h1; // @[InputUnit.scala 240:53]
  wire  _T_26 = vcalloc_vals_0 | vcalloc_vals_1 | vcalloc_vals_2 | vcalloc_vals_3; // @[package.scala 73:59]
  wire [1:0] _mask_T_12 = vcalloc_sel[1] ? 2'h3 : 2'h0; // @[Mux.scala 27:73]
  wire [2:0] _mask_T_13 = vcalloc_sel[2] ? 3'h7 : 3'h0; // @[Mux.scala 27:73]
  wire [3:0] _mask_T_14 = vcalloc_sel[3] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [1:0] _GEN_60 = {{1'd0}, vcalloc_sel[0]}; // @[Mux.scala 27:73]
  wire [1:0] _mask_T_15 = _GEN_60 | _mask_T_12; // @[Mux.scala 27:73]
  wire [2:0] _GEN_61 = {{1'd0}, _mask_T_15}; // @[Mux.scala 27:73]
  wire [2:0] _mask_T_16 = _GEN_61 | _mask_T_13; // @[Mux.scala 27:73]
  wire [3:0] _GEN_62 = {{1'd0}, _mask_T_16}; // @[Mux.scala 27:73]
  wire [3:0] _mask_T_17 = _GEN_62 | _mask_T_14; // @[Mux.scala 27:73]
  wire [2:0] _GEN_222 = vcalloc_vals_0 & vcalloc_sel[0] & io_vcalloc_req_ready ? 3'h3 : _GEN_180; // @[InputUnit.scala 253:{76,82}]
  wire [2:0] _GEN_223 = vcalloc_vals_1 & vcalloc_sel[1] & io_vcalloc_req_ready ? 3'h3 : _GEN_181; // @[InputUnit.scala 253:{76,82}]
  wire [2:0] _GEN_224 = vcalloc_vals_2 & vcalloc_sel[2] & io_vcalloc_req_ready ? 3'h3 : _GEN_182; // @[InputUnit.scala 253:{76,82}]
  wire [2:0] _GEN_225 = vcalloc_vals_3 & vcalloc_sel[3] & io_vcalloc_req_ready ? 3'h3 : _GEN_183; // @[InputUnit.scala 253:{76,82}]
  wire [1:0] _io_debug_va_stall_T = vcalloc_vals_0 + vcalloc_vals_1; // @[Bitwise.scala 51:90]
  wire [1:0] _io_debug_va_stall_T_2 = vcalloc_vals_2 + vcalloc_vals_3; // @[Bitwise.scala 51:90]
  wire [2:0] _io_debug_va_stall_T_4 = _io_debug_va_stall_T + _io_debug_va_stall_T_2; // @[Bitwise.scala 51:90]
  wire [2:0] _GEN_63 = {{2'd0}, io_vcalloc_req_ready}; // @[InputUnit.scala 266:47]
  wire [2:0] _io_debug_va_stall_T_7 = _io_debug_va_stall_T_4 - _GEN_63; // @[InputUnit.scala 266:47]
  wire  _T_39 = io_vcalloc_req_ready & io_vcalloc_req_valid; // @[Decoupled.scala 51:35]
  wire [8:0] _credit_available_T = {states_0_vc_sel_2_0,1'h0,1'h0,1'h0,states_0_vc_sel_1_0,2'h0,1'h0,states_0_vc_sel_0_0
    }; // @[InputUnit.scala 287:40]
  wire [8:0] _credit_available_T_1 = {io_out_credit_available_2_0,io_out_credit_available_1_3,
    io_out_credit_available_1_2,io_out_credit_available_1_1,io_out_credit_available_1_0,io_out_credit_available_0_3,
    io_out_credit_available_0_2,io_out_credit_available_0_1,io_out_credit_available_0_0}; // @[InputUnit.scala 287:73]
  wire [8:0] _credit_available_T_2 = _credit_available_T & _credit_available_T_1; // @[InputUnit.scala 287:47]
  wire  credit_available = _credit_available_T_2 != 9'h0; // @[InputUnit.scala 287:81]
  wire  _T_60 = salloc_arb_io_in_0_ready & salloc_arb_io_in_0_valid; // @[Decoupled.scala 51:35]
  wire [8:0] _credit_available_T_3 = {states_1_vc_sel_2_0,1'h0,1'h0,states_1_vc_sel_1_1,1'h0,2'h0,states_1_vc_sel_0_1,
    states_1_vc_sel_0_0}; // @[InputUnit.scala 287:40]
  wire [8:0] _credit_available_T_5 = _credit_available_T_3 & _credit_available_T_1; // @[InputUnit.scala 287:47]
  wire  credit_available_1 = _credit_available_T_5 != 9'h0; // @[InputUnit.scala 287:81]
  wire  _T_62 = salloc_arb_io_in_1_ready & salloc_arb_io_in_1_valid; // @[Decoupled.scala 51:35]
  wire [8:0] _credit_available_T_6 = {states_2_vc_sel_2_0,1'h0,states_2_vc_sel_1_2,states_2_vc_sel_1_1,1'h0,1'h0,
    states_2_vc_sel_0_2,states_2_vc_sel_0_1,states_2_vc_sel_0_0}; // @[InputUnit.scala 287:40]
  wire [8:0] _credit_available_T_8 = _credit_available_T_6 & _credit_available_T_1; // @[InputUnit.scala 287:47]
  wire  credit_available_2 = _credit_available_T_8 != 9'h0; // @[InputUnit.scala 287:81]
  wire  _T_64 = salloc_arb_io_in_2_ready & salloc_arb_io_in_2_valid; // @[Decoupled.scala 51:35]
  wire [8:0] _credit_available_T_9 = {states_3_vc_sel_2_0,states_3_vc_sel_1_3,states_3_vc_sel_1_2,states_3_vc_sel_1_1,1'h0
    ,states_3_vc_sel_0_3,states_3_vc_sel_0_2,states_3_vc_sel_0_1,states_3_vc_sel_0_0}; // @[InputUnit.scala 287:40]
  wire [8:0] _credit_available_T_11 = _credit_available_T_9 & _credit_available_T_1; // @[InputUnit.scala 287:47]
  wire  credit_available_3 = _credit_available_T_11 != 9'h0; // @[InputUnit.scala 287:81]
  wire  _T_66 = salloc_arb_io_in_3_ready & salloc_arb_io_in_3_valid; // @[Decoupled.scala 51:35]
  wire  _io_debug_sa_stall_T_1 = salloc_arb_io_in_0_valid & ~salloc_arb_io_in_0_ready; // @[InputUnit.scala 301:67]
  wire  _io_debug_sa_stall_T_3 = salloc_arb_io_in_1_valid & ~salloc_arb_io_in_1_ready; // @[InputUnit.scala 301:67]
  wire  _io_debug_sa_stall_T_5 = salloc_arb_io_in_2_valid & ~salloc_arb_io_in_2_ready; // @[InputUnit.scala 301:67]
  wire  _io_debug_sa_stall_T_7 = salloc_arb_io_in_3_valid & ~salloc_arb_io_in_3_ready; // @[InputUnit.scala 301:67]
  wire [1:0] _io_debug_sa_stall_T_8 = _io_debug_sa_stall_T_1 + _io_debug_sa_stall_T_3; // @[Bitwise.scala 51:90]
  wire [1:0] _io_debug_sa_stall_T_10 = _io_debug_sa_stall_T_5 + _io_debug_sa_stall_T_7; // @[Bitwise.scala 51:90]
  wire [2:0] _io_debug_sa_stall_T_12 = _io_debug_sa_stall_T_8 + _io_debug_sa_stall_T_10; // @[Bitwise.scala 51:90]
  reg  salloc_outs_0_valid; // @[InputUnit.scala 318:8]
  reg [1:0] salloc_outs_0_out_vid; // @[InputUnit.scala 318:8]
  reg  salloc_outs_0_flit_head; // @[InputUnit.scala 318:8]
  reg  salloc_outs_0_flit_tail; // @[InputUnit.scala 318:8]
  reg [63:0] salloc_outs_0_flit_payload; // @[InputUnit.scala 318:8]
  reg [1:0] salloc_outs_0_flit_flow_ingress_node; // @[InputUnit.scala 318:8]
  reg [1:0] salloc_outs_0_flit_flow_egress_node; // @[InputUnit.scala 318:8]
  wire  _io_in_credit_return_T = salloc_arb_io_out_0_ready & salloc_arb_io_out_0_valid; // @[Decoupled.scala 51:35]
  wire  _io_in_vc_free_T_11 = salloc_arb_io_chosen_oh_0[0] & input_buffer_io_deq_0_bits_tail | salloc_arb_io_chosen_oh_0
    [1] & input_buffer_io_deq_1_bits_tail | salloc_arb_io_chosen_oh_0[2] & input_buffer_io_deq_2_bits_tail |
    salloc_arb_io_chosen_oh_0[3] & input_buffer_io_deq_3_bits_tail; // @[Mux.scala 27:73]
  wire  vc_sel_0_0 = salloc_arb_io_chosen_oh_0[0] & states_0_vc_sel_0_0 | salloc_arb_io_chosen_oh_0[1] &
    states_1_vc_sel_0_0 | salloc_arb_io_chosen_oh_0[2] & states_2_vc_sel_0_0 | salloc_arb_io_chosen_oh_0[3] &
    states_3_vc_sel_0_0; // @[Mux.scala 27:73]
  wire  vc_sel_0_1 = salloc_arb_io_chosen_oh_0[1] & states_1_vc_sel_0_1 | salloc_arb_io_chosen_oh_0[2] &
    states_2_vc_sel_0_1 | salloc_arb_io_chosen_oh_0[3] & states_3_vc_sel_0_1; // @[Mux.scala 27:73]
  wire  vc_sel_0_2 = salloc_arb_io_chosen_oh_0[2] & states_2_vc_sel_0_2 | salloc_arb_io_chosen_oh_0[3] &
    states_3_vc_sel_0_2; // @[Mux.scala 27:73]
  wire  vc_sel_0_3 = salloc_arb_io_chosen_oh_0[3] & states_3_vc_sel_0_3; // @[Mux.scala 27:73]
  wire  vc_sel_1_0 = salloc_arb_io_chosen_oh_0[0] & states_0_vc_sel_1_0; // @[Mux.scala 27:73]
  wire  vc_sel_1_1 = salloc_arb_io_chosen_oh_0[1] & states_1_vc_sel_1_1 | salloc_arb_io_chosen_oh_0[2] &
    states_2_vc_sel_1_1 | salloc_arb_io_chosen_oh_0[3] & states_3_vc_sel_1_1; // @[Mux.scala 27:73]
  wire  vc_sel_1_2 = salloc_arb_io_chosen_oh_0[2] & states_2_vc_sel_1_2 | salloc_arb_io_chosen_oh_0[3] &
    states_3_vc_sel_1_2; // @[Mux.scala 27:73]
  wire  vc_sel_1_3 = salloc_arb_io_chosen_oh_0[3] & states_3_vc_sel_1_3; // @[Mux.scala 27:73]
  wire  channel_oh_0 = vc_sel_0_0 | vc_sel_0_1 | vc_sel_0_2 | vc_sel_0_3; // @[InputUnit.scala 334:43]
  wire  channel_oh_1 = vc_sel_1_0 | vc_sel_1_1 | vc_sel_1_2 | vc_sel_1_3; // @[InputUnit.scala 334:43]
  wire [3:0] _virt_channel_T = {vc_sel_0_3,vc_sel_0_2,vc_sel_0_1,vc_sel_0_0}; // @[OneHot.scala 22:45]
  wire [1:0] virt_channel_hi_1 = _virt_channel_T[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] virt_channel_lo_1 = _virt_channel_T[1:0]; // @[OneHot.scala 31:18]
  wire  _virt_channel_T_1 = |virt_channel_hi_1; // @[OneHot.scala 32:14]
  wire [1:0] _virt_channel_T_2 = virt_channel_hi_1 | virt_channel_lo_1; // @[OneHot.scala 32:28]
  wire [1:0] _virt_channel_T_4 = {_virt_channel_T_1,_virt_channel_T_2[1]}; // @[Cat.scala 33:92]
  wire [3:0] _virt_channel_T_5 = {vc_sel_1_3,vc_sel_1_2,vc_sel_1_1,vc_sel_1_0}; // @[OneHot.scala 22:45]
  wire [1:0] virt_channel_hi_3 = _virt_channel_T_5[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] virt_channel_lo_3 = _virt_channel_T_5[1:0]; // @[OneHot.scala 31:18]
  wire  _virt_channel_T_6 = |virt_channel_hi_3; // @[OneHot.scala 32:14]
  wire [1:0] _virt_channel_T_7 = virt_channel_hi_3 | virt_channel_lo_3; // @[OneHot.scala 32:28]
  wire [1:0] _virt_channel_T_9 = {_virt_channel_T_6,_virt_channel_T_7[1]}; // @[Cat.scala 33:92]
  wire [1:0] _virt_channel_T_10 = channel_oh_0 ? _virt_channel_T_4 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _virt_channel_T_11 = channel_oh_1 ? _virt_channel_T_9 : 2'h0; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_4 = salloc_arb_io_chosen_oh_0[0] ? input_buffer_io_deq_0_bits_payload : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_5 = salloc_arb_io_chosen_oh_0[1] ? input_buffer_io_deq_1_bits_payload : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_6 = salloc_arb_io_chosen_oh_0[2] ? input_buffer_io_deq_2_bits_payload : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_7 = salloc_arb_io_chosen_oh_0[3] ? input_buffer_io_deq_3_bits_payload : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_8 = _salloc_outs_0_flit_payload_T_4 | _salloc_outs_0_flit_payload_T_5; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_9 = _salloc_outs_0_flit_payload_T_8 | _salloc_outs_0_flit_payload_T_6; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_11 = salloc_arb_io_chosen_oh_0[0] ? states_0_flow_egress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_12 = salloc_arb_io_chosen_oh_0[1] ? states_1_flow_egress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_13 = salloc_arb_io_chosen_oh_0[2] ? states_2_flow_egress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_14 = salloc_arb_io_chosen_oh_0[3] ? states_3_flow_egress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_15 = _salloc_outs_0_flit_flow_T_11 | _salloc_outs_0_flit_flow_T_12; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_16 = _salloc_outs_0_flit_flow_T_15 | _salloc_outs_0_flit_flow_T_13; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_25 = salloc_arb_io_chosen_oh_0[0] ? states_0_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_26 = salloc_arb_io_chosen_oh_0[1] ? states_1_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_27 = salloc_arb_io_chosen_oh_0[2] ? states_2_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_28 = salloc_arb_io_chosen_oh_0[3] ? states_3_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_29 = _salloc_outs_0_flit_flow_T_25 | _salloc_outs_0_flit_flow_T_26; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_30 = _salloc_outs_0_flit_flow_T_29 | _salloc_outs_0_flit_flow_T_27; // @[Mux.scala 27:73]
  InputBuffer input_buffer ( // @[InputUnit.scala 180:28]
    .clock(input_buffer_clock),
    .reset(input_buffer_reset),
    .io_enq_0_valid(input_buffer_io_enq_0_valid),
    .io_enq_0_bits_head(input_buffer_io_enq_0_bits_head),
    .io_enq_0_bits_tail(input_buffer_io_enq_0_bits_tail),
    .io_enq_0_bits_payload(input_buffer_io_enq_0_bits_payload),
    .io_enq_0_bits_virt_channel_id(input_buffer_io_enq_0_bits_virt_channel_id),
    .io_deq_0_ready(input_buffer_io_deq_0_ready),
    .io_deq_0_valid(input_buffer_io_deq_0_valid),
    .io_deq_0_bits_head(input_buffer_io_deq_0_bits_head),
    .io_deq_0_bits_tail(input_buffer_io_deq_0_bits_tail),
    .io_deq_0_bits_payload(input_buffer_io_deq_0_bits_payload),
    .io_deq_1_ready(input_buffer_io_deq_1_ready),
    .io_deq_1_valid(input_buffer_io_deq_1_valid),
    .io_deq_1_bits_head(input_buffer_io_deq_1_bits_head),
    .io_deq_1_bits_tail(input_buffer_io_deq_1_bits_tail),
    .io_deq_1_bits_payload(input_buffer_io_deq_1_bits_payload),
    .io_deq_2_ready(input_buffer_io_deq_2_ready),
    .io_deq_2_valid(input_buffer_io_deq_2_valid),
    .io_deq_2_bits_head(input_buffer_io_deq_2_bits_head),
    .io_deq_2_bits_tail(input_buffer_io_deq_2_bits_tail),
    .io_deq_2_bits_payload(input_buffer_io_deq_2_bits_payload),
    .io_deq_3_ready(input_buffer_io_deq_3_ready),
    .io_deq_3_valid(input_buffer_io_deq_3_valid),
    .io_deq_3_bits_head(input_buffer_io_deq_3_bits_head),
    .io_deq_3_bits_tail(input_buffer_io_deq_3_bits_tail),
    .io_deq_3_bits_payload(input_buffer_io_deq_3_bits_payload)
  );
  Arbiter route_arbiter ( // @[InputUnit.scala 186:29]
    .io_in_0_valid(route_arbiter_io_in_0_valid),
    .io_in_0_bits_flow_ingress_node(route_arbiter_io_in_0_bits_flow_ingress_node),
    .io_in_0_bits_flow_egress_node(route_arbiter_io_in_0_bits_flow_egress_node),
    .io_in_1_ready(route_arbiter_io_in_1_ready),
    .io_in_1_valid(route_arbiter_io_in_1_valid),
    .io_in_1_bits_flow_ingress_node(route_arbiter_io_in_1_bits_flow_ingress_node),
    .io_in_1_bits_flow_egress_node(route_arbiter_io_in_1_bits_flow_egress_node),
    .io_in_2_ready(route_arbiter_io_in_2_ready),
    .io_in_2_valid(route_arbiter_io_in_2_valid),
    .io_in_2_bits_flow_ingress_node(route_arbiter_io_in_2_bits_flow_ingress_node),
    .io_in_2_bits_flow_egress_node(route_arbiter_io_in_2_bits_flow_egress_node),
    .io_in_3_ready(route_arbiter_io_in_3_ready),
    .io_in_3_valid(route_arbiter_io_in_3_valid),
    .io_in_3_bits_flow_ingress_node(route_arbiter_io_in_3_bits_flow_ingress_node),
    .io_in_3_bits_flow_egress_node(route_arbiter_io_in_3_bits_flow_egress_node),
    .io_out_valid(route_arbiter_io_out_valid),
    .io_out_bits_src_virt_id(route_arbiter_io_out_bits_src_virt_id),
    .io_out_bits_flow_ingress_node(route_arbiter_io_out_bits_flow_ingress_node),
    .io_out_bits_flow_egress_node(route_arbiter_io_out_bits_flow_egress_node)
  );
  SwitchArbiter salloc_arb ( // @[InputUnit.scala 279:26]
    .clock(salloc_arb_clock),
    .reset(salloc_arb_reset),
    .io_in_0_ready(salloc_arb_io_in_0_ready),
    .io_in_0_valid(salloc_arb_io_in_0_valid),
    .io_in_0_bits_vc_sel_2_0(salloc_arb_io_in_0_bits_vc_sel_2_0),
    .io_in_0_bits_vc_sel_1_0(salloc_arb_io_in_0_bits_vc_sel_1_0),
    .io_in_0_bits_vc_sel_0_0(salloc_arb_io_in_0_bits_vc_sel_0_0),
    .io_in_0_bits_tail(salloc_arb_io_in_0_bits_tail),
    .io_in_1_ready(salloc_arb_io_in_1_ready),
    .io_in_1_valid(salloc_arb_io_in_1_valid),
    .io_in_1_bits_vc_sel_2_0(salloc_arb_io_in_1_bits_vc_sel_2_0),
    .io_in_1_bits_vc_sel_1_0(salloc_arb_io_in_1_bits_vc_sel_1_0),
    .io_in_1_bits_vc_sel_1_1(salloc_arb_io_in_1_bits_vc_sel_1_1),
    .io_in_1_bits_vc_sel_0_0(salloc_arb_io_in_1_bits_vc_sel_0_0),
    .io_in_1_bits_vc_sel_0_1(salloc_arb_io_in_1_bits_vc_sel_0_1),
    .io_in_1_bits_tail(salloc_arb_io_in_1_bits_tail),
    .io_in_2_ready(salloc_arb_io_in_2_ready),
    .io_in_2_valid(salloc_arb_io_in_2_valid),
    .io_in_2_bits_vc_sel_2_0(salloc_arb_io_in_2_bits_vc_sel_2_0),
    .io_in_2_bits_vc_sel_1_0(salloc_arb_io_in_2_bits_vc_sel_1_0),
    .io_in_2_bits_vc_sel_1_1(salloc_arb_io_in_2_bits_vc_sel_1_1),
    .io_in_2_bits_vc_sel_1_2(salloc_arb_io_in_2_bits_vc_sel_1_2),
    .io_in_2_bits_vc_sel_0_0(salloc_arb_io_in_2_bits_vc_sel_0_0),
    .io_in_2_bits_vc_sel_0_1(salloc_arb_io_in_2_bits_vc_sel_0_1),
    .io_in_2_bits_vc_sel_0_2(salloc_arb_io_in_2_bits_vc_sel_0_2),
    .io_in_2_bits_tail(salloc_arb_io_in_2_bits_tail),
    .io_in_3_ready(salloc_arb_io_in_3_ready),
    .io_in_3_valid(salloc_arb_io_in_3_valid),
    .io_in_3_bits_vc_sel_2_0(salloc_arb_io_in_3_bits_vc_sel_2_0),
    .io_in_3_bits_vc_sel_1_0(salloc_arb_io_in_3_bits_vc_sel_1_0),
    .io_in_3_bits_vc_sel_1_1(salloc_arb_io_in_3_bits_vc_sel_1_1),
    .io_in_3_bits_vc_sel_1_2(salloc_arb_io_in_3_bits_vc_sel_1_2),
    .io_in_3_bits_vc_sel_1_3(salloc_arb_io_in_3_bits_vc_sel_1_3),
    .io_in_3_bits_vc_sel_0_0(salloc_arb_io_in_3_bits_vc_sel_0_0),
    .io_in_3_bits_vc_sel_0_1(salloc_arb_io_in_3_bits_vc_sel_0_1),
    .io_in_3_bits_vc_sel_0_2(salloc_arb_io_in_3_bits_vc_sel_0_2),
    .io_in_3_bits_vc_sel_0_3(salloc_arb_io_in_3_bits_vc_sel_0_3),
    .io_in_3_bits_tail(salloc_arb_io_in_3_bits_tail),
    .io_out_0_ready(salloc_arb_io_out_0_ready),
    .io_out_0_valid(salloc_arb_io_out_0_valid),
    .io_out_0_bits_vc_sel_2_0(salloc_arb_io_out_0_bits_vc_sel_2_0),
    .io_out_0_bits_vc_sel_1_0(salloc_arb_io_out_0_bits_vc_sel_1_0),
    .io_out_0_bits_vc_sel_1_1(salloc_arb_io_out_0_bits_vc_sel_1_1),
    .io_out_0_bits_vc_sel_1_2(salloc_arb_io_out_0_bits_vc_sel_1_2),
    .io_out_0_bits_vc_sel_1_3(salloc_arb_io_out_0_bits_vc_sel_1_3),
    .io_out_0_bits_vc_sel_0_0(salloc_arb_io_out_0_bits_vc_sel_0_0),
    .io_out_0_bits_vc_sel_0_1(salloc_arb_io_out_0_bits_vc_sel_0_1),
    .io_out_0_bits_vc_sel_0_2(salloc_arb_io_out_0_bits_vc_sel_0_2),
    .io_out_0_bits_vc_sel_0_3(salloc_arb_io_out_0_bits_vc_sel_0_3),
    .io_out_0_bits_tail(salloc_arb_io_out_0_bits_tail),
    .io_chosen_oh_0(salloc_arb_io_chosen_oh_0)
  );
  assign io_router_req_valid = route_arbiter_io_out_valid; // @[InputUnit.scala 189:17]
  assign io_router_req_bits_src_virt_id = route_arbiter_io_out_bits_src_virt_id; // @[InputUnit.scala 189:17]
  assign io_router_req_bits_flow_ingress_node = route_arbiter_io_out_bits_flow_ingress_node; // @[InputUnit.scala 189:17]
  assign io_router_req_bits_flow_egress_node = route_arbiter_io_out_bits_flow_egress_node; // @[InputUnit.scala 189:17]
  assign io_vcalloc_req_valid = vcalloc_vals_0 | vcalloc_vals_1 | vcalloc_vals_2 | vcalloc_vals_3; // @[package.scala 73:59]
  assign io_vcalloc_req_bits_vc_sel_2_0 = vcalloc_sel[0] & states_0_vc_sel_2_0 | vcalloc_sel[1] & states_1_vc_sel_2_0 |
    vcalloc_sel[2] & states_2_vc_sel_2_0 | vcalloc_sel[3] & states_3_vc_sel_2_0; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_1_0 = vcalloc_sel[0] & states_0_vc_sel_1_0; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_1_1 = vcalloc_sel[1] & states_1_vc_sel_1_1 | vcalloc_sel[2] & states_2_vc_sel_1_1 |
    vcalloc_sel[3] & states_3_vc_sel_1_1; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_1_2 = vcalloc_sel[2] & states_2_vc_sel_1_2 | vcalloc_sel[3] & states_3_vc_sel_1_2; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_1_3 = vcalloc_sel[3] & states_3_vc_sel_1_3; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_0_0 = vcalloc_sel[0] & states_0_vc_sel_0_0 | vcalloc_sel[1] & states_1_vc_sel_0_0 |
    vcalloc_sel[2] & states_2_vc_sel_0_0 | vcalloc_sel[3] & states_3_vc_sel_0_0; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_0_1 = vcalloc_sel[1] & states_1_vc_sel_0_1 | vcalloc_sel[2] & states_2_vc_sel_0_1 |
    vcalloc_sel[3] & states_3_vc_sel_0_1; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_0_2 = vcalloc_sel[2] & states_2_vc_sel_0_2 | vcalloc_sel[3] & states_3_vc_sel_0_2; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_0_3 = vcalloc_sel[3] & states_3_vc_sel_0_3; // @[Mux.scala 27:73]
  assign io_salloc_req_0_valid = salloc_arb_io_out_0_valid; // @[InputUnit.scala 302:17 303:19 305:35]
  assign io_salloc_req_0_bits_vc_sel_2_0 = salloc_arb_io_out_0_bits_vc_sel_2_0; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_1_0 = salloc_arb_io_out_0_bits_vc_sel_1_0; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_1_1 = salloc_arb_io_out_0_bits_vc_sel_1_1; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_1_2 = salloc_arb_io_out_0_bits_vc_sel_1_2; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_1_3 = salloc_arb_io_out_0_bits_vc_sel_1_3; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_0_0 = salloc_arb_io_out_0_bits_vc_sel_0_0; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_0_1 = salloc_arb_io_out_0_bits_vc_sel_0_1; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_0_2 = salloc_arb_io_out_0_bits_vc_sel_0_2; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_0_3 = salloc_arb_io_out_0_bits_vc_sel_0_3; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_tail = salloc_arb_io_out_0_bits_tail; // @[InputUnit.scala 302:17]
  assign io_out_0_valid = salloc_outs_0_valid; // @[InputUnit.scala 349:21]
  assign io_out_0_bits_flit_head = salloc_outs_0_flit_head; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_flit_tail = salloc_outs_0_flit_tail; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_flit_payload = salloc_outs_0_flit_payload; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_flit_flow_ingress_node = salloc_outs_0_flit_flow_ingress_node; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_flit_flow_egress_node = salloc_outs_0_flit_flow_egress_node; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_out_virt_channel = salloc_outs_0_out_vid; // @[InputUnit.scala 351:37]
  assign io_debug_va_stall = _io_debug_va_stall_T_7[1:0]; // @[InputUnit.scala 266:21]
  assign io_debug_sa_stall = _io_debug_sa_stall_T_12[1:0]; // @[InputUnit.scala 301:21]
  assign io_in_credit_return = _io_in_credit_return_T ? salloc_arb_io_chosen_oh_0 : 4'h0; // @[InputUnit.scala 322:8]
  assign io_in_vc_free = _io_in_credit_return_T & _io_in_vc_free_T_11 ? salloc_arb_io_chosen_oh_0 : 4'h0; // @[InputUnit.scala 325:8]
  assign input_buffer_clock = clock;
  assign input_buffer_reset = reset;
  assign input_buffer_io_enq_0_valid = io_in_flit_0_valid; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_head = io_in_flit_0_bits_head; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_tail = io_in_flit_0_bits_tail; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_payload = io_in_flit_0_bits_payload; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_virt_channel_id = io_in_flit_0_bits_virt_channel_id; // @[InputUnit.scala 182:28]
  assign input_buffer_io_deq_0_ready = salloc_arb_io_in_0_ready; // @[InputUnit.scala 295:36]
  assign input_buffer_io_deq_1_ready = salloc_arb_io_in_1_ready; // @[InputUnit.scala 295:36]
  assign input_buffer_io_deq_2_ready = salloc_arb_io_in_2_ready; // @[InputUnit.scala 295:36]
  assign input_buffer_io_deq_3_ready = salloc_arb_io_in_3_ready; // @[InputUnit.scala 295:36]
  assign route_arbiter_io_in_0_valid = states_0_g == 3'h1; // @[InputUnit.scala 212:22]
  assign route_arbiter_io_in_0_bits_flow_ingress_node = states_0_flow_ingress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_0_bits_flow_egress_node = states_0_flow_egress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_1_valid = states_1_g == 3'h1; // @[InputUnit.scala 212:22]
  assign route_arbiter_io_in_1_bits_flow_ingress_node = states_1_flow_ingress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_1_bits_flow_egress_node = states_1_flow_egress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_2_valid = states_2_g == 3'h1; // @[InputUnit.scala 212:22]
  assign route_arbiter_io_in_2_bits_flow_ingress_node = states_2_flow_ingress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_2_bits_flow_egress_node = states_2_flow_egress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_3_valid = states_3_g == 3'h1; // @[InputUnit.scala 212:22]
  assign route_arbiter_io_in_3_bits_flow_ingress_node = states_3_flow_ingress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_3_bits_flow_egress_node = states_3_flow_egress_node; // @[InputUnit.scala 213:19]
  assign salloc_arb_clock = clock;
  assign salloc_arb_reset = reset;
  assign salloc_arb_io_in_0_valid = states_0_g == 3'h3 & credit_available & input_buffer_io_deq_0_valid; // @[InputUnit.scala 288:50]
  assign salloc_arb_io_in_0_bits_vc_sel_2_0 = states_0_vc_sel_2_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_0_bits_vc_sel_1_0 = states_0_vc_sel_1_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_0_bits_vc_sel_0_0 = states_0_vc_sel_0_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_0_bits_tail = input_buffer_io_deq_0_bits_tail; // @[InputUnit.scala 291:19]
  assign salloc_arb_io_in_1_valid = states_1_g == 3'h3 & credit_available_1 & input_buffer_io_deq_1_valid; // @[InputUnit.scala 288:50]
  assign salloc_arb_io_in_1_bits_vc_sel_2_0 = states_1_vc_sel_2_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_1_bits_vc_sel_1_0 = 1'h0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_1_bits_vc_sel_1_1 = states_1_vc_sel_1_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_1_bits_vc_sel_0_0 = states_1_vc_sel_0_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_1_bits_vc_sel_0_1 = states_1_vc_sel_0_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_1_bits_tail = input_buffer_io_deq_1_bits_tail; // @[InputUnit.scala 291:19]
  assign salloc_arb_io_in_2_valid = states_2_g == 3'h3 & credit_available_2 & input_buffer_io_deq_2_valid; // @[InputUnit.scala 288:50]
  assign salloc_arb_io_in_2_bits_vc_sel_2_0 = states_2_vc_sel_2_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_1_0 = 1'h0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_1_1 = states_2_vc_sel_1_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_1_2 = states_2_vc_sel_1_2; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_0_0 = states_2_vc_sel_0_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_0_1 = states_2_vc_sel_0_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_0_2 = states_2_vc_sel_0_2; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_tail = input_buffer_io_deq_2_bits_tail; // @[InputUnit.scala 291:19]
  assign salloc_arb_io_in_3_valid = states_3_g == 3'h3 & credit_available_3 & input_buffer_io_deq_3_valid; // @[InputUnit.scala 288:50]
  assign salloc_arb_io_in_3_bits_vc_sel_2_0 = states_3_vc_sel_2_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_1_0 = 1'h0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_1_1 = states_3_vc_sel_1_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_1_2 = states_3_vc_sel_1_2; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_1_3 = states_3_vc_sel_1_3; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_0_0 = states_3_vc_sel_0_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_0_1 = states_3_vc_sel_0_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_0_2 = states_3_vc_sel_0_2; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_0_3 = states_3_vc_sel_0_3; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_tail = input_buffer_io_deq_3_bits_tail; // @[InputUnit.scala 291:19]
  assign salloc_arb_io_out_0_ready = io_salloc_req_0_ready; // @[InputUnit.scala 302:17 303:19 304:39]
  always @(posedge clock) begin
    if (reset) begin // @[InputUnit.scala 377:23]
      states_0_g <= 3'h0; // @[InputUnit.scala 378:24]
    end else if (_T_60 & input_buffer_io_deq_0_bits_tail) begin // @[InputUnit.scala 292:35]
      states_0_g <= 3'h0; // @[InputUnit.scala 293:13]
    end else if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[0]) begin // @[InputUnit.scala 270:29]
        states_0_g <= 3'h3; // @[InputUnit.scala 272:21]
      end else begin
        states_0_g <= _GEN_222;
      end
    end else begin
      states_0_g <= _GEN_222;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[0]) begin // @[InputUnit.scala 270:29]
        states_0_vc_sel_2_0 <= io_vcalloc_resp_vc_sel_2_0; // @[InputUnit.scala 271:26]
      end else begin
        states_0_vc_sel_2_0 <= _GEN_184;
      end
    end else begin
      states_0_vc_sel_2_0 <= _GEN_184;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[0]) begin // @[InputUnit.scala 270:29]
        states_0_vc_sel_1_0 <= io_vcalloc_resp_vc_sel_1_0; // @[InputUnit.scala 271:26]
      end else begin
        states_0_vc_sel_1_0 <= _GEN_185;
      end
    end else begin
      states_0_vc_sel_1_0 <= _GEN_185;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[0]) begin // @[InputUnit.scala 270:29]
        states_0_vc_sel_0_0 <= io_vcalloc_resp_vc_sel_0_0; // @[InputUnit.scala 271:26]
      end else begin
        states_0_vc_sel_0_0 <= _GEN_189;
      end
    end else begin
      states_0_vc_sel_0_0 <= _GEN_189;
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h0 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_0_flow_ingress_node <= io_in_flit_0_bits_flow_ingress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h0 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_0_flow_egress_node <= io_in_flit_0_bits_flow_egress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (reset) begin // @[InputUnit.scala 377:23]
      states_1_g <= 3'h0; // @[InputUnit.scala 378:24]
    end else if (_T_62 & input_buffer_io_deq_1_bits_tail) begin // @[InputUnit.scala 292:35]
      states_1_g <= 3'h0; // @[InputUnit.scala 293:13]
    end else if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_g <= 3'h3; // @[InputUnit.scala 272:21]
      end else begin
        states_1_g <= _GEN_223;
      end
    end else begin
      states_1_g <= _GEN_223;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_vc_sel_2_0 <= io_vcalloc_resp_vc_sel_2_0; // @[InputUnit.scala 271:26]
      end else begin
        states_1_vc_sel_2_0 <= _GEN_193;
      end
    end else begin
      states_1_vc_sel_2_0 <= _GEN_193;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_vc_sel_1_1 <= io_vcalloc_resp_vc_sel_1_1; // @[InputUnit.scala 271:26]
      end else begin
        states_1_vc_sel_1_1 <= _GEN_195;
      end
    end else begin
      states_1_vc_sel_1_1 <= _GEN_195;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_vc_sel_0_0 <= io_vcalloc_resp_vc_sel_0_0; // @[InputUnit.scala 271:26]
      end else begin
        states_1_vc_sel_0_0 <= _GEN_198;
      end
    end else begin
      states_1_vc_sel_0_0 <= _GEN_198;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_vc_sel_0_1 <= io_vcalloc_resp_vc_sel_0_1; // @[InputUnit.scala 271:26]
      end else begin
        states_1_vc_sel_0_1 <= _GEN_199;
      end
    end else begin
      states_1_vc_sel_0_1 <= _GEN_199;
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h1 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_1_flow_ingress_node <= io_in_flit_0_bits_flow_ingress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h1 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_1_flow_egress_node <= io_in_flit_0_bits_flow_egress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (reset) begin // @[InputUnit.scala 377:23]
      states_2_g <= 3'h0; // @[InputUnit.scala 378:24]
    end else if (_T_64 & input_buffer_io_deq_2_bits_tail) begin // @[InputUnit.scala 292:35]
      states_2_g <= 3'h0; // @[InputUnit.scala 293:13]
    end else if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_g <= 3'h3; // @[InputUnit.scala 272:21]
      end else begin
        states_2_g <= _GEN_224;
      end
    end else begin
      states_2_g <= _GEN_224;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_2_0 <= io_vcalloc_resp_vc_sel_2_0; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_2_0 <= _GEN_202;
      end
    end else begin
      states_2_vc_sel_2_0 <= _GEN_202;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_1_1 <= io_vcalloc_resp_vc_sel_1_1; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_1_1 <= _GEN_204;
      end
    end else begin
      states_2_vc_sel_1_1 <= _GEN_204;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_1_2 <= io_vcalloc_resp_vc_sel_1_2; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_1_2 <= _GEN_205;
      end
    end else begin
      states_2_vc_sel_1_2 <= _GEN_205;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_0_0 <= io_vcalloc_resp_vc_sel_0_0; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_0_0 <= _GEN_207;
      end
    end else begin
      states_2_vc_sel_0_0 <= _GEN_207;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_0_1 <= io_vcalloc_resp_vc_sel_0_1; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_0_1 <= _GEN_208;
      end
    end else begin
      states_2_vc_sel_0_1 <= _GEN_208;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_0_2 <= io_vcalloc_resp_vc_sel_0_2; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_0_2 <= _GEN_209;
      end
    end else begin
      states_2_vc_sel_0_2 <= _GEN_209;
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h2 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_2_flow_ingress_node <= io_in_flit_0_bits_flow_ingress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h2 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_2_flow_egress_node <= io_in_flit_0_bits_flow_egress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (reset) begin // @[InputUnit.scala 377:23]
      states_3_g <= 3'h0; // @[InputUnit.scala 378:24]
    end else if (_T_66 & input_buffer_io_deq_3_bits_tail) begin // @[InputUnit.scala 292:35]
      states_3_g <= 3'h0; // @[InputUnit.scala 293:13]
    end else if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_g <= 3'h3; // @[InputUnit.scala 272:21]
      end else begin
        states_3_g <= _GEN_225;
      end
    end else begin
      states_3_g <= _GEN_225;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_2_0 <= io_vcalloc_resp_vc_sel_2_0; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_2_0 <= _GEN_211;
      end
    end else begin
      states_3_vc_sel_2_0 <= _GEN_211;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_1_1 <= io_vcalloc_resp_vc_sel_1_1; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_1_1 <= _GEN_213;
      end
    end else begin
      states_3_vc_sel_1_1 <= _GEN_213;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_1_2 <= io_vcalloc_resp_vc_sel_1_2; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_1_2 <= _GEN_214;
      end
    end else begin
      states_3_vc_sel_1_2 <= _GEN_214;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_1_3 <= io_vcalloc_resp_vc_sel_1_3; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_1_3 <= _GEN_215;
      end
    end else begin
      states_3_vc_sel_1_3 <= _GEN_215;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_0_0 <= io_vcalloc_resp_vc_sel_0_0; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_0_0 <= _GEN_216;
      end
    end else begin
      states_3_vc_sel_0_0 <= _GEN_216;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_0_1 <= io_vcalloc_resp_vc_sel_0_1; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_0_1 <= _GEN_217;
      end
    end else begin
      states_3_vc_sel_0_1 <= _GEN_217;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_0_2 <= io_vcalloc_resp_vc_sel_0_2; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_0_2 <= _GEN_218;
      end
    end else begin
      states_3_vc_sel_0_2 <= _GEN_218;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_0_3 <= io_vcalloc_resp_vc_sel_0_3; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_0_3 <= _GEN_219;
      end
    end else begin
      states_3_vc_sel_0_3 <= _GEN_219;
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h3 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_3_flow_ingress_node <= io_in_flit_0_bits_flow_ingress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h3 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_3_flow_egress_node <= io_in_flit_0_bits_flow_egress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (reset) begin // @[InputUnit.scala 233:21]
      mask <= 4'h0; // @[InputUnit.scala 233:21]
    end else if (io_router_req_valid) begin // @[InputUnit.scala 239:31]
      mask <= _mask_T_2; // @[InputUnit.scala 240:10]
    end else if (_T_26) begin // @[InputUnit.scala 241:34]
      mask <= _mask_T_17; // @[InputUnit.scala 242:10]
    end
    salloc_outs_0_valid <= salloc_arb_io_out_0_ready & salloc_arb_io_out_0_valid; // @[Decoupled.scala 51:35]
    salloc_outs_0_out_vid <= _virt_channel_T_10 | _virt_channel_T_11; // @[Mux.scala 27:73]
    salloc_outs_0_flit_head <= salloc_arb_io_chosen_oh_0[0] & input_buffer_io_deq_0_bits_head |
      salloc_arb_io_chosen_oh_0[1] & input_buffer_io_deq_1_bits_head | salloc_arb_io_chosen_oh_0[2] &
      input_buffer_io_deq_2_bits_head | salloc_arb_io_chosen_oh_0[3] & input_buffer_io_deq_3_bits_head; // @[Mux.scala 27:73]
    salloc_outs_0_flit_tail <= salloc_arb_io_chosen_oh_0[0] & input_buffer_io_deq_0_bits_tail |
      salloc_arb_io_chosen_oh_0[1] & input_buffer_io_deq_1_bits_tail | salloc_arb_io_chosen_oh_0[2] &
      input_buffer_io_deq_2_bits_tail | salloc_arb_io_chosen_oh_0[3] & input_buffer_io_deq_3_bits_tail; // @[Mux.scala 27:73]
    salloc_outs_0_flit_payload <= _salloc_outs_0_flit_payload_T_9 | _salloc_outs_0_flit_payload_T_7; // @[Mux.scala 27:73]
    salloc_outs_0_flit_flow_ingress_node <= _salloc_outs_0_flit_flow_T_30 | _salloc_outs_0_flit_flow_T_28; // @[Mux.scala 27:73]
    salloc_outs_0_flit_flow_egress_node <= _salloc_outs_0_flit_flow_T_16 | _salloc_outs_0_flit_flow_T_14; // @[Mux.scala 27:73]
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T & _T_3 & ~(_GEN_3 == 3'h0)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:197 assert(states(id).g === g_i)\n"); // @[InputUnit.scala 197:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_router_req_valid & _T_3 & ~(_GEN_139 == 3'h1)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:224 assert(states(id).g === g_r)\n"); // @[InputUnit.scala 224:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_39 & vcalloc_sel[0] & _T_3 & ~vcalloc_vals_0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:274 assert(states(i).g === g_v)\n"); // @[InputUnit.scala 274:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_39 & vcalloc_sel[1] & _T_3 & ~vcalloc_vals_1) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:274 assert(states(i).g === g_v)\n"); // @[InputUnit.scala 274:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_39 & vcalloc_sel[2] & _T_3 & ~vcalloc_vals_2) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:274 assert(states(i).g === g_v)\n"); // @[InputUnit.scala 274:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_39 & vcalloc_sel[3] & _T_3 & ~vcalloc_vals_3) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:274 assert(states(i).g === g_v)\n"); // @[InputUnit.scala 274:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  states_0_g = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  states_0_vc_sel_2_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  states_0_vc_sel_1_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  states_0_vc_sel_0_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  states_0_flow_ingress_node = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  states_0_flow_egress_node = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  states_1_g = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  states_1_vc_sel_2_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  states_1_vc_sel_1_1 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  states_1_vc_sel_0_0 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  states_1_vc_sel_0_1 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  states_1_flow_ingress_node = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  states_1_flow_egress_node = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  states_2_g = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  states_2_vc_sel_2_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  states_2_vc_sel_1_1 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  states_2_vc_sel_1_2 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  states_2_vc_sel_0_0 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  states_2_vc_sel_0_1 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  states_2_vc_sel_0_2 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  states_2_flow_ingress_node = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  states_2_flow_egress_node = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  states_3_g = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  states_3_vc_sel_2_0 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  states_3_vc_sel_1_1 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  states_3_vc_sel_1_2 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  states_3_vc_sel_1_3 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  states_3_vc_sel_0_0 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  states_3_vc_sel_0_1 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  states_3_vc_sel_0_2 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  states_3_vc_sel_0_3 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  states_3_flow_ingress_node = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  states_3_flow_egress_node = _RAND_32[1:0];
  _RAND_33 = {1{`RANDOM}};
  mask = _RAND_33[3:0];
  _RAND_34 = {1{`RANDOM}};
  salloc_outs_0_valid = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  salloc_outs_0_out_vid = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  salloc_outs_0_flit_head = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  salloc_outs_0_flit_tail = _RAND_37[0:0];
  _RAND_38 = {2{`RANDOM}};
  salloc_outs_0_flit_payload = _RAND_38[63:0];
  _RAND_39 = {1{`RANDOM}};
  salloc_outs_0_flit_flow_ingress_node = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  salloc_outs_0_flit_flow_egress_node = _RAND_40[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (_T & ~reset) begin
      assert(1'h1); // @[InputUnit.scala 196:13]
    end
    //
    if (_T & _T_3) begin
      assert(_GEN_3 == 3'h0); // @[InputUnit.scala 197:13]
    end
    //
    if (io_router_req_valid & _T_3) begin
      assert(_GEN_139 == 3'h1); // @[InputUnit.scala 224:11]
    end
    //
    if (_T_39 & vcalloc_sel[0] & _T_3) begin
      assert(vcalloc_vals_0); // @[InputUnit.scala 274:17]
    end
    //
    if (_T_39 & vcalloc_sel[1] & _T_3) begin
      assert(vcalloc_vals_1); // @[InputUnit.scala 274:17]
    end
    //
    if (_T_39 & vcalloc_sel[2] & _T_3) begin
      assert(vcalloc_vals_2); // @[InputUnit.scala 274:17]
    end
    //
    if (_T_39 & vcalloc_sel[3] & _T_3) begin
      assert(vcalloc_vals_3); // @[InputUnit.scala 274:17]
    end
  end
endmodule
module IngressUnit_1(
  input         clock,
  input         reset,
  output        io_router_req_valid,
  output [1:0]  io_router_req_bits_flow_ingress_node,
  output [1:0]  io_router_req_bits_flow_egress_node,
  input         io_router_resp_vc_sel_1_0,
  input         io_router_resp_vc_sel_1_1,
  input         io_router_resp_vc_sel_1_2,
  input         io_router_resp_vc_sel_1_3,
  input         io_router_resp_vc_sel_0_0,
  input         io_router_resp_vc_sel_0_1,
  input         io_router_resp_vc_sel_0_2,
  input         io_router_resp_vc_sel_0_3,
  input         io_vcalloc_req_ready,
  output        io_vcalloc_req_valid,
  output        io_vcalloc_req_bits_vc_sel_2_0,
  output        io_vcalloc_req_bits_vc_sel_1_0,
  output        io_vcalloc_req_bits_vc_sel_1_1,
  output        io_vcalloc_req_bits_vc_sel_1_2,
  output        io_vcalloc_req_bits_vc_sel_1_3,
  output        io_vcalloc_req_bits_vc_sel_0_0,
  output        io_vcalloc_req_bits_vc_sel_0_1,
  output        io_vcalloc_req_bits_vc_sel_0_2,
  output        io_vcalloc_req_bits_vc_sel_0_3,
  input         io_vcalloc_resp_vc_sel_2_0,
  input         io_vcalloc_resp_vc_sel_1_0,
  input         io_vcalloc_resp_vc_sel_1_1,
  input         io_vcalloc_resp_vc_sel_1_2,
  input         io_vcalloc_resp_vc_sel_1_3,
  input         io_vcalloc_resp_vc_sel_0_0,
  input         io_vcalloc_resp_vc_sel_0_1,
  input         io_vcalloc_resp_vc_sel_0_2,
  input         io_vcalloc_resp_vc_sel_0_3,
  input         io_out_credit_available_2_0,
  input         io_out_credit_available_1_0,
  input         io_out_credit_available_1_1,
  input         io_out_credit_available_1_2,
  input         io_out_credit_available_1_3,
  input         io_out_credit_available_0_0,
  input         io_out_credit_available_0_1,
  input         io_out_credit_available_0_2,
  input         io_out_credit_available_0_3,
  input         io_salloc_req_0_ready,
  output        io_salloc_req_0_valid,
  output        io_salloc_req_0_bits_vc_sel_2_0,
  output        io_salloc_req_0_bits_vc_sel_1_0,
  output        io_salloc_req_0_bits_vc_sel_1_1,
  output        io_salloc_req_0_bits_vc_sel_1_2,
  output        io_salloc_req_0_bits_vc_sel_1_3,
  output        io_salloc_req_0_bits_vc_sel_0_0,
  output        io_salloc_req_0_bits_vc_sel_0_1,
  output        io_salloc_req_0_bits_vc_sel_0_2,
  output        io_salloc_req_0_bits_vc_sel_0_3,
  output        io_salloc_req_0_bits_tail,
  output        io_out_0_valid,
  output        io_out_0_bits_flit_head,
  output        io_out_0_bits_flit_tail,
  output [63:0] io_out_0_bits_flit_payload,
  output [1:0]  io_out_0_bits_flit_flow_ingress_node,
  output [1:0]  io_out_0_bits_flit_flow_egress_node,
  output [1:0]  io_out_0_bits_out_virt_channel,
  output        io_in_ready,
  input         io_in_valid,
  input         io_in_bits_head,
  input         io_in_bits_tail,
  input  [63:0] io_in_bits_payload,
  input  [1:0]  io_in_bits_egress_id
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  route_buffer_clock; // @[IngressUnit.scala 26:28]
  wire  route_buffer_reset; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_enq_ready; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_enq_valid; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_enq_bits_head; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_enq_bits_tail; // @[IngressUnit.scala 26:28]
  wire [63:0] route_buffer_io_enq_bits_payload; // @[IngressUnit.scala 26:28]
  wire [1:0] route_buffer_io_enq_bits_flow_ingress_node; // @[IngressUnit.scala 26:28]
  wire [1:0] route_buffer_io_enq_bits_flow_egress_node; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_deq_ready; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_deq_valid; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_deq_bits_head; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_deq_bits_tail; // @[IngressUnit.scala 26:28]
  wire [63:0] route_buffer_io_deq_bits_payload; // @[IngressUnit.scala 26:28]
  wire [1:0] route_buffer_io_deq_bits_flow_ingress_node; // @[IngressUnit.scala 26:28]
  wire [1:0] route_buffer_io_deq_bits_flow_egress_node; // @[IngressUnit.scala 26:28]
  wire  route_q_clock; // @[IngressUnit.scala 27:23]
  wire  route_q_reset; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_ready; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_valid; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_2_0; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_1_0; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_1_1; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_1_2; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_1_3; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_0_0; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_0_1; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_0_2; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_0_3; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_ready; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_valid; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_2_0; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_1_0; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_1_1; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_1_2; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_1_3; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_0_0; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_0_1; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_0_2; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_0_3; // @[IngressUnit.scala 27:23]
  wire  vcalloc_buffer_clock; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_reset; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_enq_ready; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_enq_valid; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_enq_bits_head; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_enq_bits_tail; // @[IngressUnit.scala 75:30]
  wire [63:0] vcalloc_buffer_io_enq_bits_payload; // @[IngressUnit.scala 75:30]
  wire [1:0] vcalloc_buffer_io_enq_bits_flow_ingress_node; // @[IngressUnit.scala 75:30]
  wire [1:0] vcalloc_buffer_io_enq_bits_flow_egress_node; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_deq_ready; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_deq_valid; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_deq_bits_head; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_deq_bits_tail; // @[IngressUnit.scala 75:30]
  wire [63:0] vcalloc_buffer_io_deq_bits_payload; // @[IngressUnit.scala 75:30]
  wire [1:0] vcalloc_buffer_io_deq_bits_flow_ingress_node; // @[IngressUnit.scala 75:30]
  wire [1:0] vcalloc_buffer_io_deq_bits_flow_egress_node; // @[IngressUnit.scala 75:30]
  wire  vcalloc_q_clock; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_reset; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_ready; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_valid; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_2_0; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_1_0; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_1_1; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_1_2; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_1_3; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_0_0; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_0_1; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_0_2; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_0_3; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_ready; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_valid; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_2_0; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_1_0; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_1_1; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_1_2; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_1_3; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_0_0; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_0_1; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_0_2; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_0_3; // @[IngressUnit.scala 76:25]
  wire  _T = 2'h0 == io_in_bits_egress_id; // @[IngressUnit.scala 30:72]
  wire  _T_1 = 2'h1 == io_in_bits_egress_id; // @[IngressUnit.scala 30:72]
  wire  _T_2 = 2'h2 == io_in_bits_egress_id; // @[IngressUnit.scala 30:72]
  wire  _T_3 = 2'h3 == io_in_bits_egress_id; // @[IngressUnit.scala 30:72]
  wire  _T_6 = _T | _T_1 | _T_2 | _T_3; // @[package.scala 73:59]
  wire  _T_11 = ~reset; // @[IngressUnit.scala 30:9]
  wire [1:0] _route_buffer_io_enq_bits_flow_egress_node_T_6 = _T_2 ? 2'h2 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _route_buffer_io_enq_bits_flow_egress_node_T_7 = _T_3 ? 2'h3 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _GEN_11 = {{1'd0}, _T_1}; // @[Mux.scala 27:73]
  wire [1:0] _route_buffer_io_enq_bits_flow_egress_node_T_9 = _GEN_11 | _route_buffer_io_enq_bits_flow_egress_node_T_6; // @[Mux.scala 27:73]
  wire  at_dest = route_buffer_io_enq_bits_flow_egress_node == 2'h1; // @[IngressUnit.scala 55:59]
  wire  _T_13 = io_in_ready & io_in_valid; // @[Decoupled.scala 51:35]
  wire  _vcalloc_buffer_io_enq_valid_T = ~route_buffer_io_deq_bits_head; // @[IngressUnit.scala 88:30]
  wire  _vcalloc_buffer_io_enq_valid_T_1 = route_q_io_deq_valid | ~route_buffer_io_deq_bits_head; // @[IngressUnit.scala 88:27]
  wire  _vcalloc_buffer_io_enq_valid_T_2 = route_buffer_io_deq_valid & _vcalloc_buffer_io_enq_valid_T_1; // @[IngressUnit.scala 87:61]
  wire  _vcalloc_buffer_io_enq_valid_T_4 = io_vcalloc_req_ready | _vcalloc_buffer_io_enq_valid_T; // @[IngressUnit.scala 89:27]
  wire  _io_vcalloc_req_valid_T_1 = route_buffer_io_deq_valid & route_q_io_deq_valid & route_buffer_io_deq_bits_head; // @[IngressUnit.scala 91:78]
  wire  _route_buffer_io_deq_ready_T_2 = vcalloc_buffer_io_enq_ready & _vcalloc_buffer_io_enq_valid_T_1; // @[IngressUnit.scala 93:61]
  wire  _route_buffer_io_deq_ready_T_5 = _route_buffer_io_deq_ready_T_2 & _vcalloc_buffer_io_enq_valid_T_4; // @[IngressUnit.scala 94:37]
  wire  _route_buffer_io_deq_ready_T_7 = vcalloc_q_io_enq_ready | _vcalloc_buffer_io_enq_valid_T; // @[IngressUnit.scala 96:29]
  wire  _route_q_io_deq_ready_T = route_buffer_io_deq_ready & route_buffer_io_deq_valid; // @[Decoupled.scala 51:35]
  wire [3:0] c_lo = {vcalloc_q_io_deq_bits_vc_sel_0_3,vcalloc_q_io_deq_bits_vc_sel_0_2,vcalloc_q_io_deq_bits_vc_sel_0_1,
    vcalloc_q_io_deq_bits_vc_sel_0_0}; // @[IngressUnit.scala 107:41]
  wire [8:0] _c_T = {vcalloc_q_io_deq_bits_vc_sel_2_0,vcalloc_q_io_deq_bits_vc_sel_1_3,vcalloc_q_io_deq_bits_vc_sel_1_2,
    vcalloc_q_io_deq_bits_vc_sel_1_1,vcalloc_q_io_deq_bits_vc_sel_1_0,vcalloc_q_io_deq_bits_vc_sel_0_3,
    vcalloc_q_io_deq_bits_vc_sel_0_2,vcalloc_q_io_deq_bits_vc_sel_0_1,vcalloc_q_io_deq_bits_vc_sel_0_0}; // @[IngressUnit.scala 107:41]
  wire [8:0] _c_T_1 = {io_out_credit_available_2_0,io_out_credit_available_1_3,io_out_credit_available_1_2,
    io_out_credit_available_1_1,io_out_credit_available_1_0,io_out_credit_available_0_3,io_out_credit_available_0_2,
    io_out_credit_available_0_1,io_out_credit_available_0_0}; // @[IngressUnit.scala 107:74]
  wire [8:0] _c_T_2 = _c_T & _c_T_1; // @[IngressUnit.scala 107:48]
  wire  c = _c_T_2 != 9'h0; // @[IngressUnit.scala 107:82]
  wire  _vcalloc_q_io_deq_ready_T = vcalloc_buffer_io_deq_ready & vcalloc_buffer_io_deq_valid; // @[Decoupled.scala 51:35]
  reg  out_bundle_valid; // @[IngressUnit.scala 116:8]
  reg  out_bundle_bits_flit_head; // @[IngressUnit.scala 116:8]
  reg  out_bundle_bits_flit_tail; // @[IngressUnit.scala 116:8]
  reg [63:0] out_bundle_bits_flit_payload; // @[IngressUnit.scala 116:8]
  reg [1:0] out_bundle_bits_flit_flow_ingress_node; // @[IngressUnit.scala 116:8]
  reg [1:0] out_bundle_bits_flit_flow_egress_node; // @[IngressUnit.scala 116:8]
  reg [1:0] out_bundle_bits_out_virt_channel; // @[IngressUnit.scala 116:8]
  wire  out_channel_oh_0 = vcalloc_q_io_deq_bits_vc_sel_0_0 | vcalloc_q_io_deq_bits_vc_sel_0_1 |
    vcalloc_q_io_deq_bits_vc_sel_0_2 | vcalloc_q_io_deq_bits_vc_sel_0_3; // @[IngressUnit.scala 123:67]
  wire  out_channel_oh_1 = vcalloc_q_io_deq_bits_vc_sel_1_0 | vcalloc_q_io_deq_bits_vc_sel_1_1 |
    vcalloc_q_io_deq_bits_vc_sel_1_2 | vcalloc_q_io_deq_bits_vc_sel_1_3; // @[IngressUnit.scala 123:67]
  wire [1:0] out_bundle_bits_out_virt_channel_hi_1 = c_lo[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] out_bundle_bits_out_virt_channel_lo_1 = c_lo[1:0]; // @[OneHot.scala 31:18]
  wire  _out_bundle_bits_out_virt_channel_T_1 = |out_bundle_bits_out_virt_channel_hi_1; // @[OneHot.scala 32:14]
  wire [1:0] _out_bundle_bits_out_virt_channel_T_2 = out_bundle_bits_out_virt_channel_hi_1 |
    out_bundle_bits_out_virt_channel_lo_1; // @[OneHot.scala 32:28]
  wire [1:0] _out_bundle_bits_out_virt_channel_T_4 = {_out_bundle_bits_out_virt_channel_T_1,
    _out_bundle_bits_out_virt_channel_T_2[1]}; // @[Cat.scala 33:92]
  wire [3:0] _out_bundle_bits_out_virt_channel_T_5 = {vcalloc_q_io_deq_bits_vc_sel_1_3,vcalloc_q_io_deq_bits_vc_sel_1_2,
    vcalloc_q_io_deq_bits_vc_sel_1_1,vcalloc_q_io_deq_bits_vc_sel_1_0}; // @[OneHot.scala 22:45]
  wire [1:0] out_bundle_bits_out_virt_channel_hi_3 = _out_bundle_bits_out_virt_channel_T_5[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] out_bundle_bits_out_virt_channel_lo_3 = _out_bundle_bits_out_virt_channel_T_5[1:0]; // @[OneHot.scala 31:18]
  wire  _out_bundle_bits_out_virt_channel_T_6 = |out_bundle_bits_out_virt_channel_hi_3; // @[OneHot.scala 32:14]
  wire [1:0] _out_bundle_bits_out_virt_channel_T_7 = out_bundle_bits_out_virt_channel_hi_3 |
    out_bundle_bits_out_virt_channel_lo_3; // @[OneHot.scala 32:28]
  wire [1:0] _out_bundle_bits_out_virt_channel_T_9 = {_out_bundle_bits_out_virt_channel_T_6,
    _out_bundle_bits_out_virt_channel_T_7[1]}; // @[Cat.scala 33:92]
  wire [1:0] _out_bundle_bits_out_virt_channel_T_10 = out_channel_oh_0 ? _out_bundle_bits_out_virt_channel_T_4 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _out_bundle_bits_out_virt_channel_T_11 = out_channel_oh_1 ? _out_bundle_bits_out_virt_channel_T_9 : 2'h0; // @[Mux.scala 27:73]
  Queue_8 route_buffer ( // @[IngressUnit.scala 26:28]
    .clock(route_buffer_clock),
    .reset(route_buffer_reset),
    .io_enq_ready(route_buffer_io_enq_ready),
    .io_enq_valid(route_buffer_io_enq_valid),
    .io_enq_bits_head(route_buffer_io_enq_bits_head),
    .io_enq_bits_tail(route_buffer_io_enq_bits_tail),
    .io_enq_bits_payload(route_buffer_io_enq_bits_payload),
    .io_enq_bits_flow_ingress_node(route_buffer_io_enq_bits_flow_ingress_node),
    .io_enq_bits_flow_egress_node(route_buffer_io_enq_bits_flow_egress_node),
    .io_deq_ready(route_buffer_io_deq_ready),
    .io_deq_valid(route_buffer_io_deq_valid),
    .io_deq_bits_head(route_buffer_io_deq_bits_head),
    .io_deq_bits_tail(route_buffer_io_deq_bits_tail),
    .io_deq_bits_payload(route_buffer_io_deq_bits_payload),
    .io_deq_bits_flow_ingress_node(route_buffer_io_deq_bits_flow_ingress_node),
    .io_deq_bits_flow_egress_node(route_buffer_io_deq_bits_flow_egress_node)
  );
  Queue_9 route_q ( // @[IngressUnit.scala 27:23]
    .clock(route_q_clock),
    .reset(route_q_reset),
    .io_enq_ready(route_q_io_enq_ready),
    .io_enq_valid(route_q_io_enq_valid),
    .io_enq_bits_vc_sel_2_0(route_q_io_enq_bits_vc_sel_2_0),
    .io_enq_bits_vc_sel_1_0(route_q_io_enq_bits_vc_sel_1_0),
    .io_enq_bits_vc_sel_1_1(route_q_io_enq_bits_vc_sel_1_1),
    .io_enq_bits_vc_sel_1_2(route_q_io_enq_bits_vc_sel_1_2),
    .io_enq_bits_vc_sel_1_3(route_q_io_enq_bits_vc_sel_1_3),
    .io_enq_bits_vc_sel_0_0(route_q_io_enq_bits_vc_sel_0_0),
    .io_enq_bits_vc_sel_0_1(route_q_io_enq_bits_vc_sel_0_1),
    .io_enq_bits_vc_sel_0_2(route_q_io_enq_bits_vc_sel_0_2),
    .io_enq_bits_vc_sel_0_3(route_q_io_enq_bits_vc_sel_0_3),
    .io_deq_ready(route_q_io_deq_ready),
    .io_deq_valid(route_q_io_deq_valid),
    .io_deq_bits_vc_sel_2_0(route_q_io_deq_bits_vc_sel_2_0),
    .io_deq_bits_vc_sel_1_0(route_q_io_deq_bits_vc_sel_1_0),
    .io_deq_bits_vc_sel_1_1(route_q_io_deq_bits_vc_sel_1_1),
    .io_deq_bits_vc_sel_1_2(route_q_io_deq_bits_vc_sel_1_2),
    .io_deq_bits_vc_sel_1_3(route_q_io_deq_bits_vc_sel_1_3),
    .io_deq_bits_vc_sel_0_0(route_q_io_deq_bits_vc_sel_0_0),
    .io_deq_bits_vc_sel_0_1(route_q_io_deq_bits_vc_sel_0_1),
    .io_deq_bits_vc_sel_0_2(route_q_io_deq_bits_vc_sel_0_2),
    .io_deq_bits_vc_sel_0_3(route_q_io_deq_bits_vc_sel_0_3)
  );
  Queue_8 vcalloc_buffer ( // @[IngressUnit.scala 75:30]
    .clock(vcalloc_buffer_clock),
    .reset(vcalloc_buffer_reset),
    .io_enq_ready(vcalloc_buffer_io_enq_ready),
    .io_enq_valid(vcalloc_buffer_io_enq_valid),
    .io_enq_bits_head(vcalloc_buffer_io_enq_bits_head),
    .io_enq_bits_tail(vcalloc_buffer_io_enq_bits_tail),
    .io_enq_bits_payload(vcalloc_buffer_io_enq_bits_payload),
    .io_enq_bits_flow_ingress_node(vcalloc_buffer_io_enq_bits_flow_ingress_node),
    .io_enq_bits_flow_egress_node(vcalloc_buffer_io_enq_bits_flow_egress_node),
    .io_deq_ready(vcalloc_buffer_io_deq_ready),
    .io_deq_valid(vcalloc_buffer_io_deq_valid),
    .io_deq_bits_head(vcalloc_buffer_io_deq_bits_head),
    .io_deq_bits_tail(vcalloc_buffer_io_deq_bits_tail),
    .io_deq_bits_payload(vcalloc_buffer_io_deq_bits_payload),
    .io_deq_bits_flow_ingress_node(vcalloc_buffer_io_deq_bits_flow_ingress_node),
    .io_deq_bits_flow_egress_node(vcalloc_buffer_io_deq_bits_flow_egress_node)
  );
  Queue_11 vcalloc_q ( // @[IngressUnit.scala 76:25]
    .clock(vcalloc_q_clock),
    .reset(vcalloc_q_reset),
    .io_enq_ready(vcalloc_q_io_enq_ready),
    .io_enq_valid(vcalloc_q_io_enq_valid),
    .io_enq_bits_vc_sel_2_0(vcalloc_q_io_enq_bits_vc_sel_2_0),
    .io_enq_bits_vc_sel_1_0(vcalloc_q_io_enq_bits_vc_sel_1_0),
    .io_enq_bits_vc_sel_1_1(vcalloc_q_io_enq_bits_vc_sel_1_1),
    .io_enq_bits_vc_sel_1_2(vcalloc_q_io_enq_bits_vc_sel_1_2),
    .io_enq_bits_vc_sel_1_3(vcalloc_q_io_enq_bits_vc_sel_1_3),
    .io_enq_bits_vc_sel_0_0(vcalloc_q_io_enq_bits_vc_sel_0_0),
    .io_enq_bits_vc_sel_0_1(vcalloc_q_io_enq_bits_vc_sel_0_1),
    .io_enq_bits_vc_sel_0_2(vcalloc_q_io_enq_bits_vc_sel_0_2),
    .io_enq_bits_vc_sel_0_3(vcalloc_q_io_enq_bits_vc_sel_0_3),
    .io_deq_ready(vcalloc_q_io_deq_ready),
    .io_deq_valid(vcalloc_q_io_deq_valid),
    .io_deq_bits_vc_sel_2_0(vcalloc_q_io_deq_bits_vc_sel_2_0),
    .io_deq_bits_vc_sel_1_0(vcalloc_q_io_deq_bits_vc_sel_1_0),
    .io_deq_bits_vc_sel_1_1(vcalloc_q_io_deq_bits_vc_sel_1_1),
    .io_deq_bits_vc_sel_1_2(vcalloc_q_io_deq_bits_vc_sel_1_2),
    .io_deq_bits_vc_sel_1_3(vcalloc_q_io_deq_bits_vc_sel_1_3),
    .io_deq_bits_vc_sel_0_0(vcalloc_q_io_deq_bits_vc_sel_0_0),
    .io_deq_bits_vc_sel_0_1(vcalloc_q_io_deq_bits_vc_sel_0_1),
    .io_deq_bits_vc_sel_0_2(vcalloc_q_io_deq_bits_vc_sel_0_2),
    .io_deq_bits_vc_sel_0_3(vcalloc_q_io_deq_bits_vc_sel_0_3)
  );
  assign io_router_req_valid = io_in_valid & route_buffer_io_enq_ready & io_in_bits_head & ~at_dest; // @[IngressUnit.scala 58:86]
  assign io_router_req_bits_flow_ingress_node = route_buffer_io_enq_bits_flow_ingress_node; // @[IngressUnit.scala 53:27]
  assign io_router_req_bits_flow_egress_node = route_buffer_io_enq_bits_flow_egress_node; // @[IngressUnit.scala 53:27]
  assign io_vcalloc_req_valid = _io_vcalloc_req_valid_T_1 & vcalloc_buffer_io_enq_ready & vcalloc_q_io_enq_ready; // @[IngressUnit.scala 92:41]
  assign io_vcalloc_req_bits_vc_sel_2_0 = route_q_io_deq_bits_vc_sel_2_0; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_1_0 = route_q_io_deq_bits_vc_sel_1_0; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_1_1 = route_q_io_deq_bits_vc_sel_1_1; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_1_2 = route_q_io_deq_bits_vc_sel_1_2; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_1_3 = route_q_io_deq_bits_vc_sel_1_3; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_0_0 = route_q_io_deq_bits_vc_sel_0_0; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_0_1 = route_q_io_deq_bits_vc_sel_0_1; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_0_2 = route_q_io_deq_bits_vc_sel_0_2; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_0_3 = route_q_io_deq_bits_vc_sel_0_3; // @[IngressUnit.scala 81:30]
  assign io_salloc_req_0_valid = vcalloc_buffer_io_deq_valid & vcalloc_q_io_deq_valid & c; // @[IngressUnit.scala 109:83]
  assign io_salloc_req_0_bits_vc_sel_2_0 = vcalloc_q_io_deq_bits_vc_sel_2_0; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_1_0 = vcalloc_q_io_deq_bits_vc_sel_1_0; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_1_1 = vcalloc_q_io_deq_bits_vc_sel_1_1; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_1_2 = vcalloc_q_io_deq_bits_vc_sel_1_2; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_1_3 = vcalloc_q_io_deq_bits_vc_sel_1_3; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_0_0 = vcalloc_q_io_deq_bits_vc_sel_0_0; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_0_1 = vcalloc_q_io_deq_bits_vc_sel_0_1; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_0_2 = vcalloc_q_io_deq_bits_vc_sel_0_2; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_0_3 = vcalloc_q_io_deq_bits_vc_sel_0_3; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_tail = vcalloc_buffer_io_deq_bits_tail; // @[IngressUnit.scala 105:30]
  assign io_out_0_valid = out_bundle_valid; // @[IngressUnit.scala 118:13]
  assign io_out_0_bits_flit_head = out_bundle_bits_flit_head; // @[IngressUnit.scala 118:13]
  assign io_out_0_bits_flit_tail = out_bundle_bits_flit_tail; // @[IngressUnit.scala 118:13]
  assign io_out_0_bits_flit_payload = out_bundle_bits_flit_payload; // @[IngressUnit.scala 118:13]
  assign io_out_0_bits_flit_flow_ingress_node = out_bundle_bits_flit_flow_ingress_node; // @[IngressUnit.scala 118:13]
  assign io_out_0_bits_flit_flow_egress_node = out_bundle_bits_flit_flow_egress_node; // @[IngressUnit.scala 118:13]
  assign io_out_0_bits_out_virt_channel = out_bundle_bits_out_virt_channel; // @[IngressUnit.scala 118:13]
  assign io_in_ready = route_buffer_io_enq_ready; // @[IngressUnit.scala 59:44]
  assign route_buffer_clock = clock;
  assign route_buffer_reset = reset;
  assign route_buffer_io_enq_valid = io_in_valid; // @[IngressUnit.scala 56:44]
  assign route_buffer_io_enq_bits_head = io_in_bits_head; // @[IngressUnit.scala 32:33]
  assign route_buffer_io_enq_bits_tail = io_in_bits_tail; // @[IngressUnit.scala 33:33]
  assign route_buffer_io_enq_bits_payload = io_in_bits_payload; // @[IngressUnit.scala 50:36]
  assign route_buffer_io_enq_bits_flow_ingress_node = 2'h1; // @[IngressUnit.scala 38:51]
  assign route_buffer_io_enq_bits_flow_egress_node = _route_buffer_io_enq_bits_flow_egress_node_T_9 |
    _route_buffer_io_enq_bits_flow_egress_node_T_7; // @[Mux.scala 27:73]
  assign route_buffer_io_deq_ready = _route_buffer_io_deq_ready_T_5 & _route_buffer_io_deq_ready_T_7; // @[IngressUnit.scala 95:37]
  assign route_q_clock = clock;
  assign route_q_reset = reset;
  assign route_q_io_enq_valid = _T_13 & io_in_bits_head & at_dest | io_router_req_valid; // @[IngressUnit.scala 62:24 64:53 65:26]
  assign route_q_io_enq_bits_vc_sel_2_0 = _T_13 & io_in_bits_head & at_dest & _T_1; // @[IngressUnit.scala 63:23 64:53]
  assign route_q_io_enq_bits_vc_sel_1_0 = _T_13 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_1_0; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_1_1 = _T_13 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_1_1; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_1_2 = _T_13 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_1_2; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_1_3 = _T_13 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_1_3; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_0_0 = _T_13 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_0_0; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_0_1 = _T_13 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_0_1; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_0_2 = _T_13 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_0_2; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_0_3 = _T_13 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_0_3; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_deq_ready = _route_q_io_deq_ready_T & route_buffer_io_deq_bits_tail; // @[IngressUnit.scala 97:55]
  assign vcalloc_buffer_clock = clock;
  assign vcalloc_buffer_reset = reset;
  assign vcalloc_buffer_io_enq_valid = _vcalloc_buffer_io_enq_valid_T_2 & _vcalloc_buffer_io_enq_valid_T_4; // @[IngressUnit.scala 88:37]
  assign vcalloc_buffer_io_enq_bits_head = route_buffer_io_deq_bits_head; // @[IngressUnit.scala 79:30]
  assign vcalloc_buffer_io_enq_bits_tail = route_buffer_io_deq_bits_tail; // @[IngressUnit.scala 79:30]
  assign vcalloc_buffer_io_enq_bits_payload = route_buffer_io_deq_bits_payload; // @[IngressUnit.scala 79:30]
  assign vcalloc_buffer_io_enq_bits_flow_ingress_node = route_buffer_io_deq_bits_flow_ingress_node; // @[IngressUnit.scala 79:30]
  assign vcalloc_buffer_io_enq_bits_flow_egress_node = route_buffer_io_deq_bits_flow_egress_node; // @[IngressUnit.scala 79:30]
  assign vcalloc_buffer_io_deq_ready = io_salloc_req_0_ready & vcalloc_q_io_deq_valid & c; // @[IngressUnit.scala 110:83]
  assign vcalloc_q_clock = clock;
  assign vcalloc_q_reset = reset;
  assign vcalloc_q_io_enq_valid = io_vcalloc_req_ready & io_vcalloc_req_valid; // @[Decoupled.scala 51:35]
  assign vcalloc_q_io_enq_bits_vc_sel_2_0 = io_vcalloc_resp_vc_sel_2_0; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_1_0 = io_vcalloc_resp_vc_sel_1_0; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_1_1 = io_vcalloc_resp_vc_sel_1_1; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_1_2 = io_vcalloc_resp_vc_sel_1_2; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_1_3 = io_vcalloc_resp_vc_sel_1_3; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_0_0 = io_vcalloc_resp_vc_sel_0_0; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_0_1 = io_vcalloc_resp_vc_sel_0_1; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_0_2 = io_vcalloc_resp_vc_sel_0_2; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_0_3 = io_vcalloc_resp_vc_sel_0_3; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_deq_ready = vcalloc_buffer_io_deq_bits_tail & _vcalloc_q_io_deq_ready_T; // @[IngressUnit.scala 111:42]
  always @(posedge clock) begin
    out_bundle_valid <= vcalloc_buffer_io_deq_ready & vcalloc_buffer_io_deq_valid; // @[Decoupled.scala 51:35]
    out_bundle_bits_flit_head <= vcalloc_buffer_io_deq_bits_head; // @[IngressUnit.scala 121:24]
    out_bundle_bits_flit_tail <= vcalloc_buffer_io_deq_bits_tail; // @[IngressUnit.scala 121:24]
    out_bundle_bits_flit_payload <= vcalloc_buffer_io_deq_bits_payload; // @[IngressUnit.scala 121:24]
    out_bundle_bits_flit_flow_ingress_node <= vcalloc_buffer_io_deq_bits_flow_ingress_node; // @[IngressUnit.scala 121:24]
    out_bundle_bits_flit_flow_egress_node <= vcalloc_buffer_io_deq_bits_flow_egress_node; // @[IngressUnit.scala 121:24]
    out_bundle_bits_out_virt_channel <= _out_bundle_bits_out_virt_channel_T_10 | _out_bundle_bits_out_virt_channel_T_11; // @[Mux.scala 27:73]
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~(io_in_valid & ~_T_6))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at IngressUnit.scala:30 assert(!(io.in.valid && !cParam.possibleFlows.toSeq.map(_.egressId.U === io.in.bits.egress_id).orR))\n"
            ); // @[IngressUnit.scala 30:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_11 & ~(~(route_q_io_enq_valid & ~route_q_io_enq_ready))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at IngressUnit.scala:73 assert(!(route_q.io.enq.valid && !route_q.io.enq.ready))\n"); // @[IngressUnit.scala 73:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_11 & ~(~(vcalloc_q_io_enq_valid & ~vcalloc_q_io_enq_ready))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at IngressUnit.scala:102 assert(!(vcalloc_q.io.enq.valid && !vcalloc_q.io.enq.ready))\n"
            ); // @[IngressUnit.scala 102:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  out_bundle_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  out_bundle_bits_flit_head = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  out_bundle_bits_flit_tail = _RAND_2[0:0];
  _RAND_3 = {2{`RANDOM}};
  out_bundle_bits_flit_payload = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  out_bundle_bits_flit_flow_ingress_node = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  out_bundle_bits_flit_flow_egress_node = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  out_bundle_bits_out_virt_channel = _RAND_6[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(~(io_in_valid & ~_T_6)); // @[IngressUnit.scala 30:9]
    end
    //
    if (_T_11) begin
      assert(~(route_q_io_enq_valid & ~route_q_io_enq_ready)); // @[IngressUnit.scala 73:9]
    end
    //
    if (_T_11) begin
      assert(~(vcalloc_q_io_enq_valid & ~vcalloc_q_io_enq_ready)); // @[IngressUnit.scala 102:9]
    end
  end
endmodule
module RouteComputer_1(
  input  [1:0] io_req_2_bits_flow_ingress_node,
  input  [1:0] io_req_2_bits_flow_egress_node,
  input  [1:0] io_req_1_bits_src_virt_id,
  input  [1:0] io_req_1_bits_flow_ingress_node,
  input  [1:0] io_req_1_bits_flow_egress_node,
  input  [1:0] io_req_0_bits_src_virt_id,
  input  [1:0] io_req_0_bits_flow_ingress_node,
  input  [1:0] io_req_0_bits_flow_egress_node,
  output       io_resp_2_vc_sel_1_0,
  output       io_resp_2_vc_sel_1_1,
  output       io_resp_2_vc_sel_1_2,
  output       io_resp_2_vc_sel_1_3,
  output       io_resp_2_vc_sel_0_0,
  output       io_resp_2_vc_sel_0_1,
  output       io_resp_2_vc_sel_0_2,
  output       io_resp_2_vc_sel_0_3,
  output       io_resp_1_vc_sel_1_0,
  output       io_resp_1_vc_sel_1_1,
  output       io_resp_1_vc_sel_1_2,
  output       io_resp_1_vc_sel_1_3,
  output       io_resp_1_vc_sel_0_0,
  output       io_resp_1_vc_sel_0_1,
  output       io_resp_1_vc_sel_0_2,
  output       io_resp_1_vc_sel_0_3,
  output       io_resp_0_vc_sel_1_0,
  output       io_resp_0_vc_sel_1_1,
  output       io_resp_0_vc_sel_1_2,
  output       io_resp_0_vc_sel_1_3,
  output       io_resp_0_vc_sel_0_0,
  output       io_resp_0_vc_sel_0_1,
  output       io_resp_0_vc_sel_0_2,
  output       io_resp_0_vc_sel_0_3
);
  wire [5:0] addr = {io_req_0_bits_src_virt_id,io_req_0_bits_flow_ingress_node,io_req_0_bits_flow_egress_node}; // @[RouteComputer.scala 74:27]
  wire [5:0] decoded_invInputs = ~addr; // @[pla.scala 78:21]
  wire  decoded_andMatrixInput_0 = decoded_invInputs[4]; // @[pla.scala 91:29]
  wire  decoded_andMatrixInput_1 = decoded_invInputs[5]; // @[pla.scala 91:29]
  wire [1:0] _decoded_T = {decoded_andMatrixInput_0,decoded_andMatrixInput_1}; // @[Cat.scala 33:92]
  wire  _decoded_T_1 = &_decoded_T; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_0_1 = decoded_invInputs[1]; // @[pla.scala 91:29]
  wire  decoded_andMatrixInput_1_1 = decoded_invInputs[2]; // @[pla.scala 91:29]
  wire  decoded_andMatrixInput_2 = decoded_invInputs[3]; // @[pla.scala 91:29]
  wire [4:0] _decoded_T_2 = {decoded_andMatrixInput_0_1,decoded_andMatrixInput_1_1,decoded_andMatrixInput_2,
    decoded_andMatrixInput_0,decoded_andMatrixInput_1}; // @[Cat.scala 33:92]
  wire  _decoded_T_3 = &_decoded_T_2; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_0_2 = decoded_invInputs[0]; // @[pla.scala 91:29]
  wire  decoded_andMatrixInput_1_2 = addr[1]; // @[pla.scala 90:45]
  wire [1:0] _decoded_T_4 = {decoded_andMatrixInput_0_2,decoded_andMatrixInput_1_2}; // @[Cat.scala 33:92]
  wire  _decoded_T_5 = &_decoded_T_4; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_0_3 = addr[3]; // @[pla.scala 90:45]
  wire [2:0] _decoded_T_6 = {decoded_andMatrixInput_0_3,decoded_andMatrixInput_0,decoded_andMatrixInput_1}; // @[Cat.scala 33:92]
  wire  _decoded_T_7 = &_decoded_T_6; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_1_4 = addr[4]; // @[pla.scala 90:45]
  wire [1:0] _decoded_T_8 = {decoded_andMatrixInput_1_1,decoded_andMatrixInput_1_4}; // @[Cat.scala 33:92]
  wire  _decoded_T_9 = &_decoded_T_8; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_0_5 = addr[0]; // @[pla.scala 90:45]
  wire [1:0] _decoded_T_10 = {decoded_andMatrixInput_0_5,decoded_andMatrixInput_1_4}; // @[Cat.scala 33:92]
  wire  _decoded_T_11 = &_decoded_T_10; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_1_6 = addr[5]; // @[pla.scala 90:45]
  wire [1:0] _decoded_T_12 = {decoded_andMatrixInput_1_1,decoded_andMatrixInput_1_6}; // @[Cat.scala 33:92]
  wire  _decoded_T_13 = &_decoded_T_12; // @[pla.scala 98:74]
  wire [1:0] _decoded_T_14 = {decoded_andMatrixInput_0_5,decoded_andMatrixInput_1_6}; // @[Cat.scala 33:92]
  wire  _decoded_T_15 = &_decoded_T_14; // @[pla.scala 98:74]
  wire [1:0] _decoded_T_16 = {decoded_andMatrixInput_1_4,decoded_andMatrixInput_1_6}; // @[Cat.scala 33:92]
  wire  _decoded_T_17 = &_decoded_T_16; // @[pla.scala 98:74]
  wire [4:0] _decoded_T_18 = {decoded_andMatrixInput_0_1,decoded_andMatrixInput_1_1,decoded_andMatrixInput_2,
    decoded_andMatrixInput_1_4,decoded_andMatrixInput_1_6}; // @[Cat.scala 33:92]
  wire  _decoded_T_19 = &_decoded_T_18; // @[pla.scala 98:74]
  wire [2:0] _decoded_T_20 = {decoded_andMatrixInput_0_3,decoded_andMatrixInput_1_4,decoded_andMatrixInput_1_6}; // @[Cat.scala 33:92]
  wire  _decoded_T_21 = &_decoded_T_20; // @[pla.scala 98:74]
  wire  _decoded_orMatrixOutputs_T = |_decoded_T_17; // @[pla.scala 114:39]
  wire [1:0] _decoded_orMatrixOutputs_T_1 = {_decoded_T_13,_decoded_T_15}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_2 = |_decoded_orMatrixOutputs_T_1; // @[pla.scala 114:39]
  wire [3:0] _decoded_orMatrixOutputs_T_3 = {_decoded_T_9,_decoded_T_11,_decoded_T_13,_decoded_T_15}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_4 = |_decoded_orMatrixOutputs_T_3; // @[pla.scala 114:39]
  wire [1:0] _decoded_orMatrixOutputs_T_5 = {_decoded_T_1,_decoded_T_5}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_6 = |_decoded_orMatrixOutputs_T_5; // @[pla.scala 114:39]
  wire [1:0] _decoded_orMatrixOutputs_T_7 = {_decoded_T_19,_decoded_T_21}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_8 = |_decoded_orMatrixOutputs_T_7; // @[pla.scala 114:39]
  wire  _decoded_orMatrixOutputs_T_9 = |_decoded_T_15; // @[pla.scala 114:39]
  wire [1:0] _decoded_orMatrixOutputs_T_10 = {_decoded_T_11,_decoded_T_15}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_11 = |_decoded_orMatrixOutputs_T_10; // @[pla.scala 114:39]
  wire [1:0] _decoded_orMatrixOutputs_T_12 = {_decoded_T_3,_decoded_T_7}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_13 = |_decoded_orMatrixOutputs_T_12; // @[pla.scala 114:39]
  wire [7:0] decoded_orMatrixOutputs = {_decoded_orMatrixOutputs_T_13,_decoded_orMatrixOutputs_T_11,
    _decoded_orMatrixOutputs_T_9,_decoded_orMatrixOutputs_T_8,_decoded_orMatrixOutputs_T_6,_decoded_orMatrixOutputs_T_4,
    _decoded_orMatrixOutputs_T_2,_decoded_orMatrixOutputs_T}; // @[Cat.scala 33:92]
  wire [7:0] decoded_invMatrixOutputs = {decoded_orMatrixOutputs[7],decoded_orMatrixOutputs[6],decoded_orMatrixOutputs[5
    ],decoded_orMatrixOutputs[4],decoded_orMatrixOutputs[3],decoded_orMatrixOutputs[2],decoded_orMatrixOutputs[1],
    decoded_orMatrixOutputs[0]}; // @[Cat.scala 33:92]
  wire [7:0] _GEN_0 = {{4'd0}, decoded_invMatrixOutputs[7:4]}; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_25 = _GEN_0 & 8'hf; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_27 = {decoded_invMatrixOutputs[3:0], 4'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _decoded_T_29 = _decoded_T_27 & 8'hf0; // @[Bitwise.scala 108:80]
  wire [7:0] _decoded_T_30 = _decoded_T_25 | _decoded_T_29; // @[Bitwise.scala 108:39]
  wire [7:0] _GEN_1 = {{2'd0}, _decoded_T_30[7:2]}; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_35 = _GEN_1 & 8'h33; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_37 = {_decoded_T_30[5:0], 2'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _decoded_T_39 = _decoded_T_37 & 8'hcc; // @[Bitwise.scala 108:80]
  wire [7:0] _decoded_T_40 = _decoded_T_35 | _decoded_T_39; // @[Bitwise.scala 108:39]
  wire [7:0] _GEN_2 = {{1'd0}, _decoded_T_40[7:1]}; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_45 = _GEN_2 & 8'h55; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_47 = {_decoded_T_40[6:0], 1'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _decoded_T_49 = _decoded_T_47 & 8'haa; // @[Bitwise.scala 108:80]
  wire [7:0] decoded = _decoded_T_45 | _decoded_T_49; // @[Bitwise.scala 108:39]
  wire [5:0] addr_1 = {io_req_1_bits_src_virt_id,io_req_1_bits_flow_ingress_node,io_req_1_bits_flow_egress_node}; // @[RouteComputer.scala 74:27]
  wire [5:0] decoded_invInputs_1 = ~addr_1; // @[pla.scala 78:21]
  wire  decoded_andMatrixInput_0_11 = decoded_invInputs_1[0]; // @[pla.scala 91:29]
  wire  decoded_andMatrixInput_1_11 = decoded_invInputs_1[1]; // @[pla.scala 91:29]
  wire [1:0] _decoded_T_50 = {decoded_andMatrixInput_0_11,decoded_andMatrixInput_1_11}; // @[Cat.scala 33:92]
  wire  _decoded_T_51 = &_decoded_T_50; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_0_12 = decoded_invInputs_1[4]; // @[pla.scala 91:29]
  wire  decoded_andMatrixInput_1_12 = decoded_invInputs_1[5]; // @[pla.scala 91:29]
  wire [1:0] _decoded_T_52 = {decoded_andMatrixInput_0_12,decoded_andMatrixInput_1_12}; // @[Cat.scala 33:92]
  wire  _decoded_T_53 = &_decoded_T_52; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_0_13 = addr_1[0]; // @[pla.scala 90:45]
  wire  decoded_andMatrixInput_1_13 = addr_1[3]; // @[pla.scala 90:45]
  wire [3:0] _decoded_T_54 = {decoded_andMatrixInput_0_13,decoded_andMatrixInput_1_13,decoded_andMatrixInput_0_12,
    decoded_andMatrixInput_1_12}; // @[Cat.scala 33:92]
  wire  _decoded_T_55 = &_decoded_T_54; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_1_14 = addr_1[4]; // @[pla.scala 90:45]
  wire [1:0] _decoded_T_56 = {decoded_andMatrixInput_1_11,decoded_andMatrixInput_1_14}; // @[Cat.scala 33:92]
  wire  _decoded_T_57 = &_decoded_T_56; // @[pla.scala 98:74]
  wire [3:0] _decoded_T_58 = {decoded_andMatrixInput_0_13,decoded_andMatrixInput_1_11,decoded_andMatrixInput_1_13,
    decoded_andMatrixInput_1_14}; // @[Cat.scala 33:92]
  wire  _decoded_T_59 = &_decoded_T_58; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_1_16 = addr_1[5]; // @[pla.scala 90:45]
  wire [1:0] _decoded_T_60 = {decoded_andMatrixInput_1_11,decoded_andMatrixInput_1_16}; // @[Cat.scala 33:92]
  wire  _decoded_T_61 = &_decoded_T_60; // @[pla.scala 98:74]
  wire [3:0] _decoded_T_62 = {decoded_andMatrixInput_0_13,decoded_andMatrixInput_1_11,decoded_andMatrixInput_1_13,
    decoded_andMatrixInput_1_16}; // @[Cat.scala 33:92]
  wire  _decoded_T_63 = &_decoded_T_62; // @[pla.scala 98:74]
  wire [1:0] _decoded_T_64 = {decoded_andMatrixInput_1_14,decoded_andMatrixInput_1_16}; // @[Cat.scala 33:92]
  wire  _decoded_T_65 = &_decoded_T_64; // @[pla.scala 98:74]
  wire [3:0] _decoded_T_66 = {decoded_andMatrixInput_0_13,decoded_andMatrixInput_1_13,decoded_andMatrixInput_1_14,
    decoded_andMatrixInput_1_16}; // @[Cat.scala 33:92]
  wire  _decoded_T_67 = &_decoded_T_66; // @[pla.scala 98:74]
  wire  _decoded_orMatrixOutputs_T_14 = |_decoded_T_67; // @[pla.scala 114:39]
  wire  _decoded_orMatrixOutputs_T_15 = |_decoded_T_63; // @[pla.scala 114:39]
  wire [1:0] _decoded_orMatrixOutputs_T_16 = {_decoded_T_59,_decoded_T_63}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_17 = |_decoded_orMatrixOutputs_T_16; // @[pla.scala 114:39]
  wire  _decoded_orMatrixOutputs_T_18 = |_decoded_T_55; // @[pla.scala 114:39]
  wire  _decoded_orMatrixOutputs_T_19 = |_decoded_T_65; // @[pla.scala 114:39]
  wire  _decoded_orMatrixOutputs_T_20 = |_decoded_T_61; // @[pla.scala 114:39]
  wire [1:0] _decoded_orMatrixOutputs_T_21 = {_decoded_T_57,_decoded_T_61}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_22 = |_decoded_orMatrixOutputs_T_21; // @[pla.scala 114:39]
  wire [1:0] _decoded_orMatrixOutputs_T_23 = {_decoded_T_51,_decoded_T_53}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_24 = |_decoded_orMatrixOutputs_T_23; // @[pla.scala 114:39]
  wire [7:0] decoded_orMatrixOutputs_1 = {_decoded_orMatrixOutputs_T_24,_decoded_orMatrixOutputs_T_22,
    _decoded_orMatrixOutputs_T_20,_decoded_orMatrixOutputs_T_19,_decoded_orMatrixOutputs_T_18,
    _decoded_orMatrixOutputs_T_17,_decoded_orMatrixOutputs_T_15,_decoded_orMatrixOutputs_T_14}; // @[Cat.scala 33:92]
  wire [7:0] decoded_invMatrixOutputs_1 = {decoded_orMatrixOutputs_1[7],decoded_orMatrixOutputs_1[6],
    decoded_orMatrixOutputs_1[5],decoded_orMatrixOutputs_1[4],decoded_orMatrixOutputs_1[3],decoded_orMatrixOutputs_1[2],
    decoded_orMatrixOutputs_1[1],decoded_orMatrixOutputs_1[0]}; // @[Cat.scala 33:92]
  wire [7:0] _GEN_3 = {{4'd0}, decoded_invMatrixOutputs_1[7:4]}; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_71 = _GEN_3 & 8'hf; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_73 = {decoded_invMatrixOutputs_1[3:0], 4'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _decoded_T_75 = _decoded_T_73 & 8'hf0; // @[Bitwise.scala 108:80]
  wire [7:0] _decoded_T_76 = _decoded_T_71 | _decoded_T_75; // @[Bitwise.scala 108:39]
  wire [7:0] _GEN_4 = {{2'd0}, _decoded_T_76[7:2]}; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_81 = _GEN_4 & 8'h33; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_83 = {_decoded_T_76[5:0], 2'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _decoded_T_85 = _decoded_T_83 & 8'hcc; // @[Bitwise.scala 108:80]
  wire [7:0] _decoded_T_86 = _decoded_T_81 | _decoded_T_85; // @[Bitwise.scala 108:39]
  wire [7:0] _GEN_5 = {{1'd0}, _decoded_T_86[7:1]}; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_91 = _GEN_5 & 8'h55; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_93 = {_decoded_T_86[6:0], 1'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _decoded_T_95 = _decoded_T_93 & 8'haa; // @[Bitwise.scala 108:80]
  wire [7:0] decoded_1 = _decoded_T_91 | _decoded_T_95; // @[Bitwise.scala 108:39]
  wire [5:0] addr_2 = {2'h0,io_req_2_bits_flow_ingress_node,io_req_2_bits_flow_egress_node}; // @[RouteComputer.scala 74:27]
  wire [5:0] decoded_invInputs_2 = ~addr_2; // @[pla.scala 78:21]
  wire  decoded_andMatrixInput_0_20 = decoded_invInputs_2[1]; // @[pla.scala 91:29]
  wire  decoded_andMatrixInput_1_20 = addr_2[2]; // @[pla.scala 90:45]
  wire  decoded_andMatrixInput_2_8 = decoded_invInputs_2[3]; // @[pla.scala 91:29]
  wire  decoded_andMatrixInput_3_6 = decoded_invInputs_2[4]; // @[pla.scala 91:29]
  wire  decoded_andMatrixInput_4_2 = decoded_invInputs_2[5]; // @[pla.scala 91:29]
  wire [4:0] _decoded_T_96 = {decoded_andMatrixInput_0_20,decoded_andMatrixInput_1_20,decoded_andMatrixInput_2_8,
    decoded_andMatrixInput_3_6,decoded_andMatrixInput_4_2}; // @[Cat.scala 33:92]
  wire  _decoded_T_97 = &_decoded_T_96; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_0_21 = addr_2[0]; // @[pla.scala 90:45]
  wire [4:0] _decoded_T_98 = {decoded_andMatrixInput_0_21,decoded_andMatrixInput_1_20,decoded_andMatrixInput_2_8,
    decoded_andMatrixInput_3_6,decoded_andMatrixInput_4_2}; // @[Cat.scala 33:92]
  wire  _decoded_T_99 = &_decoded_T_98; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_0_22 = addr_2[1]; // @[pla.scala 90:45]
  wire [4:0] _decoded_T_100 = {decoded_andMatrixInput_0_22,decoded_andMatrixInput_1_20,decoded_andMatrixInput_2_8,
    decoded_andMatrixInput_3_6,decoded_andMatrixInput_4_2}; // @[Cat.scala 33:92]
  wire  _decoded_T_101 = &_decoded_T_100; // @[pla.scala 98:74]
  wire [1:0] _decoded_orMatrixOutputs_T_25 = {_decoded_T_99,_decoded_T_101}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_26 = |_decoded_orMatrixOutputs_T_25; // @[pla.scala 114:39]
  wire [1:0] _decoded_orMatrixOutputs_T_31 = {_decoded_T_97,_decoded_T_99}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_32 = |_decoded_orMatrixOutputs_T_31; // @[pla.scala 114:39]
  wire [7:0] decoded_orMatrixOutputs_2 = {1'h0,_decoded_orMatrixOutputs_T_32,_decoded_orMatrixOutputs_T_32,
    _decoded_orMatrixOutputs_T_32,1'h0,_decoded_orMatrixOutputs_T_26,_decoded_orMatrixOutputs_T_26,
    _decoded_orMatrixOutputs_T_26}; // @[Cat.scala 33:92]
  wire [7:0] decoded_invMatrixOutputs_2 = {decoded_orMatrixOutputs_2[7],decoded_orMatrixOutputs_2[6],
    decoded_orMatrixOutputs_2[5],decoded_orMatrixOutputs_2[4],decoded_orMatrixOutputs_2[3],decoded_orMatrixOutputs_2[2],
    decoded_orMatrixOutputs_2[1],decoded_orMatrixOutputs_2[0]}; // @[Cat.scala 33:92]
  wire [7:0] _GEN_6 = {{4'd0}, decoded_invMatrixOutputs_2[7:4]}; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_105 = _GEN_6 & 8'hf; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_107 = {decoded_invMatrixOutputs_2[3:0], 4'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _decoded_T_109 = _decoded_T_107 & 8'hf0; // @[Bitwise.scala 108:80]
  wire [7:0] _decoded_T_110 = _decoded_T_105 | _decoded_T_109; // @[Bitwise.scala 108:39]
  wire [7:0] _GEN_7 = {{2'd0}, _decoded_T_110[7:2]}; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_115 = _GEN_7 & 8'h33; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_117 = {_decoded_T_110[5:0], 2'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _decoded_T_119 = _decoded_T_117 & 8'hcc; // @[Bitwise.scala 108:80]
  wire [7:0] _decoded_T_120 = _decoded_T_115 | _decoded_T_119; // @[Bitwise.scala 108:39]
  wire [7:0] _GEN_8 = {{1'd0}, _decoded_T_120[7:1]}; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_125 = _GEN_8 & 8'h55; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_127 = {_decoded_T_120[6:0], 1'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _decoded_T_129 = _decoded_T_127 & 8'haa; // @[Bitwise.scala 108:80]
  wire [7:0] decoded_2 = _decoded_T_125 | _decoded_T_129; // @[Bitwise.scala 108:39]
  assign io_resp_2_vc_sel_1_0 = decoded_2[4]; // @[RouteComputer.scala 90:46]
  assign io_resp_2_vc_sel_1_1 = decoded_2[5]; // @[RouteComputer.scala 90:46]
  assign io_resp_2_vc_sel_1_2 = decoded_2[6]; // @[RouteComputer.scala 90:46]
  assign io_resp_2_vc_sel_1_3 = decoded_2[7]; // @[RouteComputer.scala 90:46]
  assign io_resp_2_vc_sel_0_0 = decoded_2[0]; // @[RouteComputer.scala 90:46]
  assign io_resp_2_vc_sel_0_1 = decoded_2[1]; // @[RouteComputer.scala 90:46]
  assign io_resp_2_vc_sel_0_2 = decoded_2[2]; // @[RouteComputer.scala 90:46]
  assign io_resp_2_vc_sel_0_3 = decoded_2[3]; // @[RouteComputer.scala 90:46]
  assign io_resp_1_vc_sel_1_0 = decoded_1[4]; // @[RouteComputer.scala 90:46]
  assign io_resp_1_vc_sel_1_1 = decoded_1[5]; // @[RouteComputer.scala 90:46]
  assign io_resp_1_vc_sel_1_2 = decoded_1[6]; // @[RouteComputer.scala 90:46]
  assign io_resp_1_vc_sel_1_3 = decoded_1[7]; // @[RouteComputer.scala 90:46]
  assign io_resp_1_vc_sel_0_0 = decoded_1[0]; // @[RouteComputer.scala 90:46]
  assign io_resp_1_vc_sel_0_1 = decoded_1[1]; // @[RouteComputer.scala 90:46]
  assign io_resp_1_vc_sel_0_2 = decoded_1[2]; // @[RouteComputer.scala 90:46]
  assign io_resp_1_vc_sel_0_3 = decoded_1[3]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_1_0 = decoded[4]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_1_1 = decoded[5]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_1_2 = decoded[6]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_1_3 = decoded[7]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_0_0 = decoded[0]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_0_1 = decoded[1]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_0_2 = decoded[2]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_0_3 = decoded[3]; // @[RouteComputer.scala 90:46]
endmodule
module Router_1(
  input         clock,
  input         reset,
  output [1:0]  auto_debug_out_va_stall_0,
  output [1:0]  auto_debug_out_va_stall_1,
  output [1:0]  auto_debug_out_sa_stall_0,
  output [1:0]  auto_debug_out_sa_stall_1,
  output        auto_egress_nodes_out_flit_valid,
  output        auto_egress_nodes_out_flit_bits_head,
  output        auto_egress_nodes_out_flit_bits_tail,
  output [63:0] auto_egress_nodes_out_flit_bits_payload,
  output [1:0]  auto_egress_nodes_out_flit_bits_ingress_id,
  output        auto_ingress_nodes_in_flit_ready,
  input         auto_ingress_nodes_in_flit_valid,
  input         auto_ingress_nodes_in_flit_bits_head,
  input         auto_ingress_nodes_in_flit_bits_tail,
  input  [63:0] auto_ingress_nodes_in_flit_bits_payload,
  input  [1:0]  auto_ingress_nodes_in_flit_bits_egress_id,
  output        auto_source_nodes_out_1_flit_0_valid,
  output        auto_source_nodes_out_1_flit_0_bits_head,
  output        auto_source_nodes_out_1_flit_0_bits_tail,
  output [63:0] auto_source_nodes_out_1_flit_0_bits_payload,
  output [1:0]  auto_source_nodes_out_1_flit_0_bits_flow_ingress_node,
  output [1:0]  auto_source_nodes_out_1_flit_0_bits_flow_egress_node,
  output [1:0]  auto_source_nodes_out_1_flit_0_bits_virt_channel_id,
  input  [3:0]  auto_source_nodes_out_1_credit_return,
  input  [3:0]  auto_source_nodes_out_1_vc_free,
  output        auto_source_nodes_out_0_flit_0_valid,
  output        auto_source_nodes_out_0_flit_0_bits_head,
  output        auto_source_nodes_out_0_flit_0_bits_tail,
  output [63:0] auto_source_nodes_out_0_flit_0_bits_payload,
  output [1:0]  auto_source_nodes_out_0_flit_0_bits_flow_ingress_node,
  output [1:0]  auto_source_nodes_out_0_flit_0_bits_flow_egress_node,
  output [1:0]  auto_source_nodes_out_0_flit_0_bits_virt_channel_id,
  input  [3:0]  auto_source_nodes_out_0_credit_return,
  input  [3:0]  auto_source_nodes_out_0_vc_free,
  input         auto_dest_nodes_in_1_flit_0_valid,
  input         auto_dest_nodes_in_1_flit_0_bits_head,
  input         auto_dest_nodes_in_1_flit_0_bits_tail,
  input  [63:0] auto_dest_nodes_in_1_flit_0_bits_payload,
  input  [1:0]  auto_dest_nodes_in_1_flit_0_bits_flow_ingress_node,
  input  [1:0]  auto_dest_nodes_in_1_flit_0_bits_flow_egress_node,
  input  [1:0]  auto_dest_nodes_in_1_flit_0_bits_virt_channel_id,
  output [3:0]  auto_dest_nodes_in_1_credit_return,
  output [3:0]  auto_dest_nodes_in_1_vc_free,
  input         auto_dest_nodes_in_0_flit_0_valid,
  input         auto_dest_nodes_in_0_flit_0_bits_head,
  input         auto_dest_nodes_in_0_flit_0_bits_tail,
  input  [63:0] auto_dest_nodes_in_0_flit_0_bits_payload,
  input  [1:0]  auto_dest_nodes_in_0_flit_0_bits_flow_ingress_node,
  input  [1:0]  auto_dest_nodes_in_0_flit_0_bits_flow_egress_node,
  input  [1:0]  auto_dest_nodes_in_0_flit_0_bits_virt_channel_id,
  output [3:0]  auto_dest_nodes_in_0_credit_return,
  output [3:0]  auto_dest_nodes_in_0_vc_free
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_REG_INIT
  wire  monitor_clock; // @[Nodes.scala 24:25]
  wire  monitor_reset; // @[Nodes.scala 24:25]
  wire  monitor_io_in_flit_0_valid; // @[Nodes.scala 24:25]
  wire  monitor_io_in_flit_0_bits_head; // @[Nodes.scala 24:25]
  wire  monitor_io_in_flit_0_bits_tail; // @[Nodes.scala 24:25]
  wire [1:0] monitor_io_in_flit_0_bits_flow_ingress_node; // @[Nodes.scala 24:25]
  wire [1:0] monitor_io_in_flit_0_bits_flow_egress_node; // @[Nodes.scala 24:25]
  wire [1:0] monitor_io_in_flit_0_bits_virt_channel_id; // @[Nodes.scala 24:25]
  wire  monitor_1_clock; // @[Nodes.scala 24:25]
  wire  monitor_1_reset; // @[Nodes.scala 24:25]
  wire  monitor_1_io_in_flit_0_valid; // @[Nodes.scala 24:25]
  wire  monitor_1_io_in_flit_0_bits_head; // @[Nodes.scala 24:25]
  wire  monitor_1_io_in_flit_0_bits_tail; // @[Nodes.scala 24:25]
  wire [1:0] monitor_1_io_in_flit_0_bits_flow_ingress_node; // @[Nodes.scala 24:25]
  wire [1:0] monitor_1_io_in_flit_0_bits_flow_egress_node; // @[Nodes.scala 24:25]
  wire [1:0] monitor_1_io_in_flit_0_bits_virt_channel_id; // @[Nodes.scala 24:25]
  wire  input_unit_0_from_0_clock; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_reset; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_router_req_valid; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_0_io_router_req_bits_src_virt_id; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_0_io_router_req_bits_flow_ingress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_0_io_router_req_bits_flow_egress_node; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_router_resp_vc_sel_1_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_router_resp_vc_sel_1_1; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_router_resp_vc_sel_1_2; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_router_resp_vc_sel_1_3; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_router_resp_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_router_resp_vc_sel_0_1; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_router_resp_vc_sel_0_2; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_router_resp_vc_sel_0_3; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_req_ready; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_req_valid; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_2_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_1_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_1_1; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_1_2; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_1_3; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_1; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_2; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_3; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_resp_vc_sel_2_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_resp_vc_sel_1_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_resp_vc_sel_1_1; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_resp_vc_sel_1_2; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_resp_vc_sel_1_3; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_resp_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_resp_vc_sel_0_1; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_resp_vc_sel_0_2; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_resp_vc_sel_0_3; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_out_credit_available_2_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_out_credit_available_1_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_out_credit_available_1_1; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_out_credit_available_1_2; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_out_credit_available_1_3; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_out_credit_available_0_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_out_credit_available_0_1; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_out_credit_available_0_2; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_out_credit_available_0_3; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_salloc_req_0_ready; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_salloc_req_0_valid; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_2_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_1_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_1_1; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_1_2; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_1_3; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_1; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_2; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_3; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_salloc_req_0_bits_tail; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_out_0_valid; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_out_0_bits_flit_head; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_out_0_bits_flit_tail; // @[Router.scala 112:13]
  wire [63:0] input_unit_0_from_0_io_out_0_bits_flit_payload; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_0_io_out_0_bits_flit_flow_ingress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_0_io_out_0_bits_flit_flow_egress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_0_io_out_0_bits_out_virt_channel; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_0_io_debug_va_stall; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_0_io_debug_sa_stall; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_in_flit_0_valid; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_in_flit_0_bits_head; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_in_flit_0_bits_tail; // @[Router.scala 112:13]
  wire [63:0] input_unit_0_from_0_io_in_flit_0_bits_payload; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_0_io_in_flit_0_bits_flow_ingress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_0_io_in_flit_0_bits_flow_egress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_0_io_in_flit_0_bits_virt_channel_id; // @[Router.scala 112:13]
  wire [3:0] input_unit_0_from_0_io_in_credit_return; // @[Router.scala 112:13]
  wire [3:0] input_unit_0_from_0_io_in_vc_free; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_clock; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_reset; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_router_req_valid; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_2_io_router_req_bits_src_virt_id; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_2_io_router_req_bits_flow_ingress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_2_io_router_req_bits_flow_egress_node; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_router_resp_vc_sel_1_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_router_resp_vc_sel_1_1; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_router_resp_vc_sel_1_2; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_router_resp_vc_sel_1_3; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_router_resp_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_router_resp_vc_sel_0_1; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_router_resp_vc_sel_0_2; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_router_resp_vc_sel_0_3; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_req_ready; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_req_valid; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_2_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_1_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_1_1; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_1_2; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_1_3; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_0_1; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_0_2; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_0_3; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_resp_vc_sel_2_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_resp_vc_sel_1_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_resp_vc_sel_1_1; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_resp_vc_sel_1_2; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_resp_vc_sel_1_3; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_resp_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_resp_vc_sel_0_1; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_resp_vc_sel_0_2; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_resp_vc_sel_0_3; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_out_credit_available_2_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_out_credit_available_1_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_out_credit_available_1_1; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_out_credit_available_1_2; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_out_credit_available_1_3; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_out_credit_available_0_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_out_credit_available_0_1; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_out_credit_available_0_2; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_out_credit_available_0_3; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_salloc_req_0_ready; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_salloc_req_0_valid; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_2_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_1_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_1_1; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_1_2; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_1_3; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_0_1; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_0_2; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_0_3; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_salloc_req_0_bits_tail; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_out_0_valid; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_out_0_bits_flit_head; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_out_0_bits_flit_tail; // @[Router.scala 112:13]
  wire [63:0] input_unit_1_from_2_io_out_0_bits_flit_payload; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_2_io_out_0_bits_flit_flow_ingress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_2_io_out_0_bits_flit_flow_egress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_2_io_out_0_bits_out_virt_channel; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_2_io_debug_va_stall; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_2_io_debug_sa_stall; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_in_flit_0_valid; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_in_flit_0_bits_head; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_in_flit_0_bits_tail; // @[Router.scala 112:13]
  wire [63:0] input_unit_1_from_2_io_in_flit_0_bits_payload; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_2_io_in_flit_0_bits_flow_ingress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_2_io_in_flit_0_bits_flow_egress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_2_io_in_flit_0_bits_virt_channel_id; // @[Router.scala 112:13]
  wire [3:0] input_unit_1_from_2_io_in_credit_return; // @[Router.scala 112:13]
  wire [3:0] input_unit_1_from_2_io_in_vc_free; // @[Router.scala 112:13]
  wire  ingress_unit_2_from_1_clock; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_reset; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_router_req_valid; // @[Router.scala 116:13]
  wire [1:0] ingress_unit_2_from_1_io_router_req_bits_flow_ingress_node; // @[Router.scala 116:13]
  wire [1:0] ingress_unit_2_from_1_io_router_req_bits_flow_egress_node; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_router_resp_vc_sel_1_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_router_resp_vc_sel_1_1; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_router_resp_vc_sel_1_2; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_router_resp_vc_sel_1_3; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_router_resp_vc_sel_0_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_router_resp_vc_sel_0_1; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_router_resp_vc_sel_0_2; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_router_resp_vc_sel_0_3; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_vcalloc_req_ready; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_vcalloc_req_valid; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_vcalloc_req_bits_vc_sel_2_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_vcalloc_req_bits_vc_sel_1_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_vcalloc_req_bits_vc_sel_1_1; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_vcalloc_req_bits_vc_sel_1_2; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_vcalloc_req_bits_vc_sel_1_3; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_vcalloc_req_bits_vc_sel_0_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_vcalloc_req_bits_vc_sel_0_1; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_vcalloc_req_bits_vc_sel_0_2; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_vcalloc_req_bits_vc_sel_0_3; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_vcalloc_resp_vc_sel_2_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_vcalloc_resp_vc_sel_1_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_vcalloc_resp_vc_sel_1_1; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_vcalloc_resp_vc_sel_1_2; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_vcalloc_resp_vc_sel_1_3; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_vcalloc_resp_vc_sel_0_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_vcalloc_resp_vc_sel_0_1; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_vcalloc_resp_vc_sel_0_2; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_vcalloc_resp_vc_sel_0_3; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_out_credit_available_2_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_out_credit_available_1_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_out_credit_available_1_1; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_out_credit_available_1_2; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_out_credit_available_1_3; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_out_credit_available_0_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_out_credit_available_0_1; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_out_credit_available_0_2; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_out_credit_available_0_3; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_salloc_req_0_ready; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_salloc_req_0_valid; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_salloc_req_0_bits_vc_sel_2_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_salloc_req_0_bits_vc_sel_1_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_salloc_req_0_bits_vc_sel_1_1; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_salloc_req_0_bits_vc_sel_1_2; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_salloc_req_0_bits_vc_sel_1_3; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_salloc_req_0_bits_vc_sel_0_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_salloc_req_0_bits_vc_sel_0_1; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_salloc_req_0_bits_vc_sel_0_2; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_salloc_req_0_bits_vc_sel_0_3; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_salloc_req_0_bits_tail; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_out_0_valid; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_out_0_bits_flit_head; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_out_0_bits_flit_tail; // @[Router.scala 116:13]
  wire [63:0] ingress_unit_2_from_1_io_out_0_bits_flit_payload; // @[Router.scala 116:13]
  wire [1:0] ingress_unit_2_from_1_io_out_0_bits_flit_flow_ingress_node; // @[Router.scala 116:13]
  wire [1:0] ingress_unit_2_from_1_io_out_0_bits_flit_flow_egress_node; // @[Router.scala 116:13]
  wire [1:0] ingress_unit_2_from_1_io_out_0_bits_out_virt_channel; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_in_ready; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_in_valid; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_in_bits_head; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_1_io_in_bits_tail; // @[Router.scala 116:13]
  wire [63:0] ingress_unit_2_from_1_io_in_bits_payload; // @[Router.scala 116:13]
  wire [1:0] ingress_unit_2_from_1_io_in_bits_egress_id; // @[Router.scala 116:13]
  wire  output_unit_0_to_0_clock; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_reset; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_in_0_valid; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_in_0_bits_head; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_in_0_bits_tail; // @[Router.scala 122:13]
  wire [63:0] output_unit_0_to_0_io_in_0_bits_payload; // @[Router.scala 122:13]
  wire [1:0] output_unit_0_to_0_io_in_0_bits_flow_ingress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_0_to_0_io_in_0_bits_flow_egress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_0_to_0_io_in_0_bits_virt_channel_id; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_credit_available_0; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_credit_available_1; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_credit_available_2; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_credit_available_3; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_channel_status_0_occupied; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_channel_status_1_occupied; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_channel_status_2_occupied; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_channel_status_3_occupied; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_allocs_0_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_allocs_1_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_allocs_2_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_allocs_3_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_credit_alloc_0_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_credit_alloc_1_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_credit_alloc_2_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_credit_alloc_3_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_out_flit_0_valid; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_out_flit_0_bits_head; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_out_flit_0_bits_tail; // @[Router.scala 122:13]
  wire [63:0] output_unit_0_to_0_io_out_flit_0_bits_payload; // @[Router.scala 122:13]
  wire [1:0] output_unit_0_to_0_io_out_flit_0_bits_flow_ingress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_0_to_0_io_out_flit_0_bits_flow_egress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_0_to_0_io_out_flit_0_bits_virt_channel_id; // @[Router.scala 122:13]
  wire [3:0] output_unit_0_to_0_io_out_credit_return; // @[Router.scala 122:13]
  wire [3:0] output_unit_0_to_0_io_out_vc_free; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_clock; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_reset; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_in_0_valid; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_in_0_bits_head; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_in_0_bits_tail; // @[Router.scala 122:13]
  wire [63:0] output_unit_1_to_2_io_in_0_bits_payload; // @[Router.scala 122:13]
  wire [1:0] output_unit_1_to_2_io_in_0_bits_flow_ingress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_1_to_2_io_in_0_bits_flow_egress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_1_to_2_io_in_0_bits_virt_channel_id; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_credit_available_0; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_credit_available_1; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_credit_available_2; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_credit_available_3; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_channel_status_0_occupied; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_channel_status_1_occupied; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_channel_status_2_occupied; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_channel_status_3_occupied; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_allocs_0_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_allocs_1_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_allocs_2_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_allocs_3_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_credit_alloc_0_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_credit_alloc_1_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_credit_alloc_2_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_credit_alloc_3_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_out_flit_0_valid; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_out_flit_0_bits_head; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_out_flit_0_bits_tail; // @[Router.scala 122:13]
  wire [63:0] output_unit_1_to_2_io_out_flit_0_bits_payload; // @[Router.scala 122:13]
  wire [1:0] output_unit_1_to_2_io_out_flit_0_bits_flow_ingress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_1_to_2_io_out_flit_0_bits_flow_egress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_1_to_2_io_out_flit_0_bits_virt_channel_id; // @[Router.scala 122:13]
  wire [3:0] output_unit_1_to_2_io_out_credit_return; // @[Router.scala 122:13]
  wire [3:0] output_unit_1_to_2_io_out_vc_free; // @[Router.scala 122:13]
  wire  egress_unit_2_to_1_clock; // @[Router.scala 125:13]
  wire  egress_unit_2_to_1_reset; // @[Router.scala 125:13]
  wire  egress_unit_2_to_1_io_in_0_valid; // @[Router.scala 125:13]
  wire  egress_unit_2_to_1_io_in_0_bits_head; // @[Router.scala 125:13]
  wire  egress_unit_2_to_1_io_in_0_bits_tail; // @[Router.scala 125:13]
  wire [63:0] egress_unit_2_to_1_io_in_0_bits_payload; // @[Router.scala 125:13]
  wire [1:0] egress_unit_2_to_1_io_in_0_bits_flow_ingress_node; // @[Router.scala 125:13]
  wire  egress_unit_2_to_1_io_credit_available_0; // @[Router.scala 125:13]
  wire  egress_unit_2_to_1_io_channel_status_0_occupied; // @[Router.scala 125:13]
  wire  egress_unit_2_to_1_io_allocs_0_alloc; // @[Router.scala 125:13]
  wire  egress_unit_2_to_1_io_credit_alloc_0_alloc; // @[Router.scala 125:13]
  wire  egress_unit_2_to_1_io_credit_alloc_0_tail; // @[Router.scala 125:13]
  wire  egress_unit_2_to_1_io_out_valid; // @[Router.scala 125:13]
  wire  egress_unit_2_to_1_io_out_bits_head; // @[Router.scala 125:13]
  wire  egress_unit_2_to_1_io_out_bits_tail; // @[Router.scala 125:13]
  wire [63:0] egress_unit_2_to_1_io_out_bits_payload; // @[Router.scala 125:13]
  wire [1:0] egress_unit_2_to_1_io_out_bits_ingress_id; // @[Router.scala 125:13]
  wire  switch_clock; // @[Router.scala 129:24]
  wire  switch_reset; // @[Router.scala 129:24]
  wire  switch_io_in_2_0_valid; // @[Router.scala 129:24]
  wire  switch_io_in_2_0_bits_flit_head; // @[Router.scala 129:24]
  wire  switch_io_in_2_0_bits_flit_tail; // @[Router.scala 129:24]
  wire [63:0] switch_io_in_2_0_bits_flit_payload; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_2_0_bits_flit_flow_ingress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_2_0_bits_flit_flow_egress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_2_0_bits_out_virt_channel; // @[Router.scala 129:24]
  wire  switch_io_in_1_0_valid; // @[Router.scala 129:24]
  wire  switch_io_in_1_0_bits_flit_head; // @[Router.scala 129:24]
  wire  switch_io_in_1_0_bits_flit_tail; // @[Router.scala 129:24]
  wire [63:0] switch_io_in_1_0_bits_flit_payload; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_1_0_bits_flit_flow_ingress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_1_0_bits_flit_flow_egress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_1_0_bits_out_virt_channel; // @[Router.scala 129:24]
  wire  switch_io_in_0_0_valid; // @[Router.scala 129:24]
  wire  switch_io_in_0_0_bits_flit_head; // @[Router.scala 129:24]
  wire  switch_io_in_0_0_bits_flit_tail; // @[Router.scala 129:24]
  wire [63:0] switch_io_in_0_0_bits_flit_payload; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_0_0_bits_flit_flow_ingress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_0_0_bits_flit_flow_egress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_0_0_bits_out_virt_channel; // @[Router.scala 129:24]
  wire  switch_io_out_2_0_valid; // @[Router.scala 129:24]
  wire  switch_io_out_2_0_bits_head; // @[Router.scala 129:24]
  wire  switch_io_out_2_0_bits_tail; // @[Router.scala 129:24]
  wire [63:0] switch_io_out_2_0_bits_payload; // @[Router.scala 129:24]
  wire [1:0] switch_io_out_2_0_bits_flow_ingress_node; // @[Router.scala 129:24]
  wire  switch_io_out_1_0_valid; // @[Router.scala 129:24]
  wire  switch_io_out_1_0_bits_head; // @[Router.scala 129:24]
  wire  switch_io_out_1_0_bits_tail; // @[Router.scala 129:24]
  wire [63:0] switch_io_out_1_0_bits_payload; // @[Router.scala 129:24]
  wire [1:0] switch_io_out_1_0_bits_flow_ingress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_out_1_0_bits_flow_egress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_out_1_0_bits_virt_channel_id; // @[Router.scala 129:24]
  wire  switch_io_out_0_0_valid; // @[Router.scala 129:24]
  wire  switch_io_out_0_0_bits_head; // @[Router.scala 129:24]
  wire  switch_io_out_0_0_bits_tail; // @[Router.scala 129:24]
  wire [63:0] switch_io_out_0_0_bits_payload; // @[Router.scala 129:24]
  wire [1:0] switch_io_out_0_0_bits_flow_ingress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_out_0_0_bits_flow_egress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_out_0_0_bits_virt_channel_id; // @[Router.scala 129:24]
  wire  switch_io_sel_2_0_2_0; // @[Router.scala 129:24]
  wire  switch_io_sel_2_0_1_0; // @[Router.scala 129:24]
  wire  switch_io_sel_2_0_0_0; // @[Router.scala 129:24]
  wire  switch_io_sel_1_0_2_0; // @[Router.scala 129:24]
  wire  switch_io_sel_1_0_1_0; // @[Router.scala 129:24]
  wire  switch_io_sel_1_0_0_0; // @[Router.scala 129:24]
  wire  switch_io_sel_0_0_2_0; // @[Router.scala 129:24]
  wire  switch_io_sel_0_0_1_0; // @[Router.scala 129:24]
  wire  switch_io_sel_0_0_0_0; // @[Router.scala 129:24]
  wire  switch_allocator_clock; // @[Router.scala 130:34]
  wire  switch_allocator_reset; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_ready; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_valid; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_bits_vc_sel_2_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_bits_vc_sel_1_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_bits_vc_sel_1_1; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_bits_vc_sel_1_2; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_bits_vc_sel_1_3; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_bits_vc_sel_0_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_bits_vc_sel_0_1; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_bits_vc_sel_0_2; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_bits_vc_sel_0_3; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_bits_tail; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_ready; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_valid; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_vc_sel_2_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_vc_sel_1_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_vc_sel_1_1; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_vc_sel_1_2; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_vc_sel_1_3; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_vc_sel_0_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_vc_sel_0_1; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_vc_sel_0_2; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_vc_sel_0_3; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_tail; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_ready; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_valid; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_2_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_1_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_1_1; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_1_2; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_1_3; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_0_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_0_1; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_0_2; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_0_3; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_tail; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_2_0_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_2_0_tail; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_1_0_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_1_1_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_1_2_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_1_3_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_0_0_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_0_1_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_0_2_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_0_3_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_2_0_2_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_2_0_1_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_2_0_0_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_1_0_2_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_1_0_1_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_1_0_0_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_0_0_2_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_0_0_1_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_0_0_0_0; // @[Router.scala 130:34]
  wire  vc_allocator_clock; // @[Router.scala 131:30]
  wire  vc_allocator_reset; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_ready; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_valid; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_bits_vc_sel_2_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_bits_vc_sel_1_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_bits_vc_sel_1_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_bits_vc_sel_1_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_bits_vc_sel_1_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_bits_vc_sel_0_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_bits_vc_sel_0_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_bits_vc_sel_0_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_bits_vc_sel_0_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_ready; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_valid; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_bits_vc_sel_2_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_bits_vc_sel_1_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_bits_vc_sel_1_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_bits_vc_sel_1_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_bits_vc_sel_1_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_bits_vc_sel_0_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_bits_vc_sel_0_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_bits_vc_sel_0_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_bits_vc_sel_0_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_ready; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_valid; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_2_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_1_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_1_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_1_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_1_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_0_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_0_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_0_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_0_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_2_vc_sel_2_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_2_vc_sel_1_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_2_vc_sel_1_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_2_vc_sel_1_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_2_vc_sel_1_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_2_vc_sel_0_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_2_vc_sel_0_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_2_vc_sel_0_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_2_vc_sel_0_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_1_vc_sel_2_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_1_vc_sel_1_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_1_vc_sel_1_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_1_vc_sel_1_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_1_vc_sel_1_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_1_vc_sel_0_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_1_vc_sel_0_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_1_vc_sel_0_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_1_vc_sel_0_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_2_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_1_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_1_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_1_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_1_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_0_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_0_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_0_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_0_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_2_0_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_1_0_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_1_1_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_1_2_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_1_3_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_0_0_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_0_1_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_0_2_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_0_3_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_2_0_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_1_0_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_1_1_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_1_2_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_1_3_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_0_0_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_0_1_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_0_2_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_0_3_alloc; // @[Router.scala 131:30]
  wire [1:0] route_computer_io_req_2_bits_flow_ingress_node; // @[Router.scala 134:32]
  wire [1:0] route_computer_io_req_2_bits_flow_egress_node; // @[Router.scala 134:32]
  wire [1:0] route_computer_io_req_1_bits_src_virt_id; // @[Router.scala 134:32]
  wire [1:0] route_computer_io_req_1_bits_flow_ingress_node; // @[Router.scala 134:32]
  wire [1:0] route_computer_io_req_1_bits_flow_egress_node; // @[Router.scala 134:32]
  wire [1:0] route_computer_io_req_0_bits_src_virt_id; // @[Router.scala 134:32]
  wire [1:0] route_computer_io_req_0_bits_flow_ingress_node; // @[Router.scala 134:32]
  wire [1:0] route_computer_io_req_0_bits_flow_egress_node; // @[Router.scala 134:32]
  wire  route_computer_io_resp_2_vc_sel_1_0; // @[Router.scala 134:32]
  wire  route_computer_io_resp_2_vc_sel_1_1; // @[Router.scala 134:32]
  wire  route_computer_io_resp_2_vc_sel_1_2; // @[Router.scala 134:32]
  wire  route_computer_io_resp_2_vc_sel_1_3; // @[Router.scala 134:32]
  wire  route_computer_io_resp_2_vc_sel_0_0; // @[Router.scala 134:32]
  wire  route_computer_io_resp_2_vc_sel_0_1; // @[Router.scala 134:32]
  wire  route_computer_io_resp_2_vc_sel_0_2; // @[Router.scala 134:32]
  wire  route_computer_io_resp_2_vc_sel_0_3; // @[Router.scala 134:32]
  wire  route_computer_io_resp_1_vc_sel_1_0; // @[Router.scala 134:32]
  wire  route_computer_io_resp_1_vc_sel_1_1; // @[Router.scala 134:32]
  wire  route_computer_io_resp_1_vc_sel_1_2; // @[Router.scala 134:32]
  wire  route_computer_io_resp_1_vc_sel_1_3; // @[Router.scala 134:32]
  wire  route_computer_io_resp_1_vc_sel_0_0; // @[Router.scala 134:32]
  wire  route_computer_io_resp_1_vc_sel_0_1; // @[Router.scala 134:32]
  wire  route_computer_io_resp_1_vc_sel_0_2; // @[Router.scala 134:32]
  wire  route_computer_io_resp_1_vc_sel_0_3; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_1_0; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_1_1; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_1_2; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_1_3; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_0_0; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_0_1; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_0_2; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_0_3; // @[Router.scala 134:32]
  wire [19:0] plusarg_reader_out; // @[PlusArg.scala 80:11]
  wire  _fires_count_T = vc_allocator_io_req_0_ready & vc_allocator_io_req_0_valid; // @[Decoupled.scala 51:35]
  wire  _fires_count_T_1 = vc_allocator_io_req_1_ready & vc_allocator_io_req_1_valid; // @[Decoupled.scala 51:35]
  wire  _fires_count_T_2 = vc_allocator_io_req_2_ready & vc_allocator_io_req_2_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _fires_count_T_3 = _fires_count_T_1 + _fires_count_T_2; // @[Bitwise.scala 51:90]
  wire [1:0] _GEN_5 = {{1'd0}, _fires_count_T}; // @[Bitwise.scala 51:90]
  wire [2:0] _fires_count_T_5 = _GEN_5 + _fires_count_T_3; // @[Bitwise.scala 51:90]
  reg  switch_io_sel_REG_2_0_2_0; // @[Router.scala 176:14]
  reg  switch_io_sel_REG_2_0_1_0; // @[Router.scala 176:14]
  reg  switch_io_sel_REG_2_0_0_0; // @[Router.scala 176:14]
  reg  switch_io_sel_REG_1_0_2_0; // @[Router.scala 176:14]
  reg  switch_io_sel_REG_1_0_1_0; // @[Router.scala 176:14]
  reg  switch_io_sel_REG_1_0_0_0; // @[Router.scala 176:14]
  reg  switch_io_sel_REG_0_0_2_0; // @[Router.scala 176:14]
  reg  switch_io_sel_REG_0_0_1_0; // @[Router.scala 176:14]
  reg  switch_io_sel_REG_0_0_0_0; // @[Router.scala 176:14]
  reg [63:0] debug_tsc; // @[Router.scala 193:28]
  wire [63:0] _debug_tsc_T_1 = debug_tsc + 64'h1; // @[Router.scala 194:28]
  reg [63:0] debug_sample; // @[Router.scala 195:31]
  wire [63:0] _debug_sample_T_1 = debug_sample + 64'h1; // @[Router.scala 196:34]
  wire [19:0] _T_1 = plusarg_reader_out - 20'h1; // @[Router.scala 198:40]
  wire [63:0] _GEN_6 = {{44'd0}, _T_1}; // @[Router.scala 198:24]
  wire  _T_2 = debug_sample == _GEN_6; // @[Router.scala 198:24]
  reg [63:0] util_ctr; // @[Router.scala 201:29]
  reg  fired; // @[Router.scala 202:26]
  wire [63:0] _GEN_7 = {{63'd0}, auto_dest_nodes_in_0_flit_0_valid}; // @[Router.scala 203:28]
  wire [63:0] _util_ctr_T_1 = util_ctr + _GEN_7; // @[Router.scala 203:28]
  wire  _T_8 = plusarg_reader_out != 20'h0 & _T_2 & fired; // @[Router.scala 205:71]
  reg [63:0] util_ctr_1; // @[Router.scala 201:29]
  reg  fired_1; // @[Router.scala 202:26]
  wire [63:0] _GEN_9 = {{63'd0}, auto_dest_nodes_in_1_flit_0_valid}; // @[Router.scala 203:28]
  wire [63:0] _util_ctr_T_3 = util_ctr_1 + _GEN_9; // @[Router.scala 203:28]
  wire  _T_16 = plusarg_reader_out != 20'h0 & _T_2 & fired_1; // @[Router.scala 205:71]
  wire  bundleIn_0_2_flit_ready = ingress_unit_2_from_1_io_in_ready; // @[Nodes.scala 1215:84 Router.scala 142:68]
  wire  _T_19 = bundleIn_0_2_flit_ready & auto_ingress_nodes_in_flit_valid; // @[Decoupled.scala 51:35]
  reg [63:0] util_ctr_2; // @[Router.scala 201:29]
  reg  fired_2; // @[Router.scala 202:26]
  wire [63:0] _GEN_11 = {{63'd0}, _T_19}; // @[Router.scala 203:28]
  wire [63:0] _util_ctr_T_5 = util_ctr_2 + _GEN_11; // @[Router.scala 203:28]
  wire  _T_25 = plusarg_reader_out != 20'h0 & _T_2 & fired_2; // @[Router.scala 205:71]
  wire  x1_2_flit_valid = egress_unit_2_to_1_io_out_valid; // @[Nodes.scala 1212:84 Router.scala 144:65]
  reg [63:0] util_ctr_3; // @[Router.scala 201:29]
  reg  fired_3; // @[Router.scala 202:26]
  wire [63:0] _GEN_13 = {{63'd0}, x1_2_flit_valid}; // @[Router.scala 203:28]
  wire [63:0] _util_ctr_T_7 = util_ctr_3 + _GEN_13; // @[Router.scala 203:28]
  wire  _T_34 = plusarg_reader_out != 20'h0 & _T_2 & fired_3; // @[Router.scala 205:71]
  wire [1:0] fires_count = _fires_count_T_5[1:0]; // @[Bitwise.scala 51:90]
  NoCMonitor_2 monitor ( // @[Nodes.scala 24:25]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_flit_0_valid(monitor_io_in_flit_0_valid),
    .io_in_flit_0_bits_head(monitor_io_in_flit_0_bits_head),
    .io_in_flit_0_bits_tail(monitor_io_in_flit_0_bits_tail),
    .io_in_flit_0_bits_flow_ingress_node(monitor_io_in_flit_0_bits_flow_ingress_node),
    .io_in_flit_0_bits_flow_egress_node(monitor_io_in_flit_0_bits_flow_egress_node),
    .io_in_flit_0_bits_virt_channel_id(monitor_io_in_flit_0_bits_virt_channel_id)
  );
  NoCMonitor_3 monitor_1 ( // @[Nodes.scala 24:25]
    .clock(monitor_1_clock),
    .reset(monitor_1_reset),
    .io_in_flit_0_valid(monitor_1_io_in_flit_0_valid),
    .io_in_flit_0_bits_head(monitor_1_io_in_flit_0_bits_head),
    .io_in_flit_0_bits_tail(monitor_1_io_in_flit_0_bits_tail),
    .io_in_flit_0_bits_flow_ingress_node(monitor_1_io_in_flit_0_bits_flow_ingress_node),
    .io_in_flit_0_bits_flow_egress_node(monitor_1_io_in_flit_0_bits_flow_egress_node),
    .io_in_flit_0_bits_virt_channel_id(monitor_1_io_in_flit_0_bits_virt_channel_id)
  );
  InputUnit_2 input_unit_0_from_0 ( // @[Router.scala 112:13]
    .clock(input_unit_0_from_0_clock),
    .reset(input_unit_0_from_0_reset),
    .io_router_req_valid(input_unit_0_from_0_io_router_req_valid),
    .io_router_req_bits_src_virt_id(input_unit_0_from_0_io_router_req_bits_src_virt_id),
    .io_router_req_bits_flow_ingress_node(input_unit_0_from_0_io_router_req_bits_flow_ingress_node),
    .io_router_req_bits_flow_egress_node(input_unit_0_from_0_io_router_req_bits_flow_egress_node),
    .io_router_resp_vc_sel_1_0(input_unit_0_from_0_io_router_resp_vc_sel_1_0),
    .io_router_resp_vc_sel_1_1(input_unit_0_from_0_io_router_resp_vc_sel_1_1),
    .io_router_resp_vc_sel_1_2(input_unit_0_from_0_io_router_resp_vc_sel_1_2),
    .io_router_resp_vc_sel_1_3(input_unit_0_from_0_io_router_resp_vc_sel_1_3),
    .io_router_resp_vc_sel_0_0(input_unit_0_from_0_io_router_resp_vc_sel_0_0),
    .io_router_resp_vc_sel_0_1(input_unit_0_from_0_io_router_resp_vc_sel_0_1),
    .io_router_resp_vc_sel_0_2(input_unit_0_from_0_io_router_resp_vc_sel_0_2),
    .io_router_resp_vc_sel_0_3(input_unit_0_from_0_io_router_resp_vc_sel_0_3),
    .io_vcalloc_req_ready(input_unit_0_from_0_io_vcalloc_req_ready),
    .io_vcalloc_req_valid(input_unit_0_from_0_io_vcalloc_req_valid),
    .io_vcalloc_req_bits_vc_sel_2_0(input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_2_0),
    .io_vcalloc_req_bits_vc_sel_1_0(input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_1_0),
    .io_vcalloc_req_bits_vc_sel_1_1(input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_1_1),
    .io_vcalloc_req_bits_vc_sel_1_2(input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_1_2),
    .io_vcalloc_req_bits_vc_sel_1_3(input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_1_3),
    .io_vcalloc_req_bits_vc_sel_0_0(input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_0),
    .io_vcalloc_req_bits_vc_sel_0_1(input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_1),
    .io_vcalloc_req_bits_vc_sel_0_2(input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_2),
    .io_vcalloc_req_bits_vc_sel_0_3(input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_3),
    .io_vcalloc_resp_vc_sel_2_0(input_unit_0_from_0_io_vcalloc_resp_vc_sel_2_0),
    .io_vcalloc_resp_vc_sel_1_0(input_unit_0_from_0_io_vcalloc_resp_vc_sel_1_0),
    .io_vcalloc_resp_vc_sel_1_1(input_unit_0_from_0_io_vcalloc_resp_vc_sel_1_1),
    .io_vcalloc_resp_vc_sel_1_2(input_unit_0_from_0_io_vcalloc_resp_vc_sel_1_2),
    .io_vcalloc_resp_vc_sel_1_3(input_unit_0_from_0_io_vcalloc_resp_vc_sel_1_3),
    .io_vcalloc_resp_vc_sel_0_0(input_unit_0_from_0_io_vcalloc_resp_vc_sel_0_0),
    .io_vcalloc_resp_vc_sel_0_1(input_unit_0_from_0_io_vcalloc_resp_vc_sel_0_1),
    .io_vcalloc_resp_vc_sel_0_2(input_unit_0_from_0_io_vcalloc_resp_vc_sel_0_2),
    .io_vcalloc_resp_vc_sel_0_3(input_unit_0_from_0_io_vcalloc_resp_vc_sel_0_3),
    .io_out_credit_available_2_0(input_unit_0_from_0_io_out_credit_available_2_0),
    .io_out_credit_available_1_0(input_unit_0_from_0_io_out_credit_available_1_0),
    .io_out_credit_available_1_1(input_unit_0_from_0_io_out_credit_available_1_1),
    .io_out_credit_available_1_2(input_unit_0_from_0_io_out_credit_available_1_2),
    .io_out_credit_available_1_3(input_unit_0_from_0_io_out_credit_available_1_3),
    .io_out_credit_available_0_0(input_unit_0_from_0_io_out_credit_available_0_0),
    .io_out_credit_available_0_1(input_unit_0_from_0_io_out_credit_available_0_1),
    .io_out_credit_available_0_2(input_unit_0_from_0_io_out_credit_available_0_2),
    .io_out_credit_available_0_3(input_unit_0_from_0_io_out_credit_available_0_3),
    .io_salloc_req_0_ready(input_unit_0_from_0_io_salloc_req_0_ready),
    .io_salloc_req_0_valid(input_unit_0_from_0_io_salloc_req_0_valid),
    .io_salloc_req_0_bits_vc_sel_2_0(input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_2_0),
    .io_salloc_req_0_bits_vc_sel_1_0(input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_1_0),
    .io_salloc_req_0_bits_vc_sel_1_1(input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_1_1),
    .io_salloc_req_0_bits_vc_sel_1_2(input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_1_2),
    .io_salloc_req_0_bits_vc_sel_1_3(input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_1_3),
    .io_salloc_req_0_bits_vc_sel_0_0(input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_0),
    .io_salloc_req_0_bits_vc_sel_0_1(input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_1),
    .io_salloc_req_0_bits_vc_sel_0_2(input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_2),
    .io_salloc_req_0_bits_vc_sel_0_3(input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_3),
    .io_salloc_req_0_bits_tail(input_unit_0_from_0_io_salloc_req_0_bits_tail),
    .io_out_0_valid(input_unit_0_from_0_io_out_0_valid),
    .io_out_0_bits_flit_head(input_unit_0_from_0_io_out_0_bits_flit_head),
    .io_out_0_bits_flit_tail(input_unit_0_from_0_io_out_0_bits_flit_tail),
    .io_out_0_bits_flit_payload(input_unit_0_from_0_io_out_0_bits_flit_payload),
    .io_out_0_bits_flit_flow_ingress_node(input_unit_0_from_0_io_out_0_bits_flit_flow_ingress_node),
    .io_out_0_bits_flit_flow_egress_node(input_unit_0_from_0_io_out_0_bits_flit_flow_egress_node),
    .io_out_0_bits_out_virt_channel(input_unit_0_from_0_io_out_0_bits_out_virt_channel),
    .io_debug_va_stall(input_unit_0_from_0_io_debug_va_stall),
    .io_debug_sa_stall(input_unit_0_from_0_io_debug_sa_stall),
    .io_in_flit_0_valid(input_unit_0_from_0_io_in_flit_0_valid),
    .io_in_flit_0_bits_head(input_unit_0_from_0_io_in_flit_0_bits_head),
    .io_in_flit_0_bits_tail(input_unit_0_from_0_io_in_flit_0_bits_tail),
    .io_in_flit_0_bits_payload(input_unit_0_from_0_io_in_flit_0_bits_payload),
    .io_in_flit_0_bits_flow_ingress_node(input_unit_0_from_0_io_in_flit_0_bits_flow_ingress_node),
    .io_in_flit_0_bits_flow_egress_node(input_unit_0_from_0_io_in_flit_0_bits_flow_egress_node),
    .io_in_flit_0_bits_virt_channel_id(input_unit_0_from_0_io_in_flit_0_bits_virt_channel_id),
    .io_in_credit_return(input_unit_0_from_0_io_in_credit_return),
    .io_in_vc_free(input_unit_0_from_0_io_in_vc_free)
  );
  InputUnit_3 input_unit_1_from_2 ( // @[Router.scala 112:13]
    .clock(input_unit_1_from_2_clock),
    .reset(input_unit_1_from_2_reset),
    .io_router_req_valid(input_unit_1_from_2_io_router_req_valid),
    .io_router_req_bits_src_virt_id(input_unit_1_from_2_io_router_req_bits_src_virt_id),
    .io_router_req_bits_flow_ingress_node(input_unit_1_from_2_io_router_req_bits_flow_ingress_node),
    .io_router_req_bits_flow_egress_node(input_unit_1_from_2_io_router_req_bits_flow_egress_node),
    .io_router_resp_vc_sel_1_0(input_unit_1_from_2_io_router_resp_vc_sel_1_0),
    .io_router_resp_vc_sel_1_1(input_unit_1_from_2_io_router_resp_vc_sel_1_1),
    .io_router_resp_vc_sel_1_2(input_unit_1_from_2_io_router_resp_vc_sel_1_2),
    .io_router_resp_vc_sel_1_3(input_unit_1_from_2_io_router_resp_vc_sel_1_3),
    .io_router_resp_vc_sel_0_0(input_unit_1_from_2_io_router_resp_vc_sel_0_0),
    .io_router_resp_vc_sel_0_1(input_unit_1_from_2_io_router_resp_vc_sel_0_1),
    .io_router_resp_vc_sel_0_2(input_unit_1_from_2_io_router_resp_vc_sel_0_2),
    .io_router_resp_vc_sel_0_3(input_unit_1_from_2_io_router_resp_vc_sel_0_3),
    .io_vcalloc_req_ready(input_unit_1_from_2_io_vcalloc_req_ready),
    .io_vcalloc_req_valid(input_unit_1_from_2_io_vcalloc_req_valid),
    .io_vcalloc_req_bits_vc_sel_2_0(input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_2_0),
    .io_vcalloc_req_bits_vc_sel_1_0(input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_1_0),
    .io_vcalloc_req_bits_vc_sel_1_1(input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_1_1),
    .io_vcalloc_req_bits_vc_sel_1_2(input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_1_2),
    .io_vcalloc_req_bits_vc_sel_1_3(input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_1_3),
    .io_vcalloc_req_bits_vc_sel_0_0(input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_0_0),
    .io_vcalloc_req_bits_vc_sel_0_1(input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_0_1),
    .io_vcalloc_req_bits_vc_sel_0_2(input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_0_2),
    .io_vcalloc_req_bits_vc_sel_0_3(input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_0_3),
    .io_vcalloc_resp_vc_sel_2_0(input_unit_1_from_2_io_vcalloc_resp_vc_sel_2_0),
    .io_vcalloc_resp_vc_sel_1_0(input_unit_1_from_2_io_vcalloc_resp_vc_sel_1_0),
    .io_vcalloc_resp_vc_sel_1_1(input_unit_1_from_2_io_vcalloc_resp_vc_sel_1_1),
    .io_vcalloc_resp_vc_sel_1_2(input_unit_1_from_2_io_vcalloc_resp_vc_sel_1_2),
    .io_vcalloc_resp_vc_sel_1_3(input_unit_1_from_2_io_vcalloc_resp_vc_sel_1_3),
    .io_vcalloc_resp_vc_sel_0_0(input_unit_1_from_2_io_vcalloc_resp_vc_sel_0_0),
    .io_vcalloc_resp_vc_sel_0_1(input_unit_1_from_2_io_vcalloc_resp_vc_sel_0_1),
    .io_vcalloc_resp_vc_sel_0_2(input_unit_1_from_2_io_vcalloc_resp_vc_sel_0_2),
    .io_vcalloc_resp_vc_sel_0_3(input_unit_1_from_2_io_vcalloc_resp_vc_sel_0_3),
    .io_out_credit_available_2_0(input_unit_1_from_2_io_out_credit_available_2_0),
    .io_out_credit_available_1_0(input_unit_1_from_2_io_out_credit_available_1_0),
    .io_out_credit_available_1_1(input_unit_1_from_2_io_out_credit_available_1_1),
    .io_out_credit_available_1_2(input_unit_1_from_2_io_out_credit_available_1_2),
    .io_out_credit_available_1_3(input_unit_1_from_2_io_out_credit_available_1_3),
    .io_out_credit_available_0_0(input_unit_1_from_2_io_out_credit_available_0_0),
    .io_out_credit_available_0_1(input_unit_1_from_2_io_out_credit_available_0_1),
    .io_out_credit_available_0_2(input_unit_1_from_2_io_out_credit_available_0_2),
    .io_out_credit_available_0_3(input_unit_1_from_2_io_out_credit_available_0_3),
    .io_salloc_req_0_ready(input_unit_1_from_2_io_salloc_req_0_ready),
    .io_salloc_req_0_valid(input_unit_1_from_2_io_salloc_req_0_valid),
    .io_salloc_req_0_bits_vc_sel_2_0(input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_2_0),
    .io_salloc_req_0_bits_vc_sel_1_0(input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_1_0),
    .io_salloc_req_0_bits_vc_sel_1_1(input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_1_1),
    .io_salloc_req_0_bits_vc_sel_1_2(input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_1_2),
    .io_salloc_req_0_bits_vc_sel_1_3(input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_1_3),
    .io_salloc_req_0_bits_vc_sel_0_0(input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_0_0),
    .io_salloc_req_0_bits_vc_sel_0_1(input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_0_1),
    .io_salloc_req_0_bits_vc_sel_0_2(input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_0_2),
    .io_salloc_req_0_bits_vc_sel_0_3(input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_0_3),
    .io_salloc_req_0_bits_tail(input_unit_1_from_2_io_salloc_req_0_bits_tail),
    .io_out_0_valid(input_unit_1_from_2_io_out_0_valid),
    .io_out_0_bits_flit_head(input_unit_1_from_2_io_out_0_bits_flit_head),
    .io_out_0_bits_flit_tail(input_unit_1_from_2_io_out_0_bits_flit_tail),
    .io_out_0_bits_flit_payload(input_unit_1_from_2_io_out_0_bits_flit_payload),
    .io_out_0_bits_flit_flow_ingress_node(input_unit_1_from_2_io_out_0_bits_flit_flow_ingress_node),
    .io_out_0_bits_flit_flow_egress_node(input_unit_1_from_2_io_out_0_bits_flit_flow_egress_node),
    .io_out_0_bits_out_virt_channel(input_unit_1_from_2_io_out_0_bits_out_virt_channel),
    .io_debug_va_stall(input_unit_1_from_2_io_debug_va_stall),
    .io_debug_sa_stall(input_unit_1_from_2_io_debug_sa_stall),
    .io_in_flit_0_valid(input_unit_1_from_2_io_in_flit_0_valid),
    .io_in_flit_0_bits_head(input_unit_1_from_2_io_in_flit_0_bits_head),
    .io_in_flit_0_bits_tail(input_unit_1_from_2_io_in_flit_0_bits_tail),
    .io_in_flit_0_bits_payload(input_unit_1_from_2_io_in_flit_0_bits_payload),
    .io_in_flit_0_bits_flow_ingress_node(input_unit_1_from_2_io_in_flit_0_bits_flow_ingress_node),
    .io_in_flit_0_bits_flow_egress_node(input_unit_1_from_2_io_in_flit_0_bits_flow_egress_node),
    .io_in_flit_0_bits_virt_channel_id(input_unit_1_from_2_io_in_flit_0_bits_virt_channel_id),
    .io_in_credit_return(input_unit_1_from_2_io_in_credit_return),
    .io_in_vc_free(input_unit_1_from_2_io_in_vc_free)
  );
  IngressUnit_1 ingress_unit_2_from_1 ( // @[Router.scala 116:13]
    .clock(ingress_unit_2_from_1_clock),
    .reset(ingress_unit_2_from_1_reset),
    .io_router_req_valid(ingress_unit_2_from_1_io_router_req_valid),
    .io_router_req_bits_flow_ingress_node(ingress_unit_2_from_1_io_router_req_bits_flow_ingress_node),
    .io_router_req_bits_flow_egress_node(ingress_unit_2_from_1_io_router_req_bits_flow_egress_node),
    .io_router_resp_vc_sel_1_0(ingress_unit_2_from_1_io_router_resp_vc_sel_1_0),
    .io_router_resp_vc_sel_1_1(ingress_unit_2_from_1_io_router_resp_vc_sel_1_1),
    .io_router_resp_vc_sel_1_2(ingress_unit_2_from_1_io_router_resp_vc_sel_1_2),
    .io_router_resp_vc_sel_1_3(ingress_unit_2_from_1_io_router_resp_vc_sel_1_3),
    .io_router_resp_vc_sel_0_0(ingress_unit_2_from_1_io_router_resp_vc_sel_0_0),
    .io_router_resp_vc_sel_0_1(ingress_unit_2_from_1_io_router_resp_vc_sel_0_1),
    .io_router_resp_vc_sel_0_2(ingress_unit_2_from_1_io_router_resp_vc_sel_0_2),
    .io_router_resp_vc_sel_0_3(ingress_unit_2_from_1_io_router_resp_vc_sel_0_3),
    .io_vcalloc_req_ready(ingress_unit_2_from_1_io_vcalloc_req_ready),
    .io_vcalloc_req_valid(ingress_unit_2_from_1_io_vcalloc_req_valid),
    .io_vcalloc_req_bits_vc_sel_2_0(ingress_unit_2_from_1_io_vcalloc_req_bits_vc_sel_2_0),
    .io_vcalloc_req_bits_vc_sel_1_0(ingress_unit_2_from_1_io_vcalloc_req_bits_vc_sel_1_0),
    .io_vcalloc_req_bits_vc_sel_1_1(ingress_unit_2_from_1_io_vcalloc_req_bits_vc_sel_1_1),
    .io_vcalloc_req_bits_vc_sel_1_2(ingress_unit_2_from_1_io_vcalloc_req_bits_vc_sel_1_2),
    .io_vcalloc_req_bits_vc_sel_1_3(ingress_unit_2_from_1_io_vcalloc_req_bits_vc_sel_1_3),
    .io_vcalloc_req_bits_vc_sel_0_0(ingress_unit_2_from_1_io_vcalloc_req_bits_vc_sel_0_0),
    .io_vcalloc_req_bits_vc_sel_0_1(ingress_unit_2_from_1_io_vcalloc_req_bits_vc_sel_0_1),
    .io_vcalloc_req_bits_vc_sel_0_2(ingress_unit_2_from_1_io_vcalloc_req_bits_vc_sel_0_2),
    .io_vcalloc_req_bits_vc_sel_0_3(ingress_unit_2_from_1_io_vcalloc_req_bits_vc_sel_0_3),
    .io_vcalloc_resp_vc_sel_2_0(ingress_unit_2_from_1_io_vcalloc_resp_vc_sel_2_0),
    .io_vcalloc_resp_vc_sel_1_0(ingress_unit_2_from_1_io_vcalloc_resp_vc_sel_1_0),
    .io_vcalloc_resp_vc_sel_1_1(ingress_unit_2_from_1_io_vcalloc_resp_vc_sel_1_1),
    .io_vcalloc_resp_vc_sel_1_2(ingress_unit_2_from_1_io_vcalloc_resp_vc_sel_1_2),
    .io_vcalloc_resp_vc_sel_1_3(ingress_unit_2_from_1_io_vcalloc_resp_vc_sel_1_3),
    .io_vcalloc_resp_vc_sel_0_0(ingress_unit_2_from_1_io_vcalloc_resp_vc_sel_0_0),
    .io_vcalloc_resp_vc_sel_0_1(ingress_unit_2_from_1_io_vcalloc_resp_vc_sel_0_1),
    .io_vcalloc_resp_vc_sel_0_2(ingress_unit_2_from_1_io_vcalloc_resp_vc_sel_0_2),
    .io_vcalloc_resp_vc_sel_0_3(ingress_unit_2_from_1_io_vcalloc_resp_vc_sel_0_3),
    .io_out_credit_available_2_0(ingress_unit_2_from_1_io_out_credit_available_2_0),
    .io_out_credit_available_1_0(ingress_unit_2_from_1_io_out_credit_available_1_0),
    .io_out_credit_available_1_1(ingress_unit_2_from_1_io_out_credit_available_1_1),
    .io_out_credit_available_1_2(ingress_unit_2_from_1_io_out_credit_available_1_2),
    .io_out_credit_available_1_3(ingress_unit_2_from_1_io_out_credit_available_1_3),
    .io_out_credit_available_0_0(ingress_unit_2_from_1_io_out_credit_available_0_0),
    .io_out_credit_available_0_1(ingress_unit_2_from_1_io_out_credit_available_0_1),
    .io_out_credit_available_0_2(ingress_unit_2_from_1_io_out_credit_available_0_2),
    .io_out_credit_available_0_3(ingress_unit_2_from_1_io_out_credit_available_0_3),
    .io_salloc_req_0_ready(ingress_unit_2_from_1_io_salloc_req_0_ready),
    .io_salloc_req_0_valid(ingress_unit_2_from_1_io_salloc_req_0_valid),
    .io_salloc_req_0_bits_vc_sel_2_0(ingress_unit_2_from_1_io_salloc_req_0_bits_vc_sel_2_0),
    .io_salloc_req_0_bits_vc_sel_1_0(ingress_unit_2_from_1_io_salloc_req_0_bits_vc_sel_1_0),
    .io_salloc_req_0_bits_vc_sel_1_1(ingress_unit_2_from_1_io_salloc_req_0_bits_vc_sel_1_1),
    .io_salloc_req_0_bits_vc_sel_1_2(ingress_unit_2_from_1_io_salloc_req_0_bits_vc_sel_1_2),
    .io_salloc_req_0_bits_vc_sel_1_3(ingress_unit_2_from_1_io_salloc_req_0_bits_vc_sel_1_3),
    .io_salloc_req_0_bits_vc_sel_0_0(ingress_unit_2_from_1_io_salloc_req_0_bits_vc_sel_0_0),
    .io_salloc_req_0_bits_vc_sel_0_1(ingress_unit_2_from_1_io_salloc_req_0_bits_vc_sel_0_1),
    .io_salloc_req_0_bits_vc_sel_0_2(ingress_unit_2_from_1_io_salloc_req_0_bits_vc_sel_0_2),
    .io_salloc_req_0_bits_vc_sel_0_3(ingress_unit_2_from_1_io_salloc_req_0_bits_vc_sel_0_3),
    .io_salloc_req_0_bits_tail(ingress_unit_2_from_1_io_salloc_req_0_bits_tail),
    .io_out_0_valid(ingress_unit_2_from_1_io_out_0_valid),
    .io_out_0_bits_flit_head(ingress_unit_2_from_1_io_out_0_bits_flit_head),
    .io_out_0_bits_flit_tail(ingress_unit_2_from_1_io_out_0_bits_flit_tail),
    .io_out_0_bits_flit_payload(ingress_unit_2_from_1_io_out_0_bits_flit_payload),
    .io_out_0_bits_flit_flow_ingress_node(ingress_unit_2_from_1_io_out_0_bits_flit_flow_ingress_node),
    .io_out_0_bits_flit_flow_egress_node(ingress_unit_2_from_1_io_out_0_bits_flit_flow_egress_node),
    .io_out_0_bits_out_virt_channel(ingress_unit_2_from_1_io_out_0_bits_out_virt_channel),
    .io_in_ready(ingress_unit_2_from_1_io_in_ready),
    .io_in_valid(ingress_unit_2_from_1_io_in_valid),
    .io_in_bits_head(ingress_unit_2_from_1_io_in_bits_head),
    .io_in_bits_tail(ingress_unit_2_from_1_io_in_bits_tail),
    .io_in_bits_payload(ingress_unit_2_from_1_io_in_bits_payload),
    .io_in_bits_egress_id(ingress_unit_2_from_1_io_in_bits_egress_id)
  );
  OutputUnit output_unit_0_to_0 ( // @[Router.scala 122:13]
    .clock(output_unit_0_to_0_clock),
    .reset(output_unit_0_to_0_reset),
    .io_in_0_valid(output_unit_0_to_0_io_in_0_valid),
    .io_in_0_bits_head(output_unit_0_to_0_io_in_0_bits_head),
    .io_in_0_bits_tail(output_unit_0_to_0_io_in_0_bits_tail),
    .io_in_0_bits_payload(output_unit_0_to_0_io_in_0_bits_payload),
    .io_in_0_bits_flow_ingress_node(output_unit_0_to_0_io_in_0_bits_flow_ingress_node),
    .io_in_0_bits_flow_egress_node(output_unit_0_to_0_io_in_0_bits_flow_egress_node),
    .io_in_0_bits_virt_channel_id(output_unit_0_to_0_io_in_0_bits_virt_channel_id),
    .io_credit_available_0(output_unit_0_to_0_io_credit_available_0),
    .io_credit_available_1(output_unit_0_to_0_io_credit_available_1),
    .io_credit_available_2(output_unit_0_to_0_io_credit_available_2),
    .io_credit_available_3(output_unit_0_to_0_io_credit_available_3),
    .io_channel_status_0_occupied(output_unit_0_to_0_io_channel_status_0_occupied),
    .io_channel_status_1_occupied(output_unit_0_to_0_io_channel_status_1_occupied),
    .io_channel_status_2_occupied(output_unit_0_to_0_io_channel_status_2_occupied),
    .io_channel_status_3_occupied(output_unit_0_to_0_io_channel_status_3_occupied),
    .io_allocs_0_alloc(output_unit_0_to_0_io_allocs_0_alloc),
    .io_allocs_1_alloc(output_unit_0_to_0_io_allocs_1_alloc),
    .io_allocs_2_alloc(output_unit_0_to_0_io_allocs_2_alloc),
    .io_allocs_3_alloc(output_unit_0_to_0_io_allocs_3_alloc),
    .io_credit_alloc_0_alloc(output_unit_0_to_0_io_credit_alloc_0_alloc),
    .io_credit_alloc_1_alloc(output_unit_0_to_0_io_credit_alloc_1_alloc),
    .io_credit_alloc_2_alloc(output_unit_0_to_0_io_credit_alloc_2_alloc),
    .io_credit_alloc_3_alloc(output_unit_0_to_0_io_credit_alloc_3_alloc),
    .io_out_flit_0_valid(output_unit_0_to_0_io_out_flit_0_valid),
    .io_out_flit_0_bits_head(output_unit_0_to_0_io_out_flit_0_bits_head),
    .io_out_flit_0_bits_tail(output_unit_0_to_0_io_out_flit_0_bits_tail),
    .io_out_flit_0_bits_payload(output_unit_0_to_0_io_out_flit_0_bits_payload),
    .io_out_flit_0_bits_flow_ingress_node(output_unit_0_to_0_io_out_flit_0_bits_flow_ingress_node),
    .io_out_flit_0_bits_flow_egress_node(output_unit_0_to_0_io_out_flit_0_bits_flow_egress_node),
    .io_out_flit_0_bits_virt_channel_id(output_unit_0_to_0_io_out_flit_0_bits_virt_channel_id),
    .io_out_credit_return(output_unit_0_to_0_io_out_credit_return),
    .io_out_vc_free(output_unit_0_to_0_io_out_vc_free)
  );
  OutputUnit output_unit_1_to_2 ( // @[Router.scala 122:13]
    .clock(output_unit_1_to_2_clock),
    .reset(output_unit_1_to_2_reset),
    .io_in_0_valid(output_unit_1_to_2_io_in_0_valid),
    .io_in_0_bits_head(output_unit_1_to_2_io_in_0_bits_head),
    .io_in_0_bits_tail(output_unit_1_to_2_io_in_0_bits_tail),
    .io_in_0_bits_payload(output_unit_1_to_2_io_in_0_bits_payload),
    .io_in_0_bits_flow_ingress_node(output_unit_1_to_2_io_in_0_bits_flow_ingress_node),
    .io_in_0_bits_flow_egress_node(output_unit_1_to_2_io_in_0_bits_flow_egress_node),
    .io_in_0_bits_virt_channel_id(output_unit_1_to_2_io_in_0_bits_virt_channel_id),
    .io_credit_available_0(output_unit_1_to_2_io_credit_available_0),
    .io_credit_available_1(output_unit_1_to_2_io_credit_available_1),
    .io_credit_available_2(output_unit_1_to_2_io_credit_available_2),
    .io_credit_available_3(output_unit_1_to_2_io_credit_available_3),
    .io_channel_status_0_occupied(output_unit_1_to_2_io_channel_status_0_occupied),
    .io_channel_status_1_occupied(output_unit_1_to_2_io_channel_status_1_occupied),
    .io_channel_status_2_occupied(output_unit_1_to_2_io_channel_status_2_occupied),
    .io_channel_status_3_occupied(output_unit_1_to_2_io_channel_status_3_occupied),
    .io_allocs_0_alloc(output_unit_1_to_2_io_allocs_0_alloc),
    .io_allocs_1_alloc(output_unit_1_to_2_io_allocs_1_alloc),
    .io_allocs_2_alloc(output_unit_1_to_2_io_allocs_2_alloc),
    .io_allocs_3_alloc(output_unit_1_to_2_io_allocs_3_alloc),
    .io_credit_alloc_0_alloc(output_unit_1_to_2_io_credit_alloc_0_alloc),
    .io_credit_alloc_1_alloc(output_unit_1_to_2_io_credit_alloc_1_alloc),
    .io_credit_alloc_2_alloc(output_unit_1_to_2_io_credit_alloc_2_alloc),
    .io_credit_alloc_3_alloc(output_unit_1_to_2_io_credit_alloc_3_alloc),
    .io_out_flit_0_valid(output_unit_1_to_2_io_out_flit_0_valid),
    .io_out_flit_0_bits_head(output_unit_1_to_2_io_out_flit_0_bits_head),
    .io_out_flit_0_bits_tail(output_unit_1_to_2_io_out_flit_0_bits_tail),
    .io_out_flit_0_bits_payload(output_unit_1_to_2_io_out_flit_0_bits_payload),
    .io_out_flit_0_bits_flow_ingress_node(output_unit_1_to_2_io_out_flit_0_bits_flow_ingress_node),
    .io_out_flit_0_bits_flow_egress_node(output_unit_1_to_2_io_out_flit_0_bits_flow_egress_node),
    .io_out_flit_0_bits_virt_channel_id(output_unit_1_to_2_io_out_flit_0_bits_virt_channel_id),
    .io_out_credit_return(output_unit_1_to_2_io_out_credit_return),
    .io_out_vc_free(output_unit_1_to_2_io_out_vc_free)
  );
  EgressUnit egress_unit_2_to_1 ( // @[Router.scala 125:13]
    .clock(egress_unit_2_to_1_clock),
    .reset(egress_unit_2_to_1_reset),
    .io_in_0_valid(egress_unit_2_to_1_io_in_0_valid),
    .io_in_0_bits_head(egress_unit_2_to_1_io_in_0_bits_head),
    .io_in_0_bits_tail(egress_unit_2_to_1_io_in_0_bits_tail),
    .io_in_0_bits_payload(egress_unit_2_to_1_io_in_0_bits_payload),
    .io_in_0_bits_flow_ingress_node(egress_unit_2_to_1_io_in_0_bits_flow_ingress_node),
    .io_credit_available_0(egress_unit_2_to_1_io_credit_available_0),
    .io_channel_status_0_occupied(egress_unit_2_to_1_io_channel_status_0_occupied),
    .io_allocs_0_alloc(egress_unit_2_to_1_io_allocs_0_alloc),
    .io_credit_alloc_0_alloc(egress_unit_2_to_1_io_credit_alloc_0_alloc),
    .io_credit_alloc_0_tail(egress_unit_2_to_1_io_credit_alloc_0_tail),
    .io_out_valid(egress_unit_2_to_1_io_out_valid),
    .io_out_bits_head(egress_unit_2_to_1_io_out_bits_head),
    .io_out_bits_tail(egress_unit_2_to_1_io_out_bits_tail),
    .io_out_bits_payload(egress_unit_2_to_1_io_out_bits_payload),
    .io_out_bits_ingress_id(egress_unit_2_to_1_io_out_bits_ingress_id)
  );
  Switch switch ( // @[Router.scala 129:24]
    .clock(switch_clock),
    .reset(switch_reset),
    .io_in_2_0_valid(switch_io_in_2_0_valid),
    .io_in_2_0_bits_flit_head(switch_io_in_2_0_bits_flit_head),
    .io_in_2_0_bits_flit_tail(switch_io_in_2_0_bits_flit_tail),
    .io_in_2_0_bits_flit_payload(switch_io_in_2_0_bits_flit_payload),
    .io_in_2_0_bits_flit_flow_ingress_node(switch_io_in_2_0_bits_flit_flow_ingress_node),
    .io_in_2_0_bits_flit_flow_egress_node(switch_io_in_2_0_bits_flit_flow_egress_node),
    .io_in_2_0_bits_out_virt_channel(switch_io_in_2_0_bits_out_virt_channel),
    .io_in_1_0_valid(switch_io_in_1_0_valid),
    .io_in_1_0_bits_flit_head(switch_io_in_1_0_bits_flit_head),
    .io_in_1_0_bits_flit_tail(switch_io_in_1_0_bits_flit_tail),
    .io_in_1_0_bits_flit_payload(switch_io_in_1_0_bits_flit_payload),
    .io_in_1_0_bits_flit_flow_ingress_node(switch_io_in_1_0_bits_flit_flow_ingress_node),
    .io_in_1_0_bits_flit_flow_egress_node(switch_io_in_1_0_bits_flit_flow_egress_node),
    .io_in_1_0_bits_out_virt_channel(switch_io_in_1_0_bits_out_virt_channel),
    .io_in_0_0_valid(switch_io_in_0_0_valid),
    .io_in_0_0_bits_flit_head(switch_io_in_0_0_bits_flit_head),
    .io_in_0_0_bits_flit_tail(switch_io_in_0_0_bits_flit_tail),
    .io_in_0_0_bits_flit_payload(switch_io_in_0_0_bits_flit_payload),
    .io_in_0_0_bits_flit_flow_ingress_node(switch_io_in_0_0_bits_flit_flow_ingress_node),
    .io_in_0_0_bits_flit_flow_egress_node(switch_io_in_0_0_bits_flit_flow_egress_node),
    .io_in_0_0_bits_out_virt_channel(switch_io_in_0_0_bits_out_virt_channel),
    .io_out_2_0_valid(switch_io_out_2_0_valid),
    .io_out_2_0_bits_head(switch_io_out_2_0_bits_head),
    .io_out_2_0_bits_tail(switch_io_out_2_0_bits_tail),
    .io_out_2_0_bits_payload(switch_io_out_2_0_bits_payload),
    .io_out_2_0_bits_flow_ingress_node(switch_io_out_2_0_bits_flow_ingress_node),
    .io_out_1_0_valid(switch_io_out_1_0_valid),
    .io_out_1_0_bits_head(switch_io_out_1_0_bits_head),
    .io_out_1_0_bits_tail(switch_io_out_1_0_bits_tail),
    .io_out_1_0_bits_payload(switch_io_out_1_0_bits_payload),
    .io_out_1_0_bits_flow_ingress_node(switch_io_out_1_0_bits_flow_ingress_node),
    .io_out_1_0_bits_flow_egress_node(switch_io_out_1_0_bits_flow_egress_node),
    .io_out_1_0_bits_virt_channel_id(switch_io_out_1_0_bits_virt_channel_id),
    .io_out_0_0_valid(switch_io_out_0_0_valid),
    .io_out_0_0_bits_head(switch_io_out_0_0_bits_head),
    .io_out_0_0_bits_tail(switch_io_out_0_0_bits_tail),
    .io_out_0_0_bits_payload(switch_io_out_0_0_bits_payload),
    .io_out_0_0_bits_flow_ingress_node(switch_io_out_0_0_bits_flow_ingress_node),
    .io_out_0_0_bits_flow_egress_node(switch_io_out_0_0_bits_flow_egress_node),
    .io_out_0_0_bits_virt_channel_id(switch_io_out_0_0_bits_virt_channel_id),
    .io_sel_2_0_2_0(switch_io_sel_2_0_2_0),
    .io_sel_2_0_1_0(switch_io_sel_2_0_1_0),
    .io_sel_2_0_0_0(switch_io_sel_2_0_0_0),
    .io_sel_1_0_2_0(switch_io_sel_1_0_2_0),
    .io_sel_1_0_1_0(switch_io_sel_1_0_1_0),
    .io_sel_1_0_0_0(switch_io_sel_1_0_0_0),
    .io_sel_0_0_2_0(switch_io_sel_0_0_2_0),
    .io_sel_0_0_1_0(switch_io_sel_0_0_1_0),
    .io_sel_0_0_0_0(switch_io_sel_0_0_0_0)
  );
  SwitchAllocator switch_allocator ( // @[Router.scala 130:34]
    .clock(switch_allocator_clock),
    .reset(switch_allocator_reset),
    .io_req_2_0_ready(switch_allocator_io_req_2_0_ready),
    .io_req_2_0_valid(switch_allocator_io_req_2_0_valid),
    .io_req_2_0_bits_vc_sel_2_0(switch_allocator_io_req_2_0_bits_vc_sel_2_0),
    .io_req_2_0_bits_vc_sel_1_0(switch_allocator_io_req_2_0_bits_vc_sel_1_0),
    .io_req_2_0_bits_vc_sel_1_1(switch_allocator_io_req_2_0_bits_vc_sel_1_1),
    .io_req_2_0_bits_vc_sel_1_2(switch_allocator_io_req_2_0_bits_vc_sel_1_2),
    .io_req_2_0_bits_vc_sel_1_3(switch_allocator_io_req_2_0_bits_vc_sel_1_3),
    .io_req_2_0_bits_vc_sel_0_0(switch_allocator_io_req_2_0_bits_vc_sel_0_0),
    .io_req_2_0_bits_vc_sel_0_1(switch_allocator_io_req_2_0_bits_vc_sel_0_1),
    .io_req_2_0_bits_vc_sel_0_2(switch_allocator_io_req_2_0_bits_vc_sel_0_2),
    .io_req_2_0_bits_vc_sel_0_3(switch_allocator_io_req_2_0_bits_vc_sel_0_3),
    .io_req_2_0_bits_tail(switch_allocator_io_req_2_0_bits_tail),
    .io_req_1_0_ready(switch_allocator_io_req_1_0_ready),
    .io_req_1_0_valid(switch_allocator_io_req_1_0_valid),
    .io_req_1_0_bits_vc_sel_2_0(switch_allocator_io_req_1_0_bits_vc_sel_2_0),
    .io_req_1_0_bits_vc_sel_1_0(switch_allocator_io_req_1_0_bits_vc_sel_1_0),
    .io_req_1_0_bits_vc_sel_1_1(switch_allocator_io_req_1_0_bits_vc_sel_1_1),
    .io_req_1_0_bits_vc_sel_1_2(switch_allocator_io_req_1_0_bits_vc_sel_1_2),
    .io_req_1_0_bits_vc_sel_1_3(switch_allocator_io_req_1_0_bits_vc_sel_1_3),
    .io_req_1_0_bits_vc_sel_0_0(switch_allocator_io_req_1_0_bits_vc_sel_0_0),
    .io_req_1_0_bits_vc_sel_0_1(switch_allocator_io_req_1_0_bits_vc_sel_0_1),
    .io_req_1_0_bits_vc_sel_0_2(switch_allocator_io_req_1_0_bits_vc_sel_0_2),
    .io_req_1_0_bits_vc_sel_0_3(switch_allocator_io_req_1_0_bits_vc_sel_0_3),
    .io_req_1_0_bits_tail(switch_allocator_io_req_1_0_bits_tail),
    .io_req_0_0_ready(switch_allocator_io_req_0_0_ready),
    .io_req_0_0_valid(switch_allocator_io_req_0_0_valid),
    .io_req_0_0_bits_vc_sel_2_0(switch_allocator_io_req_0_0_bits_vc_sel_2_0),
    .io_req_0_0_bits_vc_sel_1_0(switch_allocator_io_req_0_0_bits_vc_sel_1_0),
    .io_req_0_0_bits_vc_sel_1_1(switch_allocator_io_req_0_0_bits_vc_sel_1_1),
    .io_req_0_0_bits_vc_sel_1_2(switch_allocator_io_req_0_0_bits_vc_sel_1_2),
    .io_req_0_0_bits_vc_sel_1_3(switch_allocator_io_req_0_0_bits_vc_sel_1_3),
    .io_req_0_0_bits_vc_sel_0_0(switch_allocator_io_req_0_0_bits_vc_sel_0_0),
    .io_req_0_0_bits_vc_sel_0_1(switch_allocator_io_req_0_0_bits_vc_sel_0_1),
    .io_req_0_0_bits_vc_sel_0_2(switch_allocator_io_req_0_0_bits_vc_sel_0_2),
    .io_req_0_0_bits_vc_sel_0_3(switch_allocator_io_req_0_0_bits_vc_sel_0_3),
    .io_req_0_0_bits_tail(switch_allocator_io_req_0_0_bits_tail),
    .io_credit_alloc_2_0_alloc(switch_allocator_io_credit_alloc_2_0_alloc),
    .io_credit_alloc_2_0_tail(switch_allocator_io_credit_alloc_2_0_tail),
    .io_credit_alloc_1_0_alloc(switch_allocator_io_credit_alloc_1_0_alloc),
    .io_credit_alloc_1_1_alloc(switch_allocator_io_credit_alloc_1_1_alloc),
    .io_credit_alloc_1_2_alloc(switch_allocator_io_credit_alloc_1_2_alloc),
    .io_credit_alloc_1_3_alloc(switch_allocator_io_credit_alloc_1_3_alloc),
    .io_credit_alloc_0_0_alloc(switch_allocator_io_credit_alloc_0_0_alloc),
    .io_credit_alloc_0_1_alloc(switch_allocator_io_credit_alloc_0_1_alloc),
    .io_credit_alloc_0_2_alloc(switch_allocator_io_credit_alloc_0_2_alloc),
    .io_credit_alloc_0_3_alloc(switch_allocator_io_credit_alloc_0_3_alloc),
    .io_switch_sel_2_0_2_0(switch_allocator_io_switch_sel_2_0_2_0),
    .io_switch_sel_2_0_1_0(switch_allocator_io_switch_sel_2_0_1_0),
    .io_switch_sel_2_0_0_0(switch_allocator_io_switch_sel_2_0_0_0),
    .io_switch_sel_1_0_2_0(switch_allocator_io_switch_sel_1_0_2_0),
    .io_switch_sel_1_0_1_0(switch_allocator_io_switch_sel_1_0_1_0),
    .io_switch_sel_1_0_0_0(switch_allocator_io_switch_sel_1_0_0_0),
    .io_switch_sel_0_0_2_0(switch_allocator_io_switch_sel_0_0_2_0),
    .io_switch_sel_0_0_1_0(switch_allocator_io_switch_sel_0_0_1_0),
    .io_switch_sel_0_0_0_0(switch_allocator_io_switch_sel_0_0_0_0)
  );
  RotatingSingleVCAllocator vc_allocator ( // @[Router.scala 131:30]
    .clock(vc_allocator_clock),
    .reset(vc_allocator_reset),
    .io_req_2_ready(vc_allocator_io_req_2_ready),
    .io_req_2_valid(vc_allocator_io_req_2_valid),
    .io_req_2_bits_vc_sel_2_0(vc_allocator_io_req_2_bits_vc_sel_2_0),
    .io_req_2_bits_vc_sel_1_0(vc_allocator_io_req_2_bits_vc_sel_1_0),
    .io_req_2_bits_vc_sel_1_1(vc_allocator_io_req_2_bits_vc_sel_1_1),
    .io_req_2_bits_vc_sel_1_2(vc_allocator_io_req_2_bits_vc_sel_1_2),
    .io_req_2_bits_vc_sel_1_3(vc_allocator_io_req_2_bits_vc_sel_1_3),
    .io_req_2_bits_vc_sel_0_0(vc_allocator_io_req_2_bits_vc_sel_0_0),
    .io_req_2_bits_vc_sel_0_1(vc_allocator_io_req_2_bits_vc_sel_0_1),
    .io_req_2_bits_vc_sel_0_2(vc_allocator_io_req_2_bits_vc_sel_0_2),
    .io_req_2_bits_vc_sel_0_3(vc_allocator_io_req_2_bits_vc_sel_0_3),
    .io_req_1_ready(vc_allocator_io_req_1_ready),
    .io_req_1_valid(vc_allocator_io_req_1_valid),
    .io_req_1_bits_vc_sel_2_0(vc_allocator_io_req_1_bits_vc_sel_2_0),
    .io_req_1_bits_vc_sel_1_0(vc_allocator_io_req_1_bits_vc_sel_1_0),
    .io_req_1_bits_vc_sel_1_1(vc_allocator_io_req_1_bits_vc_sel_1_1),
    .io_req_1_bits_vc_sel_1_2(vc_allocator_io_req_1_bits_vc_sel_1_2),
    .io_req_1_bits_vc_sel_1_3(vc_allocator_io_req_1_bits_vc_sel_1_3),
    .io_req_1_bits_vc_sel_0_0(vc_allocator_io_req_1_bits_vc_sel_0_0),
    .io_req_1_bits_vc_sel_0_1(vc_allocator_io_req_1_bits_vc_sel_0_1),
    .io_req_1_bits_vc_sel_0_2(vc_allocator_io_req_1_bits_vc_sel_0_2),
    .io_req_1_bits_vc_sel_0_3(vc_allocator_io_req_1_bits_vc_sel_0_3),
    .io_req_0_ready(vc_allocator_io_req_0_ready),
    .io_req_0_valid(vc_allocator_io_req_0_valid),
    .io_req_0_bits_vc_sel_2_0(vc_allocator_io_req_0_bits_vc_sel_2_0),
    .io_req_0_bits_vc_sel_1_0(vc_allocator_io_req_0_bits_vc_sel_1_0),
    .io_req_0_bits_vc_sel_1_1(vc_allocator_io_req_0_bits_vc_sel_1_1),
    .io_req_0_bits_vc_sel_1_2(vc_allocator_io_req_0_bits_vc_sel_1_2),
    .io_req_0_bits_vc_sel_1_3(vc_allocator_io_req_0_bits_vc_sel_1_3),
    .io_req_0_bits_vc_sel_0_0(vc_allocator_io_req_0_bits_vc_sel_0_0),
    .io_req_0_bits_vc_sel_0_1(vc_allocator_io_req_0_bits_vc_sel_0_1),
    .io_req_0_bits_vc_sel_0_2(vc_allocator_io_req_0_bits_vc_sel_0_2),
    .io_req_0_bits_vc_sel_0_3(vc_allocator_io_req_0_bits_vc_sel_0_3),
    .io_resp_2_vc_sel_2_0(vc_allocator_io_resp_2_vc_sel_2_0),
    .io_resp_2_vc_sel_1_0(vc_allocator_io_resp_2_vc_sel_1_0),
    .io_resp_2_vc_sel_1_1(vc_allocator_io_resp_2_vc_sel_1_1),
    .io_resp_2_vc_sel_1_2(vc_allocator_io_resp_2_vc_sel_1_2),
    .io_resp_2_vc_sel_1_3(vc_allocator_io_resp_2_vc_sel_1_3),
    .io_resp_2_vc_sel_0_0(vc_allocator_io_resp_2_vc_sel_0_0),
    .io_resp_2_vc_sel_0_1(vc_allocator_io_resp_2_vc_sel_0_1),
    .io_resp_2_vc_sel_0_2(vc_allocator_io_resp_2_vc_sel_0_2),
    .io_resp_2_vc_sel_0_3(vc_allocator_io_resp_2_vc_sel_0_3),
    .io_resp_1_vc_sel_2_0(vc_allocator_io_resp_1_vc_sel_2_0),
    .io_resp_1_vc_sel_1_0(vc_allocator_io_resp_1_vc_sel_1_0),
    .io_resp_1_vc_sel_1_1(vc_allocator_io_resp_1_vc_sel_1_1),
    .io_resp_1_vc_sel_1_2(vc_allocator_io_resp_1_vc_sel_1_2),
    .io_resp_1_vc_sel_1_3(vc_allocator_io_resp_1_vc_sel_1_3),
    .io_resp_1_vc_sel_0_0(vc_allocator_io_resp_1_vc_sel_0_0),
    .io_resp_1_vc_sel_0_1(vc_allocator_io_resp_1_vc_sel_0_1),
    .io_resp_1_vc_sel_0_2(vc_allocator_io_resp_1_vc_sel_0_2),
    .io_resp_1_vc_sel_0_3(vc_allocator_io_resp_1_vc_sel_0_3),
    .io_resp_0_vc_sel_2_0(vc_allocator_io_resp_0_vc_sel_2_0),
    .io_resp_0_vc_sel_1_0(vc_allocator_io_resp_0_vc_sel_1_0),
    .io_resp_0_vc_sel_1_1(vc_allocator_io_resp_0_vc_sel_1_1),
    .io_resp_0_vc_sel_1_2(vc_allocator_io_resp_0_vc_sel_1_2),
    .io_resp_0_vc_sel_1_3(vc_allocator_io_resp_0_vc_sel_1_3),
    .io_resp_0_vc_sel_0_0(vc_allocator_io_resp_0_vc_sel_0_0),
    .io_resp_0_vc_sel_0_1(vc_allocator_io_resp_0_vc_sel_0_1),
    .io_resp_0_vc_sel_0_2(vc_allocator_io_resp_0_vc_sel_0_2),
    .io_resp_0_vc_sel_0_3(vc_allocator_io_resp_0_vc_sel_0_3),
    .io_channel_status_2_0_occupied(vc_allocator_io_channel_status_2_0_occupied),
    .io_channel_status_1_0_occupied(vc_allocator_io_channel_status_1_0_occupied),
    .io_channel_status_1_1_occupied(vc_allocator_io_channel_status_1_1_occupied),
    .io_channel_status_1_2_occupied(vc_allocator_io_channel_status_1_2_occupied),
    .io_channel_status_1_3_occupied(vc_allocator_io_channel_status_1_3_occupied),
    .io_channel_status_0_0_occupied(vc_allocator_io_channel_status_0_0_occupied),
    .io_channel_status_0_1_occupied(vc_allocator_io_channel_status_0_1_occupied),
    .io_channel_status_0_2_occupied(vc_allocator_io_channel_status_0_2_occupied),
    .io_channel_status_0_3_occupied(vc_allocator_io_channel_status_0_3_occupied),
    .io_out_allocs_2_0_alloc(vc_allocator_io_out_allocs_2_0_alloc),
    .io_out_allocs_1_0_alloc(vc_allocator_io_out_allocs_1_0_alloc),
    .io_out_allocs_1_1_alloc(vc_allocator_io_out_allocs_1_1_alloc),
    .io_out_allocs_1_2_alloc(vc_allocator_io_out_allocs_1_2_alloc),
    .io_out_allocs_1_3_alloc(vc_allocator_io_out_allocs_1_3_alloc),
    .io_out_allocs_0_0_alloc(vc_allocator_io_out_allocs_0_0_alloc),
    .io_out_allocs_0_1_alloc(vc_allocator_io_out_allocs_0_1_alloc),
    .io_out_allocs_0_2_alloc(vc_allocator_io_out_allocs_0_2_alloc),
    .io_out_allocs_0_3_alloc(vc_allocator_io_out_allocs_0_3_alloc)
  );
  RouteComputer_1 route_computer ( // @[Router.scala 134:32]
    .io_req_2_bits_flow_ingress_node(route_computer_io_req_2_bits_flow_ingress_node),
    .io_req_2_bits_flow_egress_node(route_computer_io_req_2_bits_flow_egress_node),
    .io_req_1_bits_src_virt_id(route_computer_io_req_1_bits_src_virt_id),
    .io_req_1_bits_flow_ingress_node(route_computer_io_req_1_bits_flow_ingress_node),
    .io_req_1_bits_flow_egress_node(route_computer_io_req_1_bits_flow_egress_node),
    .io_req_0_bits_src_virt_id(route_computer_io_req_0_bits_src_virt_id),
    .io_req_0_bits_flow_ingress_node(route_computer_io_req_0_bits_flow_ingress_node),
    .io_req_0_bits_flow_egress_node(route_computer_io_req_0_bits_flow_egress_node),
    .io_resp_2_vc_sel_1_0(route_computer_io_resp_2_vc_sel_1_0),
    .io_resp_2_vc_sel_1_1(route_computer_io_resp_2_vc_sel_1_1),
    .io_resp_2_vc_sel_1_2(route_computer_io_resp_2_vc_sel_1_2),
    .io_resp_2_vc_sel_1_3(route_computer_io_resp_2_vc_sel_1_3),
    .io_resp_2_vc_sel_0_0(route_computer_io_resp_2_vc_sel_0_0),
    .io_resp_2_vc_sel_0_1(route_computer_io_resp_2_vc_sel_0_1),
    .io_resp_2_vc_sel_0_2(route_computer_io_resp_2_vc_sel_0_2),
    .io_resp_2_vc_sel_0_3(route_computer_io_resp_2_vc_sel_0_3),
    .io_resp_1_vc_sel_1_0(route_computer_io_resp_1_vc_sel_1_0),
    .io_resp_1_vc_sel_1_1(route_computer_io_resp_1_vc_sel_1_1),
    .io_resp_1_vc_sel_1_2(route_computer_io_resp_1_vc_sel_1_2),
    .io_resp_1_vc_sel_1_3(route_computer_io_resp_1_vc_sel_1_3),
    .io_resp_1_vc_sel_0_0(route_computer_io_resp_1_vc_sel_0_0),
    .io_resp_1_vc_sel_0_1(route_computer_io_resp_1_vc_sel_0_1),
    .io_resp_1_vc_sel_0_2(route_computer_io_resp_1_vc_sel_0_2),
    .io_resp_1_vc_sel_0_3(route_computer_io_resp_1_vc_sel_0_3),
    .io_resp_0_vc_sel_1_0(route_computer_io_resp_0_vc_sel_1_0),
    .io_resp_0_vc_sel_1_1(route_computer_io_resp_0_vc_sel_1_1),
    .io_resp_0_vc_sel_1_2(route_computer_io_resp_0_vc_sel_1_2),
    .io_resp_0_vc_sel_1_3(route_computer_io_resp_0_vc_sel_1_3),
    .io_resp_0_vc_sel_0_0(route_computer_io_resp_0_vc_sel_0_0),
    .io_resp_0_vc_sel_0_1(route_computer_io_resp_0_vc_sel_0_1),
    .io_resp_0_vc_sel_0_2(route_computer_io_resp_0_vc_sel_0_2),
    .io_resp_0_vc_sel_0_3(route_computer_io_resp_0_vc_sel_0_3)
  );
  plusarg_reader #(.FORMAT("noc_util_sample_rate=%d"), .DEFAULT(0), .WIDTH(20)) plusarg_reader ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_out)
  );
  assign auto_debug_out_va_stall_0 = input_unit_0_from_0_io_debug_va_stall; // @[Nodes.scala 1212:84 Router.scala 190:92]
  assign auto_debug_out_va_stall_1 = input_unit_1_from_2_io_debug_va_stall; // @[Nodes.scala 1212:84 Router.scala 190:92]
  assign auto_debug_out_sa_stall_0 = input_unit_0_from_0_io_debug_sa_stall; // @[Nodes.scala 1212:84 Router.scala 191:92]
  assign auto_debug_out_sa_stall_1 = input_unit_1_from_2_io_debug_sa_stall; // @[Nodes.scala 1212:84 Router.scala 191:92]
  assign auto_egress_nodes_out_flit_valid = egress_unit_2_to_1_io_out_valid; // @[Nodes.scala 1212:84 Router.scala 144:65]
  assign auto_egress_nodes_out_flit_bits_head = egress_unit_2_to_1_io_out_bits_head; // @[Nodes.scala 1212:84 Router.scala 144:65]
  assign auto_egress_nodes_out_flit_bits_tail = egress_unit_2_to_1_io_out_bits_tail; // @[Nodes.scala 1212:84 Router.scala 144:65]
  assign auto_egress_nodes_out_flit_bits_payload = egress_unit_2_to_1_io_out_bits_payload; // @[Nodes.scala 1212:84 Router.scala 144:65]
  assign auto_egress_nodes_out_flit_bits_ingress_id = egress_unit_2_to_1_io_out_bits_ingress_id; // @[Nodes.scala 1212:84 Router.scala 144:65]
  assign auto_ingress_nodes_in_flit_ready = ingress_unit_2_from_1_io_in_ready; // @[Nodes.scala 1215:84 Router.scala 142:68]
  assign auto_source_nodes_out_1_flit_0_valid = output_unit_1_to_2_io_out_flit_0_valid; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_1_flit_0_bits_head = output_unit_1_to_2_io_out_flit_0_bits_head; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_1_flit_0_bits_tail = output_unit_1_to_2_io_out_flit_0_bits_tail; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_1_flit_0_bits_payload = output_unit_1_to_2_io_out_flit_0_bits_payload; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_1_flit_0_bits_flow_ingress_node = output_unit_1_to_2_io_out_flit_0_bits_flow_ingress_node
    ; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_1_flit_0_bits_flow_egress_node = output_unit_1_to_2_io_out_flit_0_bits_flow_egress_node; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_1_flit_0_bits_virt_channel_id = output_unit_1_to_2_io_out_flit_0_bits_virt_channel_id; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_0_flit_0_valid = output_unit_0_to_0_io_out_flit_0_valid; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_0_flit_0_bits_head = output_unit_0_to_0_io_out_flit_0_bits_head; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_0_flit_0_bits_tail = output_unit_0_to_0_io_out_flit_0_bits_tail; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_0_flit_0_bits_payload = output_unit_0_to_0_io_out_flit_0_bits_payload; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_0_flit_0_bits_flow_ingress_node = output_unit_0_to_0_io_out_flit_0_bits_flow_ingress_node
    ; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_0_flit_0_bits_flow_egress_node = output_unit_0_to_0_io_out_flit_0_bits_flow_egress_node; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_0_flit_0_bits_virt_channel_id = output_unit_0_to_0_io_out_flit_0_bits_virt_channel_id; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_dest_nodes_in_1_credit_return = input_unit_1_from_2_io_in_credit_return; // @[Nodes.scala 1215:84 Router.scala 141:68]
  assign auto_dest_nodes_in_1_vc_free = input_unit_1_from_2_io_in_vc_free; // @[Nodes.scala 1215:84 Router.scala 141:68]
  assign auto_dest_nodes_in_0_credit_return = input_unit_0_from_0_io_in_credit_return; // @[Nodes.scala 1215:84 Router.scala 141:68]
  assign auto_dest_nodes_in_0_vc_free = input_unit_0_from_0_io_in_vc_free; // @[Nodes.scala 1215:84 Router.scala 141:68]
  assign monitor_clock = clock;
  assign monitor_reset = reset;
  assign monitor_io_in_flit_0_valid = auto_dest_nodes_in_0_flit_0_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_io_in_flit_0_bits_head = auto_dest_nodes_in_0_flit_0_bits_head; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_io_in_flit_0_bits_tail = auto_dest_nodes_in_0_flit_0_bits_tail; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_io_in_flit_0_bits_flow_ingress_node = auto_dest_nodes_in_0_flit_0_bits_flow_ingress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_io_in_flit_0_bits_flow_egress_node = auto_dest_nodes_in_0_flit_0_bits_flow_egress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_io_in_flit_0_bits_virt_channel_id = auto_dest_nodes_in_0_flit_0_bits_virt_channel_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_1_clock = clock;
  assign monitor_1_reset = reset;
  assign monitor_1_io_in_flit_0_valid = auto_dest_nodes_in_1_flit_0_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_1_io_in_flit_0_bits_head = auto_dest_nodes_in_1_flit_0_bits_head; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_1_io_in_flit_0_bits_tail = auto_dest_nodes_in_1_flit_0_bits_tail; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_1_io_in_flit_0_bits_flow_ingress_node = auto_dest_nodes_in_1_flit_0_bits_flow_ingress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_1_io_in_flit_0_bits_flow_egress_node = auto_dest_nodes_in_1_flit_0_bits_flow_egress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_1_io_in_flit_0_bits_virt_channel_id = auto_dest_nodes_in_1_flit_0_bits_virt_channel_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_0_clock = clock;
  assign input_unit_0_from_0_reset = reset;
  assign input_unit_0_from_0_io_router_resp_vc_sel_1_0 = route_computer_io_resp_0_vc_sel_1_0; // @[Router.scala 148:38]
  assign input_unit_0_from_0_io_router_resp_vc_sel_1_1 = route_computer_io_resp_0_vc_sel_1_1; // @[Router.scala 148:38]
  assign input_unit_0_from_0_io_router_resp_vc_sel_1_2 = route_computer_io_resp_0_vc_sel_1_2; // @[Router.scala 148:38]
  assign input_unit_0_from_0_io_router_resp_vc_sel_1_3 = route_computer_io_resp_0_vc_sel_1_3; // @[Router.scala 148:38]
  assign input_unit_0_from_0_io_router_resp_vc_sel_0_0 = route_computer_io_resp_0_vc_sel_0_0; // @[Router.scala 148:38]
  assign input_unit_0_from_0_io_router_resp_vc_sel_0_1 = route_computer_io_resp_0_vc_sel_0_1; // @[Router.scala 148:38]
  assign input_unit_0_from_0_io_router_resp_vc_sel_0_2 = route_computer_io_resp_0_vc_sel_0_2; // @[Router.scala 148:38]
  assign input_unit_0_from_0_io_router_resp_vc_sel_0_3 = route_computer_io_resp_0_vc_sel_0_3; // @[Router.scala 148:38]
  assign input_unit_0_from_0_io_vcalloc_req_ready = vc_allocator_io_req_0_ready; // @[Router.scala 151:23]
  assign input_unit_0_from_0_io_vcalloc_resp_vc_sel_2_0 = vc_allocator_io_resp_0_vc_sel_2_0; // @[Router.scala 153:39]
  assign input_unit_0_from_0_io_vcalloc_resp_vc_sel_1_0 = vc_allocator_io_resp_0_vc_sel_1_0; // @[Router.scala 153:39]
  assign input_unit_0_from_0_io_vcalloc_resp_vc_sel_1_1 = vc_allocator_io_resp_0_vc_sel_1_1; // @[Router.scala 153:39]
  assign input_unit_0_from_0_io_vcalloc_resp_vc_sel_1_2 = vc_allocator_io_resp_0_vc_sel_1_2; // @[Router.scala 153:39]
  assign input_unit_0_from_0_io_vcalloc_resp_vc_sel_1_3 = vc_allocator_io_resp_0_vc_sel_1_3; // @[Router.scala 153:39]
  assign input_unit_0_from_0_io_vcalloc_resp_vc_sel_0_0 = vc_allocator_io_resp_0_vc_sel_0_0; // @[Router.scala 153:39]
  assign input_unit_0_from_0_io_vcalloc_resp_vc_sel_0_1 = vc_allocator_io_resp_0_vc_sel_0_1; // @[Router.scala 153:39]
  assign input_unit_0_from_0_io_vcalloc_resp_vc_sel_0_2 = vc_allocator_io_resp_0_vc_sel_0_2; // @[Router.scala 153:39]
  assign input_unit_0_from_0_io_vcalloc_resp_vc_sel_0_3 = vc_allocator_io_resp_0_vc_sel_0_3; // @[Router.scala 153:39]
  assign input_unit_0_from_0_io_out_credit_available_2_0 = egress_unit_2_to_1_io_credit_available_0; // @[Router.scala 162:42]
  assign input_unit_0_from_0_io_out_credit_available_1_0 = output_unit_1_to_2_io_credit_available_0; // @[Router.scala 162:42]
  assign input_unit_0_from_0_io_out_credit_available_1_1 = output_unit_1_to_2_io_credit_available_1; // @[Router.scala 162:42]
  assign input_unit_0_from_0_io_out_credit_available_1_2 = output_unit_1_to_2_io_credit_available_2; // @[Router.scala 162:42]
  assign input_unit_0_from_0_io_out_credit_available_1_3 = output_unit_1_to_2_io_credit_available_3; // @[Router.scala 162:42]
  assign input_unit_0_from_0_io_out_credit_available_0_0 = output_unit_0_to_0_io_credit_available_0; // @[Router.scala 162:42]
  assign input_unit_0_from_0_io_out_credit_available_0_1 = output_unit_0_to_0_io_credit_available_1; // @[Router.scala 162:42]
  assign input_unit_0_from_0_io_out_credit_available_0_2 = output_unit_0_to_0_io_credit_available_2; // @[Router.scala 162:42]
  assign input_unit_0_from_0_io_out_credit_available_0_3 = output_unit_0_to_0_io_credit_available_3; // @[Router.scala 162:42]
  assign input_unit_0_from_0_io_salloc_req_0_ready = switch_allocator_io_req_0_0_ready; // @[Router.scala 165:23]
  assign input_unit_0_from_0_io_in_flit_0_valid = auto_dest_nodes_in_0_flit_0_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_0_io_in_flit_0_bits_head = auto_dest_nodes_in_0_flit_0_bits_head; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_0_io_in_flit_0_bits_tail = auto_dest_nodes_in_0_flit_0_bits_tail; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_0_io_in_flit_0_bits_payload = auto_dest_nodes_in_0_flit_0_bits_payload; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_0_io_in_flit_0_bits_flow_ingress_node = auto_dest_nodes_in_0_flit_0_bits_flow_ingress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_0_io_in_flit_0_bits_flow_egress_node = auto_dest_nodes_in_0_flit_0_bits_flow_egress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_0_io_in_flit_0_bits_virt_channel_id = auto_dest_nodes_in_0_flit_0_bits_virt_channel_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_1_from_2_clock = clock;
  assign input_unit_1_from_2_reset = reset;
  assign input_unit_1_from_2_io_router_resp_vc_sel_1_0 = route_computer_io_resp_1_vc_sel_1_0; // @[Router.scala 148:38]
  assign input_unit_1_from_2_io_router_resp_vc_sel_1_1 = route_computer_io_resp_1_vc_sel_1_1; // @[Router.scala 148:38]
  assign input_unit_1_from_2_io_router_resp_vc_sel_1_2 = route_computer_io_resp_1_vc_sel_1_2; // @[Router.scala 148:38]
  assign input_unit_1_from_2_io_router_resp_vc_sel_1_3 = route_computer_io_resp_1_vc_sel_1_3; // @[Router.scala 148:38]
  assign input_unit_1_from_2_io_router_resp_vc_sel_0_0 = route_computer_io_resp_1_vc_sel_0_0; // @[Router.scala 148:38]
  assign input_unit_1_from_2_io_router_resp_vc_sel_0_1 = route_computer_io_resp_1_vc_sel_0_1; // @[Router.scala 148:38]
  assign input_unit_1_from_2_io_router_resp_vc_sel_0_2 = route_computer_io_resp_1_vc_sel_0_2; // @[Router.scala 148:38]
  assign input_unit_1_from_2_io_router_resp_vc_sel_0_3 = route_computer_io_resp_1_vc_sel_0_3; // @[Router.scala 148:38]
  assign input_unit_1_from_2_io_vcalloc_req_ready = vc_allocator_io_req_1_ready; // @[Router.scala 151:23]
  assign input_unit_1_from_2_io_vcalloc_resp_vc_sel_2_0 = vc_allocator_io_resp_1_vc_sel_2_0; // @[Router.scala 153:39]
  assign input_unit_1_from_2_io_vcalloc_resp_vc_sel_1_0 = vc_allocator_io_resp_1_vc_sel_1_0; // @[Router.scala 153:39]
  assign input_unit_1_from_2_io_vcalloc_resp_vc_sel_1_1 = vc_allocator_io_resp_1_vc_sel_1_1; // @[Router.scala 153:39]
  assign input_unit_1_from_2_io_vcalloc_resp_vc_sel_1_2 = vc_allocator_io_resp_1_vc_sel_1_2; // @[Router.scala 153:39]
  assign input_unit_1_from_2_io_vcalloc_resp_vc_sel_1_3 = vc_allocator_io_resp_1_vc_sel_1_3; // @[Router.scala 153:39]
  assign input_unit_1_from_2_io_vcalloc_resp_vc_sel_0_0 = vc_allocator_io_resp_1_vc_sel_0_0; // @[Router.scala 153:39]
  assign input_unit_1_from_2_io_vcalloc_resp_vc_sel_0_1 = vc_allocator_io_resp_1_vc_sel_0_1; // @[Router.scala 153:39]
  assign input_unit_1_from_2_io_vcalloc_resp_vc_sel_0_2 = vc_allocator_io_resp_1_vc_sel_0_2; // @[Router.scala 153:39]
  assign input_unit_1_from_2_io_vcalloc_resp_vc_sel_0_3 = vc_allocator_io_resp_1_vc_sel_0_3; // @[Router.scala 153:39]
  assign input_unit_1_from_2_io_out_credit_available_2_0 = egress_unit_2_to_1_io_credit_available_0; // @[Router.scala 162:42]
  assign input_unit_1_from_2_io_out_credit_available_1_0 = output_unit_1_to_2_io_credit_available_0; // @[Router.scala 162:42]
  assign input_unit_1_from_2_io_out_credit_available_1_1 = output_unit_1_to_2_io_credit_available_1; // @[Router.scala 162:42]
  assign input_unit_1_from_2_io_out_credit_available_1_2 = output_unit_1_to_2_io_credit_available_2; // @[Router.scala 162:42]
  assign input_unit_1_from_2_io_out_credit_available_1_3 = output_unit_1_to_2_io_credit_available_3; // @[Router.scala 162:42]
  assign input_unit_1_from_2_io_out_credit_available_0_0 = output_unit_0_to_0_io_credit_available_0; // @[Router.scala 162:42]
  assign input_unit_1_from_2_io_out_credit_available_0_1 = output_unit_0_to_0_io_credit_available_1; // @[Router.scala 162:42]
  assign input_unit_1_from_2_io_out_credit_available_0_2 = output_unit_0_to_0_io_credit_available_2; // @[Router.scala 162:42]
  assign input_unit_1_from_2_io_out_credit_available_0_3 = output_unit_0_to_0_io_credit_available_3; // @[Router.scala 162:42]
  assign input_unit_1_from_2_io_salloc_req_0_ready = switch_allocator_io_req_1_0_ready; // @[Router.scala 165:23]
  assign input_unit_1_from_2_io_in_flit_0_valid = auto_dest_nodes_in_1_flit_0_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_1_from_2_io_in_flit_0_bits_head = auto_dest_nodes_in_1_flit_0_bits_head; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_1_from_2_io_in_flit_0_bits_tail = auto_dest_nodes_in_1_flit_0_bits_tail; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_1_from_2_io_in_flit_0_bits_payload = auto_dest_nodes_in_1_flit_0_bits_payload; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_1_from_2_io_in_flit_0_bits_flow_ingress_node = auto_dest_nodes_in_1_flit_0_bits_flow_ingress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_1_from_2_io_in_flit_0_bits_flow_egress_node = auto_dest_nodes_in_1_flit_0_bits_flow_egress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_1_from_2_io_in_flit_0_bits_virt_channel_id = auto_dest_nodes_in_1_flit_0_bits_virt_channel_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign ingress_unit_2_from_1_clock = clock;
  assign ingress_unit_2_from_1_reset = reset;
  assign ingress_unit_2_from_1_io_router_resp_vc_sel_1_0 = route_computer_io_resp_2_vc_sel_1_0; // @[Router.scala 148:38]
  assign ingress_unit_2_from_1_io_router_resp_vc_sel_1_1 = route_computer_io_resp_2_vc_sel_1_1; // @[Router.scala 148:38]
  assign ingress_unit_2_from_1_io_router_resp_vc_sel_1_2 = route_computer_io_resp_2_vc_sel_1_2; // @[Router.scala 148:38]
  assign ingress_unit_2_from_1_io_router_resp_vc_sel_1_3 = route_computer_io_resp_2_vc_sel_1_3; // @[Router.scala 148:38]
  assign ingress_unit_2_from_1_io_router_resp_vc_sel_0_0 = route_computer_io_resp_2_vc_sel_0_0; // @[Router.scala 148:38]
  assign ingress_unit_2_from_1_io_router_resp_vc_sel_0_1 = route_computer_io_resp_2_vc_sel_0_1; // @[Router.scala 148:38]
  assign ingress_unit_2_from_1_io_router_resp_vc_sel_0_2 = route_computer_io_resp_2_vc_sel_0_2; // @[Router.scala 148:38]
  assign ingress_unit_2_from_1_io_router_resp_vc_sel_0_3 = route_computer_io_resp_2_vc_sel_0_3; // @[Router.scala 148:38]
  assign ingress_unit_2_from_1_io_vcalloc_req_ready = vc_allocator_io_req_2_ready; // @[Router.scala 151:23]
  assign ingress_unit_2_from_1_io_vcalloc_resp_vc_sel_2_0 = vc_allocator_io_resp_2_vc_sel_2_0; // @[Router.scala 153:39]
  assign ingress_unit_2_from_1_io_vcalloc_resp_vc_sel_1_0 = vc_allocator_io_resp_2_vc_sel_1_0; // @[Router.scala 153:39]
  assign ingress_unit_2_from_1_io_vcalloc_resp_vc_sel_1_1 = vc_allocator_io_resp_2_vc_sel_1_1; // @[Router.scala 153:39]
  assign ingress_unit_2_from_1_io_vcalloc_resp_vc_sel_1_2 = vc_allocator_io_resp_2_vc_sel_1_2; // @[Router.scala 153:39]
  assign ingress_unit_2_from_1_io_vcalloc_resp_vc_sel_1_3 = vc_allocator_io_resp_2_vc_sel_1_3; // @[Router.scala 153:39]
  assign ingress_unit_2_from_1_io_vcalloc_resp_vc_sel_0_0 = vc_allocator_io_resp_2_vc_sel_0_0; // @[Router.scala 153:39]
  assign ingress_unit_2_from_1_io_vcalloc_resp_vc_sel_0_1 = vc_allocator_io_resp_2_vc_sel_0_1; // @[Router.scala 153:39]
  assign ingress_unit_2_from_1_io_vcalloc_resp_vc_sel_0_2 = vc_allocator_io_resp_2_vc_sel_0_2; // @[Router.scala 153:39]
  assign ingress_unit_2_from_1_io_vcalloc_resp_vc_sel_0_3 = vc_allocator_io_resp_2_vc_sel_0_3; // @[Router.scala 153:39]
  assign ingress_unit_2_from_1_io_out_credit_available_2_0 = egress_unit_2_to_1_io_credit_available_0; // @[Router.scala 162:42]
  assign ingress_unit_2_from_1_io_out_credit_available_1_0 = output_unit_1_to_2_io_credit_available_0; // @[Router.scala 162:42]
  assign ingress_unit_2_from_1_io_out_credit_available_1_1 = output_unit_1_to_2_io_credit_available_1; // @[Router.scala 162:42]
  assign ingress_unit_2_from_1_io_out_credit_available_1_2 = output_unit_1_to_2_io_credit_available_2; // @[Router.scala 162:42]
  assign ingress_unit_2_from_1_io_out_credit_available_1_3 = output_unit_1_to_2_io_credit_available_3; // @[Router.scala 162:42]
  assign ingress_unit_2_from_1_io_out_credit_available_0_0 = output_unit_0_to_0_io_credit_available_0; // @[Router.scala 162:42]
  assign ingress_unit_2_from_1_io_out_credit_available_0_1 = output_unit_0_to_0_io_credit_available_1; // @[Router.scala 162:42]
  assign ingress_unit_2_from_1_io_out_credit_available_0_2 = output_unit_0_to_0_io_credit_available_2; // @[Router.scala 162:42]
  assign ingress_unit_2_from_1_io_out_credit_available_0_3 = output_unit_0_to_0_io_credit_available_3; // @[Router.scala 162:42]
  assign ingress_unit_2_from_1_io_salloc_req_0_ready = switch_allocator_io_req_2_0_ready; // @[Router.scala 165:23]
  assign ingress_unit_2_from_1_io_in_valid = auto_ingress_nodes_in_flit_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign ingress_unit_2_from_1_io_in_bits_head = auto_ingress_nodes_in_flit_bits_head; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign ingress_unit_2_from_1_io_in_bits_tail = auto_ingress_nodes_in_flit_bits_tail; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign ingress_unit_2_from_1_io_in_bits_payload = auto_ingress_nodes_in_flit_bits_payload; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign ingress_unit_2_from_1_io_in_bits_egress_id = auto_ingress_nodes_in_flit_bits_egress_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign output_unit_0_to_0_clock = clock;
  assign output_unit_0_to_0_reset = reset;
  assign output_unit_0_to_0_io_in_0_valid = switch_io_out_0_0_valid; // @[Router.scala 172:29]
  assign output_unit_0_to_0_io_in_0_bits_head = switch_io_out_0_0_bits_head; // @[Router.scala 172:29]
  assign output_unit_0_to_0_io_in_0_bits_tail = switch_io_out_0_0_bits_tail; // @[Router.scala 172:29]
  assign output_unit_0_to_0_io_in_0_bits_payload = switch_io_out_0_0_bits_payload; // @[Router.scala 172:29]
  assign output_unit_0_to_0_io_in_0_bits_flow_ingress_node = switch_io_out_0_0_bits_flow_ingress_node; // @[Router.scala 172:29]
  assign output_unit_0_to_0_io_in_0_bits_flow_egress_node = switch_io_out_0_0_bits_flow_egress_node; // @[Router.scala 172:29]
  assign output_unit_0_to_0_io_in_0_bits_virt_channel_id = switch_io_out_0_0_bits_virt_channel_id; // @[Router.scala 172:29]
  assign output_unit_0_to_0_io_allocs_0_alloc = vc_allocator_io_out_allocs_0_0_alloc; // @[Router.scala 157:33]
  assign output_unit_0_to_0_io_allocs_1_alloc = vc_allocator_io_out_allocs_0_1_alloc; // @[Router.scala 157:33]
  assign output_unit_0_to_0_io_allocs_2_alloc = vc_allocator_io_out_allocs_0_2_alloc; // @[Router.scala 157:33]
  assign output_unit_0_to_0_io_allocs_3_alloc = vc_allocator_io_out_allocs_0_3_alloc; // @[Router.scala 157:33]
  assign output_unit_0_to_0_io_credit_alloc_0_alloc = switch_allocator_io_credit_alloc_0_0_alloc; // @[Router.scala 167:39]
  assign output_unit_0_to_0_io_credit_alloc_1_alloc = switch_allocator_io_credit_alloc_0_1_alloc; // @[Router.scala 167:39]
  assign output_unit_0_to_0_io_credit_alloc_2_alloc = switch_allocator_io_credit_alloc_0_2_alloc; // @[Router.scala 167:39]
  assign output_unit_0_to_0_io_credit_alloc_3_alloc = switch_allocator_io_credit_alloc_0_3_alloc; // @[Router.scala 167:39]
  assign output_unit_0_to_0_io_out_credit_return = auto_source_nodes_out_0_credit_return; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign output_unit_0_to_0_io_out_vc_free = auto_source_nodes_out_0_vc_free; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign output_unit_1_to_2_clock = clock;
  assign output_unit_1_to_2_reset = reset;
  assign output_unit_1_to_2_io_in_0_valid = switch_io_out_1_0_valid; // @[Router.scala 172:29]
  assign output_unit_1_to_2_io_in_0_bits_head = switch_io_out_1_0_bits_head; // @[Router.scala 172:29]
  assign output_unit_1_to_2_io_in_0_bits_tail = switch_io_out_1_0_bits_tail; // @[Router.scala 172:29]
  assign output_unit_1_to_2_io_in_0_bits_payload = switch_io_out_1_0_bits_payload; // @[Router.scala 172:29]
  assign output_unit_1_to_2_io_in_0_bits_flow_ingress_node = switch_io_out_1_0_bits_flow_ingress_node; // @[Router.scala 172:29]
  assign output_unit_1_to_2_io_in_0_bits_flow_egress_node = switch_io_out_1_0_bits_flow_egress_node; // @[Router.scala 172:29]
  assign output_unit_1_to_2_io_in_0_bits_virt_channel_id = switch_io_out_1_0_bits_virt_channel_id; // @[Router.scala 172:29]
  assign output_unit_1_to_2_io_allocs_0_alloc = vc_allocator_io_out_allocs_1_0_alloc; // @[Router.scala 157:33]
  assign output_unit_1_to_2_io_allocs_1_alloc = vc_allocator_io_out_allocs_1_1_alloc; // @[Router.scala 157:33]
  assign output_unit_1_to_2_io_allocs_2_alloc = vc_allocator_io_out_allocs_1_2_alloc; // @[Router.scala 157:33]
  assign output_unit_1_to_2_io_allocs_3_alloc = vc_allocator_io_out_allocs_1_3_alloc; // @[Router.scala 157:33]
  assign output_unit_1_to_2_io_credit_alloc_0_alloc = switch_allocator_io_credit_alloc_1_0_alloc; // @[Router.scala 167:39]
  assign output_unit_1_to_2_io_credit_alloc_1_alloc = switch_allocator_io_credit_alloc_1_1_alloc; // @[Router.scala 167:39]
  assign output_unit_1_to_2_io_credit_alloc_2_alloc = switch_allocator_io_credit_alloc_1_2_alloc; // @[Router.scala 167:39]
  assign output_unit_1_to_2_io_credit_alloc_3_alloc = switch_allocator_io_credit_alloc_1_3_alloc; // @[Router.scala 167:39]
  assign output_unit_1_to_2_io_out_credit_return = auto_source_nodes_out_1_credit_return; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign output_unit_1_to_2_io_out_vc_free = auto_source_nodes_out_1_vc_free; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign egress_unit_2_to_1_clock = clock;
  assign egress_unit_2_to_1_reset = reset;
  assign egress_unit_2_to_1_io_in_0_valid = switch_io_out_2_0_valid; // @[Router.scala 172:29]
  assign egress_unit_2_to_1_io_in_0_bits_head = switch_io_out_2_0_bits_head; // @[Router.scala 172:29]
  assign egress_unit_2_to_1_io_in_0_bits_tail = switch_io_out_2_0_bits_tail; // @[Router.scala 172:29]
  assign egress_unit_2_to_1_io_in_0_bits_payload = switch_io_out_2_0_bits_payload; // @[Router.scala 172:29]
  assign egress_unit_2_to_1_io_in_0_bits_flow_ingress_node = switch_io_out_2_0_bits_flow_ingress_node; // @[Router.scala 172:29]
  assign egress_unit_2_to_1_io_allocs_0_alloc = vc_allocator_io_out_allocs_2_0_alloc; // @[Router.scala 157:33]
  assign egress_unit_2_to_1_io_credit_alloc_0_alloc = switch_allocator_io_credit_alloc_2_0_alloc; // @[Router.scala 167:39]
  assign egress_unit_2_to_1_io_credit_alloc_0_tail = switch_allocator_io_credit_alloc_2_0_tail; // @[Router.scala 167:39]
  assign switch_clock = clock;
  assign switch_reset = reset;
  assign switch_io_in_2_0_valid = ingress_unit_2_from_1_io_out_0_valid; // @[Router.scala 170:23]
  assign switch_io_in_2_0_bits_flit_head = ingress_unit_2_from_1_io_out_0_bits_flit_head; // @[Router.scala 170:23]
  assign switch_io_in_2_0_bits_flit_tail = ingress_unit_2_from_1_io_out_0_bits_flit_tail; // @[Router.scala 170:23]
  assign switch_io_in_2_0_bits_flit_payload = ingress_unit_2_from_1_io_out_0_bits_flit_payload; // @[Router.scala 170:23]
  assign switch_io_in_2_0_bits_flit_flow_ingress_node = ingress_unit_2_from_1_io_out_0_bits_flit_flow_ingress_node; // @[Router.scala 170:23]
  assign switch_io_in_2_0_bits_flit_flow_egress_node = ingress_unit_2_from_1_io_out_0_bits_flit_flow_egress_node; // @[Router.scala 170:23]
  assign switch_io_in_2_0_bits_out_virt_channel = ingress_unit_2_from_1_io_out_0_bits_out_virt_channel; // @[Router.scala 170:23]
  assign switch_io_in_1_0_valid = input_unit_1_from_2_io_out_0_valid; // @[Router.scala 170:23]
  assign switch_io_in_1_0_bits_flit_head = input_unit_1_from_2_io_out_0_bits_flit_head; // @[Router.scala 170:23]
  assign switch_io_in_1_0_bits_flit_tail = input_unit_1_from_2_io_out_0_bits_flit_tail; // @[Router.scala 170:23]
  assign switch_io_in_1_0_bits_flit_payload = input_unit_1_from_2_io_out_0_bits_flit_payload; // @[Router.scala 170:23]
  assign switch_io_in_1_0_bits_flit_flow_ingress_node = input_unit_1_from_2_io_out_0_bits_flit_flow_ingress_node; // @[Router.scala 170:23]
  assign switch_io_in_1_0_bits_flit_flow_egress_node = input_unit_1_from_2_io_out_0_bits_flit_flow_egress_node; // @[Router.scala 170:23]
  assign switch_io_in_1_0_bits_out_virt_channel = input_unit_1_from_2_io_out_0_bits_out_virt_channel; // @[Router.scala 170:23]
  assign switch_io_in_0_0_valid = input_unit_0_from_0_io_out_0_valid; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_head = input_unit_0_from_0_io_out_0_bits_flit_head; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_tail = input_unit_0_from_0_io_out_0_bits_flit_tail; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_payload = input_unit_0_from_0_io_out_0_bits_flit_payload; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_flow_ingress_node = input_unit_0_from_0_io_out_0_bits_flit_flow_ingress_node; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_flow_egress_node = input_unit_0_from_0_io_out_0_bits_flit_flow_egress_node; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_out_virt_channel = input_unit_0_from_0_io_out_0_bits_out_virt_channel; // @[Router.scala 170:23]
  assign switch_io_sel_2_0_2_0 = switch_io_sel_REG_2_0_2_0; // @[Router.scala 173:19]
  assign switch_io_sel_2_0_1_0 = switch_io_sel_REG_2_0_1_0; // @[Router.scala 173:19]
  assign switch_io_sel_2_0_0_0 = switch_io_sel_REG_2_0_0_0; // @[Router.scala 173:19]
  assign switch_io_sel_1_0_2_0 = switch_io_sel_REG_1_0_2_0; // @[Router.scala 173:19]
  assign switch_io_sel_1_0_1_0 = switch_io_sel_REG_1_0_1_0; // @[Router.scala 173:19]
  assign switch_io_sel_1_0_0_0 = switch_io_sel_REG_1_0_0_0; // @[Router.scala 173:19]
  assign switch_io_sel_0_0_2_0 = switch_io_sel_REG_0_0_2_0; // @[Router.scala 173:19]
  assign switch_io_sel_0_0_1_0 = switch_io_sel_REG_0_0_1_0; // @[Router.scala 173:19]
  assign switch_io_sel_0_0_0_0 = switch_io_sel_REG_0_0_0_0; // @[Router.scala 173:19]
  assign switch_allocator_clock = clock;
  assign switch_allocator_reset = reset;
  assign switch_allocator_io_req_2_0_valid = ingress_unit_2_from_1_io_salloc_req_0_valid; // @[Router.scala 165:23]
  assign switch_allocator_io_req_2_0_bits_vc_sel_2_0 = ingress_unit_2_from_1_io_salloc_req_0_bits_vc_sel_2_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_2_0_bits_vc_sel_1_0 = ingress_unit_2_from_1_io_salloc_req_0_bits_vc_sel_1_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_2_0_bits_vc_sel_1_1 = ingress_unit_2_from_1_io_salloc_req_0_bits_vc_sel_1_1; // @[Router.scala 165:23]
  assign switch_allocator_io_req_2_0_bits_vc_sel_1_2 = ingress_unit_2_from_1_io_salloc_req_0_bits_vc_sel_1_2; // @[Router.scala 165:23]
  assign switch_allocator_io_req_2_0_bits_vc_sel_1_3 = ingress_unit_2_from_1_io_salloc_req_0_bits_vc_sel_1_3; // @[Router.scala 165:23]
  assign switch_allocator_io_req_2_0_bits_vc_sel_0_0 = ingress_unit_2_from_1_io_salloc_req_0_bits_vc_sel_0_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_2_0_bits_vc_sel_0_1 = ingress_unit_2_from_1_io_salloc_req_0_bits_vc_sel_0_1; // @[Router.scala 165:23]
  assign switch_allocator_io_req_2_0_bits_vc_sel_0_2 = ingress_unit_2_from_1_io_salloc_req_0_bits_vc_sel_0_2; // @[Router.scala 165:23]
  assign switch_allocator_io_req_2_0_bits_vc_sel_0_3 = ingress_unit_2_from_1_io_salloc_req_0_bits_vc_sel_0_3; // @[Router.scala 165:23]
  assign switch_allocator_io_req_2_0_bits_tail = ingress_unit_2_from_1_io_salloc_req_0_bits_tail; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_valid = input_unit_1_from_2_io_salloc_req_0_valid; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_vc_sel_2_0 = input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_2_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_vc_sel_1_0 = input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_1_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_vc_sel_1_1 = input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_1_1; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_vc_sel_1_2 = input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_1_2; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_vc_sel_1_3 = input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_1_3; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_vc_sel_0_0 = input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_0_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_vc_sel_0_1 = input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_0_1; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_vc_sel_0_2 = input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_0_2; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_vc_sel_0_3 = input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_0_3; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_tail = input_unit_1_from_2_io_salloc_req_0_bits_tail; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_valid = input_unit_0_from_0_io_salloc_req_0_valid; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_2_0 = input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_2_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_1_0 = input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_1_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_1_1 = input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_1_1; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_1_2 = input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_1_2; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_1_3 = input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_1_3; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_0_0 = input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_0_1 = input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_1; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_0_2 = input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_2; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_0_3 = input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_3; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_tail = input_unit_0_from_0_io_salloc_req_0_bits_tail; // @[Router.scala 165:23]
  assign vc_allocator_clock = clock;
  assign vc_allocator_reset = reset;
  assign vc_allocator_io_req_2_valid = ingress_unit_2_from_1_io_vcalloc_req_valid; // @[Router.scala 151:23]
  assign vc_allocator_io_req_2_bits_vc_sel_2_0 = ingress_unit_2_from_1_io_vcalloc_req_bits_vc_sel_2_0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_2_bits_vc_sel_1_0 = ingress_unit_2_from_1_io_vcalloc_req_bits_vc_sel_1_0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_2_bits_vc_sel_1_1 = ingress_unit_2_from_1_io_vcalloc_req_bits_vc_sel_1_1; // @[Router.scala 151:23]
  assign vc_allocator_io_req_2_bits_vc_sel_1_2 = ingress_unit_2_from_1_io_vcalloc_req_bits_vc_sel_1_2; // @[Router.scala 151:23]
  assign vc_allocator_io_req_2_bits_vc_sel_1_3 = ingress_unit_2_from_1_io_vcalloc_req_bits_vc_sel_1_3; // @[Router.scala 151:23]
  assign vc_allocator_io_req_2_bits_vc_sel_0_0 = ingress_unit_2_from_1_io_vcalloc_req_bits_vc_sel_0_0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_2_bits_vc_sel_0_1 = ingress_unit_2_from_1_io_vcalloc_req_bits_vc_sel_0_1; // @[Router.scala 151:23]
  assign vc_allocator_io_req_2_bits_vc_sel_0_2 = ingress_unit_2_from_1_io_vcalloc_req_bits_vc_sel_0_2; // @[Router.scala 151:23]
  assign vc_allocator_io_req_2_bits_vc_sel_0_3 = ingress_unit_2_from_1_io_vcalloc_req_bits_vc_sel_0_3; // @[Router.scala 151:23]
  assign vc_allocator_io_req_1_valid = input_unit_1_from_2_io_vcalloc_req_valid; // @[Router.scala 151:23]
  assign vc_allocator_io_req_1_bits_vc_sel_2_0 = input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_2_0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_1_bits_vc_sel_1_0 = input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_1_0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_1_bits_vc_sel_1_1 = input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_1_1; // @[Router.scala 151:23]
  assign vc_allocator_io_req_1_bits_vc_sel_1_2 = input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_1_2; // @[Router.scala 151:23]
  assign vc_allocator_io_req_1_bits_vc_sel_1_3 = input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_1_3; // @[Router.scala 151:23]
  assign vc_allocator_io_req_1_bits_vc_sel_0_0 = input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_0_0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_1_bits_vc_sel_0_1 = input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_0_1; // @[Router.scala 151:23]
  assign vc_allocator_io_req_1_bits_vc_sel_0_2 = input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_0_2; // @[Router.scala 151:23]
  assign vc_allocator_io_req_1_bits_vc_sel_0_3 = input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_0_3; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_valid = input_unit_0_from_0_io_vcalloc_req_valid; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_2_0 = input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_2_0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_1_0 = input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_1_0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_1_1 = input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_1_1; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_1_2 = input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_1_2; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_1_3 = input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_1_3; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_0_0 = input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_0_1 = input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_1; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_0_2 = input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_2; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_0_3 = input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_3; // @[Router.scala 151:23]
  assign vc_allocator_io_channel_status_2_0_occupied = egress_unit_2_to_1_io_channel_status_0_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_1_0_occupied = output_unit_1_to_2_io_channel_status_0_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_1_1_occupied = output_unit_1_to_2_io_channel_status_1_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_1_2_occupied = output_unit_1_to_2_io_channel_status_2_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_1_3_occupied = output_unit_1_to_2_io_channel_status_3_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_0_0_occupied = output_unit_0_to_0_io_channel_status_0_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_0_1_occupied = output_unit_0_to_0_io_channel_status_1_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_0_2_occupied = output_unit_0_to_0_io_channel_status_2_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_0_3_occupied = output_unit_0_to_0_io_channel_status_3_occupied; // @[Router.scala 159:23]
  assign route_computer_io_req_2_bits_flow_ingress_node = ingress_unit_2_from_1_io_router_req_bits_flow_ingress_node; // @[Router.scala 146:23]
  assign route_computer_io_req_2_bits_flow_egress_node = ingress_unit_2_from_1_io_router_req_bits_flow_egress_node; // @[Router.scala 146:23]
  assign route_computer_io_req_1_bits_src_virt_id = input_unit_1_from_2_io_router_req_bits_src_virt_id; // @[Router.scala 146:23]
  assign route_computer_io_req_1_bits_flow_ingress_node = input_unit_1_from_2_io_router_req_bits_flow_ingress_node; // @[Router.scala 146:23]
  assign route_computer_io_req_1_bits_flow_egress_node = input_unit_1_from_2_io_router_req_bits_flow_egress_node; // @[Router.scala 146:23]
  assign route_computer_io_req_0_bits_src_virt_id = input_unit_0_from_0_io_router_req_bits_src_virt_id; // @[Router.scala 146:23]
  assign route_computer_io_req_0_bits_flow_ingress_node = input_unit_0_from_0_io_router_req_bits_flow_ingress_node; // @[Router.scala 146:23]
  assign route_computer_io_req_0_bits_flow_egress_node = input_unit_0_from_0_io_router_req_bits_flow_egress_node; // @[Router.scala 146:23]
  always @(posedge clock) begin
    switch_io_sel_REG_2_0_2_0 <= switch_allocator_io_switch_sel_2_0_2_0; // @[Router.scala 176:14]
    switch_io_sel_REG_2_0_1_0 <= switch_allocator_io_switch_sel_2_0_1_0; // @[Router.scala 176:14]
    switch_io_sel_REG_2_0_0_0 <= switch_allocator_io_switch_sel_2_0_0_0; // @[Router.scala 176:14]
    switch_io_sel_REG_1_0_2_0 <= switch_allocator_io_switch_sel_1_0_2_0; // @[Router.scala 176:14]
    switch_io_sel_REG_1_0_1_0 <= switch_allocator_io_switch_sel_1_0_1_0; // @[Router.scala 176:14]
    switch_io_sel_REG_1_0_0_0 <= switch_allocator_io_switch_sel_1_0_0_0; // @[Router.scala 176:14]
    switch_io_sel_REG_0_0_2_0 <= switch_allocator_io_switch_sel_0_0_2_0; // @[Router.scala 176:14]
    switch_io_sel_REG_0_0_1_0 <= switch_allocator_io_switch_sel_0_0_1_0; // @[Router.scala 176:14]
    switch_io_sel_REG_0_0_0_0 <= switch_allocator_io_switch_sel_0_0_0_0; // @[Router.scala 176:14]
    if (reset) begin // @[Router.scala 193:28]
      debug_tsc <= 64'h0; // @[Router.scala 193:28]
    end else begin
      debug_tsc <= _debug_tsc_T_1; // @[Router.scala 194:15]
    end
    if (reset) begin // @[Router.scala 195:31]
      debug_sample <= 64'h0; // @[Router.scala 195:31]
    end else if (debug_sample == _GEN_6) begin // @[Router.scala 198:47]
      debug_sample <= 64'h0; // @[Router.scala 198:62]
    end else begin
      debug_sample <= _debug_sample_T_1; // @[Router.scala 196:18]
    end
    if (reset) begin // @[Router.scala 201:29]
      util_ctr <= 64'h0; // @[Router.scala 201:29]
    end else begin
      util_ctr <= _util_ctr_T_1; // @[Router.scala 203:16]
    end
    if (reset) begin // @[Router.scala 202:26]
      fired <= 1'h0; // @[Router.scala 202:26]
    end else if (plusarg_reader_out != 20'h0 & _T_2 & fired) begin // @[Router.scala 205:81]
      fired <= auto_dest_nodes_in_0_flit_0_valid; // @[Router.scala 208:15]
    end else begin
      fired <= fired | auto_dest_nodes_in_0_flit_0_valid; // @[Router.scala 204:13]
    end
    if (reset) begin // @[Router.scala 201:29]
      util_ctr_1 <= 64'h0; // @[Router.scala 201:29]
    end else begin
      util_ctr_1 <= _util_ctr_T_3; // @[Router.scala 203:16]
    end
    if (reset) begin // @[Router.scala 202:26]
      fired_1 <= 1'h0; // @[Router.scala 202:26]
    end else if (plusarg_reader_out != 20'h0 & _T_2 & fired_1) begin // @[Router.scala 205:81]
      fired_1 <= auto_dest_nodes_in_1_flit_0_valid; // @[Router.scala 208:15]
    end else begin
      fired_1 <= fired_1 | auto_dest_nodes_in_1_flit_0_valid; // @[Router.scala 204:13]
    end
    if (reset) begin // @[Router.scala 201:29]
      util_ctr_2 <= 64'h0; // @[Router.scala 201:29]
    end else begin
      util_ctr_2 <= _util_ctr_T_5; // @[Router.scala 203:16]
    end
    if (reset) begin // @[Router.scala 202:26]
      fired_2 <= 1'h0; // @[Router.scala 202:26]
    end else if (plusarg_reader_out != 20'h0 & _T_2 & fired_2) begin // @[Router.scala 205:81]
      fired_2 <= _T_19; // @[Router.scala 208:15]
    end else begin
      fired_2 <= fired_2 | _T_19; // @[Router.scala 204:13]
    end
    if (reset) begin // @[Router.scala 201:29]
      util_ctr_3 <= 64'h0; // @[Router.scala 201:29]
    end else begin
      util_ctr_3 <= _util_ctr_T_7; // @[Router.scala 203:16]
    end
    if (reset) begin // @[Router.scala 202:26]
      fired_3 <= 1'h0; // @[Router.scala 202:26]
    end else if (plusarg_reader_out != 20'h0 & _T_2 & fired_3) begin // @[Router.scala 205:81]
      fired_3 <= x1_2_flit_valid; // @[Router.scala 208:15]
    end else begin
      fired_3 <= fired_3 | x1_2_flit_valid; // @[Router.scala 204:13]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8 & ~reset) begin
          $fwrite(32'h80000002,"nocsample %d 0 1 %d\n",debug_tsc,util_ctr); // @[Router.scala 207:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_16 & ~reset) begin
          $fwrite(32'h80000002,"nocsample %d 2 1 %d\n",debug_tsc,util_ctr_1); // @[Router.scala 207:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_25 & ~reset) begin
          $fwrite(32'h80000002,"nocsample %d i1 1 %d\n",debug_tsc,util_ctr_2); // @[Router.scala 207:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_34 & ~reset) begin
          $fwrite(32'h80000002,"nocsample %d 1 e1 %d\n",debug_tsc,util_ctr_3); // @[Router.scala 207:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  switch_io_sel_REG_2_0_2_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  switch_io_sel_REG_2_0_1_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  switch_io_sel_REG_2_0_0_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  switch_io_sel_REG_1_0_2_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  switch_io_sel_REG_1_0_1_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  switch_io_sel_REG_1_0_0_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  switch_io_sel_REG_0_0_2_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  switch_io_sel_REG_0_0_1_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  switch_io_sel_REG_0_0_0_0 = _RAND_8[0:0];
  _RAND_9 = {2{`RANDOM}};
  debug_tsc = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  debug_sample = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  util_ctr = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  fired = _RAND_12[0:0];
  _RAND_13 = {2{`RANDOM}};
  util_ctr_1 = _RAND_13[63:0];
  _RAND_14 = {1{`RANDOM}};
  fired_1 = _RAND_14[0:0];
  _RAND_15 = {2{`RANDOM}};
  util_ctr_2 = _RAND_15[63:0];
  _RAND_16 = {1{`RANDOM}};
  fired_2 = _RAND_16[0:0];
  _RAND_17 = {2{`RANDOM}};
  util_ctr_3 = _RAND_17[63:0];
  _RAND_18 = {1{`RANDOM}};
  fired_3 = _RAND_18[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ClockSinkDomain_1(
  output [1:0]  auto_routers_debug_out_va_stall_0,
  output [1:0]  auto_routers_debug_out_va_stall_1,
  output [1:0]  auto_routers_debug_out_sa_stall_0,
  output [1:0]  auto_routers_debug_out_sa_stall_1,
  output        auto_routers_egress_nodes_out_flit_valid,
  output        auto_routers_egress_nodes_out_flit_bits_head,
  output        auto_routers_egress_nodes_out_flit_bits_tail,
  output [63:0] auto_routers_egress_nodes_out_flit_bits_payload,
  output [1:0]  auto_routers_egress_nodes_out_flit_bits_ingress_id,
  output        auto_routers_ingress_nodes_in_flit_ready,
  input         auto_routers_ingress_nodes_in_flit_valid,
  input         auto_routers_ingress_nodes_in_flit_bits_head,
  input         auto_routers_ingress_nodes_in_flit_bits_tail,
  input  [63:0] auto_routers_ingress_nodes_in_flit_bits_payload,
  input  [1:0]  auto_routers_ingress_nodes_in_flit_bits_egress_id,
  output        auto_routers_source_nodes_out_1_flit_0_valid,
  output        auto_routers_source_nodes_out_1_flit_0_bits_head,
  output        auto_routers_source_nodes_out_1_flit_0_bits_tail,
  output [63:0] auto_routers_source_nodes_out_1_flit_0_bits_payload,
  output [1:0]  auto_routers_source_nodes_out_1_flit_0_bits_flow_ingress_node,
  output [1:0]  auto_routers_source_nodes_out_1_flit_0_bits_flow_egress_node,
  output [1:0]  auto_routers_source_nodes_out_1_flit_0_bits_virt_channel_id,
  input  [3:0]  auto_routers_source_nodes_out_1_credit_return,
  input  [3:0]  auto_routers_source_nodes_out_1_vc_free,
  output        auto_routers_source_nodes_out_0_flit_0_valid,
  output        auto_routers_source_nodes_out_0_flit_0_bits_head,
  output        auto_routers_source_nodes_out_0_flit_0_bits_tail,
  output [63:0] auto_routers_source_nodes_out_0_flit_0_bits_payload,
  output [1:0]  auto_routers_source_nodes_out_0_flit_0_bits_flow_ingress_node,
  output [1:0]  auto_routers_source_nodes_out_0_flit_0_bits_flow_egress_node,
  output [1:0]  auto_routers_source_nodes_out_0_flit_0_bits_virt_channel_id,
  input  [3:0]  auto_routers_source_nodes_out_0_credit_return,
  input  [3:0]  auto_routers_source_nodes_out_0_vc_free,
  input         auto_routers_dest_nodes_in_1_flit_0_valid,
  input         auto_routers_dest_nodes_in_1_flit_0_bits_head,
  input         auto_routers_dest_nodes_in_1_flit_0_bits_tail,
  input  [63:0] auto_routers_dest_nodes_in_1_flit_0_bits_payload,
  input  [1:0]  auto_routers_dest_nodes_in_1_flit_0_bits_flow_ingress_node,
  input  [1:0]  auto_routers_dest_nodes_in_1_flit_0_bits_flow_egress_node,
  input  [1:0]  auto_routers_dest_nodes_in_1_flit_0_bits_virt_channel_id,
  output [3:0]  auto_routers_dest_nodes_in_1_credit_return,
  output [3:0]  auto_routers_dest_nodes_in_1_vc_free,
  input         auto_routers_dest_nodes_in_0_flit_0_valid,
  input         auto_routers_dest_nodes_in_0_flit_0_bits_head,
  input         auto_routers_dest_nodes_in_0_flit_0_bits_tail,
  input  [63:0] auto_routers_dest_nodes_in_0_flit_0_bits_payload,
  input  [1:0]  auto_routers_dest_nodes_in_0_flit_0_bits_flow_ingress_node,
  input  [1:0]  auto_routers_dest_nodes_in_0_flit_0_bits_flow_egress_node,
  input  [1:0]  auto_routers_dest_nodes_in_0_flit_0_bits_virt_channel_id,
  output [3:0]  auto_routers_dest_nodes_in_0_credit_return,
  output [3:0]  auto_routers_dest_nodes_in_0_vc_free,
  input         auto_clock_in_clock,
  input         auto_clock_in_reset
);
  wire  routers_clock; // @[NoC.scala 64:22]
  wire  routers_reset; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_debug_out_va_stall_0; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_debug_out_va_stall_1; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_debug_out_sa_stall_0; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_debug_out_sa_stall_1; // @[NoC.scala 64:22]
  wire  routers_auto_egress_nodes_out_flit_valid; // @[NoC.scala 64:22]
  wire  routers_auto_egress_nodes_out_flit_bits_head; // @[NoC.scala 64:22]
  wire  routers_auto_egress_nodes_out_flit_bits_tail; // @[NoC.scala 64:22]
  wire [63:0] routers_auto_egress_nodes_out_flit_bits_payload; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_egress_nodes_out_flit_bits_ingress_id; // @[NoC.scala 64:22]
  wire  routers_auto_ingress_nodes_in_flit_ready; // @[NoC.scala 64:22]
  wire  routers_auto_ingress_nodes_in_flit_valid; // @[NoC.scala 64:22]
  wire  routers_auto_ingress_nodes_in_flit_bits_head; // @[NoC.scala 64:22]
  wire  routers_auto_ingress_nodes_in_flit_bits_tail; // @[NoC.scala 64:22]
  wire [63:0] routers_auto_ingress_nodes_in_flit_bits_payload; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_ingress_nodes_in_flit_bits_egress_id; // @[NoC.scala 64:22]
  wire  routers_auto_source_nodes_out_1_flit_0_valid; // @[NoC.scala 64:22]
  wire  routers_auto_source_nodes_out_1_flit_0_bits_head; // @[NoC.scala 64:22]
  wire  routers_auto_source_nodes_out_1_flit_0_bits_tail; // @[NoC.scala 64:22]
  wire [63:0] routers_auto_source_nodes_out_1_flit_0_bits_payload; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_source_nodes_out_1_flit_0_bits_flow_ingress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_source_nodes_out_1_flit_0_bits_flow_egress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_source_nodes_out_1_flit_0_bits_virt_channel_id; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_source_nodes_out_1_credit_return; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_source_nodes_out_1_vc_free; // @[NoC.scala 64:22]
  wire  routers_auto_source_nodes_out_0_flit_0_valid; // @[NoC.scala 64:22]
  wire  routers_auto_source_nodes_out_0_flit_0_bits_head; // @[NoC.scala 64:22]
  wire  routers_auto_source_nodes_out_0_flit_0_bits_tail; // @[NoC.scala 64:22]
  wire [63:0] routers_auto_source_nodes_out_0_flit_0_bits_payload; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_source_nodes_out_0_flit_0_bits_flow_ingress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_source_nodes_out_0_flit_0_bits_flow_egress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_source_nodes_out_0_flit_0_bits_virt_channel_id; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_source_nodes_out_0_credit_return; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_source_nodes_out_0_vc_free; // @[NoC.scala 64:22]
  wire  routers_auto_dest_nodes_in_1_flit_0_valid; // @[NoC.scala 64:22]
  wire  routers_auto_dest_nodes_in_1_flit_0_bits_head; // @[NoC.scala 64:22]
  wire  routers_auto_dest_nodes_in_1_flit_0_bits_tail; // @[NoC.scala 64:22]
  wire [63:0] routers_auto_dest_nodes_in_1_flit_0_bits_payload; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_dest_nodes_in_1_flit_0_bits_flow_ingress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_dest_nodes_in_1_flit_0_bits_flow_egress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_dest_nodes_in_1_flit_0_bits_virt_channel_id; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_dest_nodes_in_1_credit_return; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_dest_nodes_in_1_vc_free; // @[NoC.scala 64:22]
  wire  routers_auto_dest_nodes_in_0_flit_0_valid; // @[NoC.scala 64:22]
  wire  routers_auto_dest_nodes_in_0_flit_0_bits_head; // @[NoC.scala 64:22]
  wire  routers_auto_dest_nodes_in_0_flit_0_bits_tail; // @[NoC.scala 64:22]
  wire [63:0] routers_auto_dest_nodes_in_0_flit_0_bits_payload; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_dest_nodes_in_0_flit_0_bits_flow_ingress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_dest_nodes_in_0_flit_0_bits_flow_egress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_dest_nodes_in_0_flit_0_bits_virt_channel_id; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_dest_nodes_in_0_credit_return; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_dest_nodes_in_0_vc_free; // @[NoC.scala 64:22]
  Router_1 routers ( // @[NoC.scala 64:22]
    .clock(routers_clock),
    .reset(routers_reset),
    .auto_debug_out_va_stall_0(routers_auto_debug_out_va_stall_0),
    .auto_debug_out_va_stall_1(routers_auto_debug_out_va_stall_1),
    .auto_debug_out_sa_stall_0(routers_auto_debug_out_sa_stall_0),
    .auto_debug_out_sa_stall_1(routers_auto_debug_out_sa_stall_1),
    .auto_egress_nodes_out_flit_valid(routers_auto_egress_nodes_out_flit_valid),
    .auto_egress_nodes_out_flit_bits_head(routers_auto_egress_nodes_out_flit_bits_head),
    .auto_egress_nodes_out_flit_bits_tail(routers_auto_egress_nodes_out_flit_bits_tail),
    .auto_egress_nodes_out_flit_bits_payload(routers_auto_egress_nodes_out_flit_bits_payload),
    .auto_egress_nodes_out_flit_bits_ingress_id(routers_auto_egress_nodes_out_flit_bits_ingress_id),
    .auto_ingress_nodes_in_flit_ready(routers_auto_ingress_nodes_in_flit_ready),
    .auto_ingress_nodes_in_flit_valid(routers_auto_ingress_nodes_in_flit_valid),
    .auto_ingress_nodes_in_flit_bits_head(routers_auto_ingress_nodes_in_flit_bits_head),
    .auto_ingress_nodes_in_flit_bits_tail(routers_auto_ingress_nodes_in_flit_bits_tail),
    .auto_ingress_nodes_in_flit_bits_payload(routers_auto_ingress_nodes_in_flit_bits_payload),
    .auto_ingress_nodes_in_flit_bits_egress_id(routers_auto_ingress_nodes_in_flit_bits_egress_id),
    .auto_source_nodes_out_1_flit_0_valid(routers_auto_source_nodes_out_1_flit_0_valid),
    .auto_source_nodes_out_1_flit_0_bits_head(routers_auto_source_nodes_out_1_flit_0_bits_head),
    .auto_source_nodes_out_1_flit_0_bits_tail(routers_auto_source_nodes_out_1_flit_0_bits_tail),
    .auto_source_nodes_out_1_flit_0_bits_payload(routers_auto_source_nodes_out_1_flit_0_bits_payload),
    .auto_source_nodes_out_1_flit_0_bits_flow_ingress_node(routers_auto_source_nodes_out_1_flit_0_bits_flow_ingress_node
      ),
    .auto_source_nodes_out_1_flit_0_bits_flow_egress_node(routers_auto_source_nodes_out_1_flit_0_bits_flow_egress_node),
    .auto_source_nodes_out_1_flit_0_bits_virt_channel_id(routers_auto_source_nodes_out_1_flit_0_bits_virt_channel_id),
    .auto_source_nodes_out_1_credit_return(routers_auto_source_nodes_out_1_credit_return),
    .auto_source_nodes_out_1_vc_free(routers_auto_source_nodes_out_1_vc_free),
    .auto_source_nodes_out_0_flit_0_valid(routers_auto_source_nodes_out_0_flit_0_valid),
    .auto_source_nodes_out_0_flit_0_bits_head(routers_auto_source_nodes_out_0_flit_0_bits_head),
    .auto_source_nodes_out_0_flit_0_bits_tail(routers_auto_source_nodes_out_0_flit_0_bits_tail),
    .auto_source_nodes_out_0_flit_0_bits_payload(routers_auto_source_nodes_out_0_flit_0_bits_payload),
    .auto_source_nodes_out_0_flit_0_bits_flow_ingress_node(routers_auto_source_nodes_out_0_flit_0_bits_flow_ingress_node
      ),
    .auto_source_nodes_out_0_flit_0_bits_flow_egress_node(routers_auto_source_nodes_out_0_flit_0_bits_flow_egress_node),
    .auto_source_nodes_out_0_flit_0_bits_virt_channel_id(routers_auto_source_nodes_out_0_flit_0_bits_virt_channel_id),
    .auto_source_nodes_out_0_credit_return(routers_auto_source_nodes_out_0_credit_return),
    .auto_source_nodes_out_0_vc_free(routers_auto_source_nodes_out_0_vc_free),
    .auto_dest_nodes_in_1_flit_0_valid(routers_auto_dest_nodes_in_1_flit_0_valid),
    .auto_dest_nodes_in_1_flit_0_bits_head(routers_auto_dest_nodes_in_1_flit_0_bits_head),
    .auto_dest_nodes_in_1_flit_0_bits_tail(routers_auto_dest_nodes_in_1_flit_0_bits_tail),
    .auto_dest_nodes_in_1_flit_0_bits_payload(routers_auto_dest_nodes_in_1_flit_0_bits_payload),
    .auto_dest_nodes_in_1_flit_0_bits_flow_ingress_node(routers_auto_dest_nodes_in_1_flit_0_bits_flow_ingress_node),
    .auto_dest_nodes_in_1_flit_0_bits_flow_egress_node(routers_auto_dest_nodes_in_1_flit_0_bits_flow_egress_node),
    .auto_dest_nodes_in_1_flit_0_bits_virt_channel_id(routers_auto_dest_nodes_in_1_flit_0_bits_virt_channel_id),
    .auto_dest_nodes_in_1_credit_return(routers_auto_dest_nodes_in_1_credit_return),
    .auto_dest_nodes_in_1_vc_free(routers_auto_dest_nodes_in_1_vc_free),
    .auto_dest_nodes_in_0_flit_0_valid(routers_auto_dest_nodes_in_0_flit_0_valid),
    .auto_dest_nodes_in_0_flit_0_bits_head(routers_auto_dest_nodes_in_0_flit_0_bits_head),
    .auto_dest_nodes_in_0_flit_0_bits_tail(routers_auto_dest_nodes_in_0_flit_0_bits_tail),
    .auto_dest_nodes_in_0_flit_0_bits_payload(routers_auto_dest_nodes_in_0_flit_0_bits_payload),
    .auto_dest_nodes_in_0_flit_0_bits_flow_ingress_node(routers_auto_dest_nodes_in_0_flit_0_bits_flow_ingress_node),
    .auto_dest_nodes_in_0_flit_0_bits_flow_egress_node(routers_auto_dest_nodes_in_0_flit_0_bits_flow_egress_node),
    .auto_dest_nodes_in_0_flit_0_bits_virt_channel_id(routers_auto_dest_nodes_in_0_flit_0_bits_virt_channel_id),
    .auto_dest_nodes_in_0_credit_return(routers_auto_dest_nodes_in_0_credit_return),
    .auto_dest_nodes_in_0_vc_free(routers_auto_dest_nodes_in_0_vc_free)
  );
  assign auto_routers_debug_out_va_stall_0 = routers_auto_debug_out_va_stall_0; // @[LazyModule.scala 368:12]
  assign auto_routers_debug_out_va_stall_1 = routers_auto_debug_out_va_stall_1; // @[LazyModule.scala 368:12]
  assign auto_routers_debug_out_sa_stall_0 = routers_auto_debug_out_sa_stall_0; // @[LazyModule.scala 368:12]
  assign auto_routers_debug_out_sa_stall_1 = routers_auto_debug_out_sa_stall_1; // @[LazyModule.scala 368:12]
  assign auto_routers_egress_nodes_out_flit_valid = routers_auto_egress_nodes_out_flit_valid; // @[LazyModule.scala 368:12]
  assign auto_routers_egress_nodes_out_flit_bits_head = routers_auto_egress_nodes_out_flit_bits_head; // @[LazyModule.scala 368:12]
  assign auto_routers_egress_nodes_out_flit_bits_tail = routers_auto_egress_nodes_out_flit_bits_tail; // @[LazyModule.scala 368:12]
  assign auto_routers_egress_nodes_out_flit_bits_payload = routers_auto_egress_nodes_out_flit_bits_payload; // @[LazyModule.scala 368:12]
  assign auto_routers_egress_nodes_out_flit_bits_ingress_id = routers_auto_egress_nodes_out_flit_bits_ingress_id; // @[LazyModule.scala 368:12]
  assign auto_routers_ingress_nodes_in_flit_ready = routers_auto_ingress_nodes_in_flit_ready; // @[LazyModule.scala 366:16]
  assign auto_routers_source_nodes_out_1_flit_0_valid = routers_auto_source_nodes_out_1_flit_0_valid; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_1_flit_0_bits_head = routers_auto_source_nodes_out_1_flit_0_bits_head; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_1_flit_0_bits_tail = routers_auto_source_nodes_out_1_flit_0_bits_tail; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_1_flit_0_bits_payload = routers_auto_source_nodes_out_1_flit_0_bits_payload; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_1_flit_0_bits_flow_ingress_node =
    routers_auto_source_nodes_out_1_flit_0_bits_flow_ingress_node; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_1_flit_0_bits_flow_egress_node =
    routers_auto_source_nodes_out_1_flit_0_bits_flow_egress_node; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_1_flit_0_bits_virt_channel_id =
    routers_auto_source_nodes_out_1_flit_0_bits_virt_channel_id; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_0_flit_0_valid = routers_auto_source_nodes_out_0_flit_0_valid; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_0_flit_0_bits_head = routers_auto_source_nodes_out_0_flit_0_bits_head; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_0_flit_0_bits_tail = routers_auto_source_nodes_out_0_flit_0_bits_tail; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_0_flit_0_bits_payload = routers_auto_source_nodes_out_0_flit_0_bits_payload; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_0_flit_0_bits_flow_ingress_node =
    routers_auto_source_nodes_out_0_flit_0_bits_flow_ingress_node; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_0_flit_0_bits_flow_egress_node =
    routers_auto_source_nodes_out_0_flit_0_bits_flow_egress_node; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_0_flit_0_bits_virt_channel_id =
    routers_auto_source_nodes_out_0_flit_0_bits_virt_channel_id; // @[LazyModule.scala 368:12]
  assign auto_routers_dest_nodes_in_1_credit_return = routers_auto_dest_nodes_in_1_credit_return; // @[LazyModule.scala 366:16]
  assign auto_routers_dest_nodes_in_1_vc_free = routers_auto_dest_nodes_in_1_vc_free; // @[LazyModule.scala 366:16]
  assign auto_routers_dest_nodes_in_0_credit_return = routers_auto_dest_nodes_in_0_credit_return; // @[LazyModule.scala 366:16]
  assign auto_routers_dest_nodes_in_0_vc_free = routers_auto_dest_nodes_in_0_vc_free; // @[LazyModule.scala 366:16]
  assign routers_clock = auto_clock_in_clock; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign routers_reset = auto_clock_in_reset; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign routers_auto_ingress_nodes_in_flit_valid = auto_routers_ingress_nodes_in_flit_valid; // @[LazyModule.scala 366:16]
  assign routers_auto_ingress_nodes_in_flit_bits_head = auto_routers_ingress_nodes_in_flit_bits_head; // @[LazyModule.scala 366:16]
  assign routers_auto_ingress_nodes_in_flit_bits_tail = auto_routers_ingress_nodes_in_flit_bits_tail; // @[LazyModule.scala 366:16]
  assign routers_auto_ingress_nodes_in_flit_bits_payload = auto_routers_ingress_nodes_in_flit_bits_payload; // @[LazyModule.scala 366:16]
  assign routers_auto_ingress_nodes_in_flit_bits_egress_id = auto_routers_ingress_nodes_in_flit_bits_egress_id; // @[LazyModule.scala 366:16]
  assign routers_auto_source_nodes_out_1_credit_return = auto_routers_source_nodes_out_1_credit_return; // @[LazyModule.scala 368:12]
  assign routers_auto_source_nodes_out_1_vc_free = auto_routers_source_nodes_out_1_vc_free; // @[LazyModule.scala 368:12]
  assign routers_auto_source_nodes_out_0_credit_return = auto_routers_source_nodes_out_0_credit_return; // @[LazyModule.scala 368:12]
  assign routers_auto_source_nodes_out_0_vc_free = auto_routers_source_nodes_out_0_vc_free; // @[LazyModule.scala 368:12]
  assign routers_auto_dest_nodes_in_1_flit_0_valid = auto_routers_dest_nodes_in_1_flit_0_valid; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_1_flit_0_bits_head = auto_routers_dest_nodes_in_1_flit_0_bits_head; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_1_flit_0_bits_tail = auto_routers_dest_nodes_in_1_flit_0_bits_tail; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_1_flit_0_bits_payload = auto_routers_dest_nodes_in_1_flit_0_bits_payload; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_1_flit_0_bits_flow_ingress_node =
    auto_routers_dest_nodes_in_1_flit_0_bits_flow_ingress_node; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_1_flit_0_bits_flow_egress_node =
    auto_routers_dest_nodes_in_1_flit_0_bits_flow_egress_node; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_1_flit_0_bits_virt_channel_id =
    auto_routers_dest_nodes_in_1_flit_0_bits_virt_channel_id; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_0_flit_0_valid = auto_routers_dest_nodes_in_0_flit_0_valid; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_0_flit_0_bits_head = auto_routers_dest_nodes_in_0_flit_0_bits_head; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_0_flit_0_bits_tail = auto_routers_dest_nodes_in_0_flit_0_bits_tail; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_0_flit_0_bits_payload = auto_routers_dest_nodes_in_0_flit_0_bits_payload; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_0_flit_0_bits_flow_ingress_node =
    auto_routers_dest_nodes_in_0_flit_0_bits_flow_ingress_node; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_0_flit_0_bits_flow_egress_node =
    auto_routers_dest_nodes_in_0_flit_0_bits_flow_egress_node; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_0_flit_0_bits_virt_channel_id =
    auto_routers_dest_nodes_in_0_flit_0_bits_virt_channel_id; // @[LazyModule.scala 366:16]
endmodule
module NoCMonitor_4(
  input        clock,
  input        reset,
  input        io_in_flit_0_valid,
  input        io_in_flit_0_bits_head,
  input        io_in_flit_0_bits_tail,
  input  [1:0] io_in_flit_0_bits_flow_ingress_node,
  input  [1:0] io_in_flit_0_bits_flow_egress_node,
  input  [1:0] io_in_flit_0_bits_virt_channel_id
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg  in_flight_0; // @[Monitor.scala 16:26]
  reg  in_flight_1; // @[Monitor.scala 16:26]
  reg  in_flight_2; // @[Monitor.scala 16:26]
  reg  in_flight_3; // @[Monitor.scala 16:26]
  wire  _GEN_0 = 2'h0 == io_in_flit_0_bits_virt_channel_id | in_flight_0; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_1 = 2'h1 == io_in_flit_0_bits_virt_channel_id | in_flight_1; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_2 = 2'h2 == io_in_flit_0_bits_virt_channel_id | in_flight_2; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_3 = 2'h3 == io_in_flit_0_bits_virt_channel_id | in_flight_3; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_5 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? in_flight_1 : in_flight_0; // @[Monitor.scala 22:{17,17}]
  wire  _GEN_6 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? in_flight_2 : _GEN_5; // @[Monitor.scala 22:{17,17}]
  wire  _GEN_7 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? in_flight_3 : _GEN_6; // @[Monitor.scala 22:{17,17}]
  wire  _T_2 = ~reset; // @[Monitor.scala 22:16]
  wire  _GEN_8 = io_in_flit_0_bits_head ? _GEN_0 : in_flight_0; // @[Monitor.scala 16:26 20:29]
  wire  _GEN_9 = io_in_flit_0_bits_head ? _GEN_1 : in_flight_1; // @[Monitor.scala 16:26 20:29]
  wire  _GEN_10 = io_in_flit_0_bits_head ? _GEN_2 : in_flight_2; // @[Monitor.scala 16:26 20:29]
  wire  _GEN_11 = io_in_flit_0_bits_head ? _GEN_3 : in_flight_3; // @[Monitor.scala 16:26 20:29]
  wire  _T_4 = io_in_flit_0_valid & io_in_flit_0_bits_head; // @[Monitor.scala 29:22]
  wire  _T_7 = io_in_flit_0_bits_flow_egress_node == 2'h2; // @[Types.scala 54:21]
  wire  _T_8 = io_in_flit_0_bits_flow_ingress_node == 2'h0 & _T_7; // @[Types.scala 53:39]
  wire  _T_27 = io_in_flit_0_bits_flow_ingress_node == 2'h1 & _T_7; // @[Types.scala 53:39]
  wire  _T_33 = io_in_flit_0_bits_flow_egress_node == 2'h3; // @[Types.scala 54:21]
  wire  _T_34 = io_in_flit_0_bits_flow_ingress_node == 2'h1 & _T_33; // @[Types.scala 53:39]
  wire  _T_40 = _T_8 | _T_27 | _T_34; // @[package.scala 73:59]
  wire  _GEN_29 = _T_4 & ~reset; // @[Monitor.scala 22:16]
  always @(posedge clock) begin
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_0 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h0 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_0 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_0 <= _GEN_8;
        end
      end else begin
        in_flight_0 <= _GEN_8;
      end
    end
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_1 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h1 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_1 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_1 <= _GEN_9;
        end
      end else begin
        in_flight_1 <= _GEN_9;
      end
    end
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_2 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h2 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_2 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_2 <= _GEN_10;
        end
      end else begin
        in_flight_2 <= _GEN_10;
      end
    end
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_3 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h3 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_3 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_3 <= _GEN_11;
        end
      end else begin
        in_flight_3 <= _GEN_11;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4 & ~reset & ~(~_GEN_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed: Flit head/tail sequencing is broken\n    at Monitor.scala:22 assert (!in_flight(flit.bits.virt_channel_id), \"Flit head/tail sequencing is broken\")\n"
            ); // @[Monitor.scala 22:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h0 | _T_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h1 | _T_40)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h2 | _T_40)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h3 | _T_40)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  in_flight_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  in_flight_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  in_flight_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  in_flight_3 = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (_T_4 & ~reset) begin
      assert(~_GEN_7); // @[Monitor.scala 22:16]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h0 | _T_8); // @[Monitor.scala 32:17]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h1 | _T_40); // @[Monitor.scala 32:17]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h2 | _T_40); // @[Monitor.scala 32:17]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h3 | _T_40); // @[Monitor.scala 32:17]
    end
  end
endmodule
module NoCMonitor_5(
  input        clock,
  input        reset,
  input        io_in_flit_0_valid,
  input        io_in_flit_0_bits_head,
  input        io_in_flit_0_bits_tail,
  input  [1:0] io_in_flit_0_bits_flow_ingress_node,
  input  [1:0] io_in_flit_0_bits_flow_egress_node,
  input  [1:0] io_in_flit_0_bits_virt_channel_id
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg  in_flight_0; // @[Monitor.scala 16:26]
  reg  in_flight_1; // @[Monitor.scala 16:26]
  reg  in_flight_2; // @[Monitor.scala 16:26]
  reg  in_flight_3; // @[Monitor.scala 16:26]
  wire  _GEN_0 = 2'h0 == io_in_flit_0_bits_virt_channel_id | in_flight_0; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_1 = 2'h1 == io_in_flit_0_bits_virt_channel_id | in_flight_1; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_2 = 2'h2 == io_in_flit_0_bits_virt_channel_id | in_flight_2; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_3 = 2'h3 == io_in_flit_0_bits_virt_channel_id | in_flight_3; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_5 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? in_flight_1 : in_flight_0; // @[Monitor.scala 22:{17,17}]
  wire  _GEN_6 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? in_flight_2 : _GEN_5; // @[Monitor.scala 22:{17,17}]
  wire  _GEN_7 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? in_flight_3 : _GEN_6; // @[Monitor.scala 22:{17,17}]
  wire  _T_2 = ~reset; // @[Monitor.scala 22:16]
  wire  _GEN_8 = io_in_flit_0_bits_head ? _GEN_0 : in_flight_0; // @[Monitor.scala 16:26 20:29]
  wire  _GEN_9 = io_in_flit_0_bits_head ? _GEN_1 : in_flight_1; // @[Monitor.scala 16:26 20:29]
  wire  _GEN_10 = io_in_flit_0_bits_head ? _GEN_2 : in_flight_2; // @[Monitor.scala 16:26 20:29]
  wire  _GEN_11 = io_in_flit_0_bits_head ? _GEN_3 : in_flight_3; // @[Monitor.scala 16:26 20:29]
  wire  _T_4 = io_in_flit_0_valid & io_in_flit_0_bits_head; // @[Monitor.scala 29:22]
  wire  _T_7 = io_in_flit_0_bits_flow_egress_node == 2'h2; // @[Types.scala 54:21]
  wire  _T_8 = io_in_flit_0_bits_flow_ingress_node == 2'h0 & _T_7; // @[Types.scala 53:39]
  wire  _T_26 = io_in_flit_0_bits_flow_egress_node == 2'h1; // @[Types.scala 54:21]
  wire  _T_27 = io_in_flit_0_bits_flow_ingress_node == 2'h3 & _T_26; // @[Types.scala 53:39]
  wire  _T_34 = io_in_flit_0_bits_flow_ingress_node == 2'h3 & _T_7; // @[Types.scala 53:39]
  wire  _T_40 = _T_8 | _T_27 | _T_34; // @[package.scala 73:59]
  wire  _GEN_29 = _T_4 & ~reset; // @[Monitor.scala 22:16]
  always @(posedge clock) begin
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_0 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h0 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_0 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_0 <= _GEN_8;
        end
      end else begin
        in_flight_0 <= _GEN_8;
      end
    end
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_1 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h1 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_1 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_1 <= _GEN_9;
        end
      end else begin
        in_flight_1 <= _GEN_9;
      end
    end
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_2 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h2 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_2 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_2 <= _GEN_10;
        end
      end else begin
        in_flight_2 <= _GEN_10;
      end
    end
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_3 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h3 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_3 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_3 <= _GEN_11;
        end
      end else begin
        in_flight_3 <= _GEN_11;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4 & ~reset & ~(~_GEN_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed: Flit head/tail sequencing is broken\n    at Monitor.scala:22 assert (!in_flight(flit.bits.virt_channel_id), \"Flit head/tail sequencing is broken\")\n"
            ); // @[Monitor.scala 22:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h0 | _T_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h1 | _T_40)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h2 | _T_40)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h3 | _T_40)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  in_flight_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  in_flight_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  in_flight_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  in_flight_3 = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (_T_4 & ~reset) begin
      assert(~_GEN_7); // @[Monitor.scala 22:16]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h0 | _T_8); // @[Monitor.scala 32:17]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h1 | _T_40); // @[Monitor.scala 32:17]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h2 | _T_40); // @[Monitor.scala 32:17]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h3 | _T_40); // @[Monitor.scala 32:17]
    end
  end
endmodule
module InputUnit_4(
  input         clock,
  input         reset,
  output        io_router_req_valid,
  output [1:0]  io_router_req_bits_src_virt_id,
  output [1:0]  io_router_req_bits_flow_ingress_node,
  output [1:0]  io_router_req_bits_flow_egress_node,
  input         io_router_resp_vc_sel_1_0,
  input         io_router_resp_vc_sel_1_1,
  input         io_router_resp_vc_sel_1_2,
  input         io_router_resp_vc_sel_1_3,
  input         io_router_resp_vc_sel_0_0,
  input         io_router_resp_vc_sel_0_1,
  input         io_router_resp_vc_sel_0_2,
  input         io_router_resp_vc_sel_0_3,
  input         io_vcalloc_req_ready,
  output        io_vcalloc_req_valid,
  output        io_vcalloc_req_bits_vc_sel_2_0,
  output        io_vcalloc_req_bits_vc_sel_1_0,
  output        io_vcalloc_req_bits_vc_sel_1_1,
  output        io_vcalloc_req_bits_vc_sel_1_2,
  output        io_vcalloc_req_bits_vc_sel_1_3,
  output        io_vcalloc_req_bits_vc_sel_0_0,
  output        io_vcalloc_req_bits_vc_sel_0_1,
  output        io_vcalloc_req_bits_vc_sel_0_2,
  output        io_vcalloc_req_bits_vc_sel_0_3,
  input         io_vcalloc_resp_vc_sel_2_0,
  input         io_vcalloc_resp_vc_sel_1_0,
  input         io_vcalloc_resp_vc_sel_1_1,
  input         io_vcalloc_resp_vc_sel_1_2,
  input         io_vcalloc_resp_vc_sel_1_3,
  input         io_vcalloc_resp_vc_sel_0_0,
  input         io_vcalloc_resp_vc_sel_0_1,
  input         io_vcalloc_resp_vc_sel_0_2,
  input         io_vcalloc_resp_vc_sel_0_3,
  input         io_out_credit_available_2_0,
  input         io_out_credit_available_1_0,
  input         io_out_credit_available_1_1,
  input         io_out_credit_available_1_2,
  input         io_out_credit_available_1_3,
  input         io_out_credit_available_0_0,
  input         io_out_credit_available_0_1,
  input         io_out_credit_available_0_2,
  input         io_out_credit_available_0_3,
  input         io_salloc_req_0_ready,
  output        io_salloc_req_0_valid,
  output        io_salloc_req_0_bits_vc_sel_2_0,
  output        io_salloc_req_0_bits_vc_sel_1_0,
  output        io_salloc_req_0_bits_vc_sel_1_1,
  output        io_salloc_req_0_bits_vc_sel_1_2,
  output        io_salloc_req_0_bits_vc_sel_1_3,
  output        io_salloc_req_0_bits_vc_sel_0_0,
  output        io_salloc_req_0_bits_vc_sel_0_1,
  output        io_salloc_req_0_bits_vc_sel_0_2,
  output        io_salloc_req_0_bits_vc_sel_0_3,
  output        io_salloc_req_0_bits_tail,
  output        io_out_0_valid,
  output        io_out_0_bits_flit_head,
  output        io_out_0_bits_flit_tail,
  output [63:0] io_out_0_bits_flit_payload,
  output [1:0]  io_out_0_bits_flit_flow_ingress_node,
  output [1:0]  io_out_0_bits_flit_flow_egress_node,
  output [1:0]  io_out_0_bits_out_virt_channel,
  output [1:0]  io_debug_va_stall,
  output [1:0]  io_debug_sa_stall,
  input         io_in_flit_0_valid,
  input         io_in_flit_0_bits_head,
  input         io_in_flit_0_bits_tail,
  input  [63:0] io_in_flit_0_bits_payload,
  input  [1:0]  io_in_flit_0_bits_flow_ingress_node,
  input  [1:0]  io_in_flit_0_bits_flow_egress_node,
  input  [1:0]  io_in_flit_0_bits_virt_channel_id,
  output [3:0]  io_in_credit_return,
  output [3:0]  io_in_vc_free
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
`endif // RANDOMIZE_REG_INIT
  wire  input_buffer_clock; // @[InputUnit.scala 180:28]
  wire  input_buffer_reset; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_enq_0_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_enq_0_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_enq_0_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_enq_0_bits_payload; // @[InputUnit.scala 180:28]
  wire [1:0] input_buffer_io_enq_0_bits_virt_channel_id; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_0_ready; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_0_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_0_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_0_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_deq_0_bits_payload; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_ready; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_deq_1_bits_payload; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_ready; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_deq_2_bits_payload; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_3_ready; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_3_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_3_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_3_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_deq_3_bits_payload; // @[InputUnit.scala 180:28]
  wire  route_arbiter_io_in_0_valid; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_0_bits_flow_ingress_node; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_0_bits_flow_egress_node; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_1_ready; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_1_valid; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_1_bits_flow_ingress_node; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_1_bits_flow_egress_node; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_2_ready; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_2_valid; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_2_bits_flow_ingress_node; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_2_bits_flow_egress_node; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_3_ready; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_3_valid; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_3_bits_flow_ingress_node; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_3_bits_flow_egress_node; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_out_valid; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_out_bits_src_virt_id; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_out_bits_flow_ingress_node; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_out_bits_flow_egress_node; // @[InputUnit.scala 186:29]
  wire  salloc_arb_clock; // @[InputUnit.scala 279:26]
  wire  salloc_arb_reset; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_bits_vc_sel_2_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_bits_vc_sel_1_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_bits_tail; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_vc_sel_2_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_vc_sel_1_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_vc_sel_1_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_vc_sel_0_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_tail; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_2_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_1_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_1_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_1_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_0_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_0_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_tail; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_2_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_1_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_1_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_1_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_1_3; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_0_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_0_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_0_3; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_tail; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_2_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_1_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_1_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_1_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_1_3; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_0_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_0_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_0_3; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_tail; // @[InputUnit.scala 279:26]
  wire [3:0] salloc_arb_io_chosen_oh_0; // @[InputUnit.scala 279:26]
  reg [2:0] states_0_g; // @[InputUnit.scala 191:19]
  reg  states_0_vc_sel_2_0; // @[InputUnit.scala 191:19]
  reg  states_0_vc_sel_1_0; // @[InputUnit.scala 191:19]
  reg  states_0_vc_sel_0_0; // @[InputUnit.scala 191:19]
  reg [1:0] states_0_flow_ingress_node; // @[InputUnit.scala 191:19]
  reg [1:0] states_0_flow_egress_node; // @[InputUnit.scala 191:19]
  reg [2:0] states_1_g; // @[InputUnit.scala 191:19]
  reg  states_1_vc_sel_2_0; // @[InputUnit.scala 191:19]
  reg  states_1_vc_sel_1_0; // @[InputUnit.scala 191:19]
  reg  states_1_vc_sel_1_1; // @[InputUnit.scala 191:19]
  reg  states_1_vc_sel_0_1; // @[InputUnit.scala 191:19]
  reg [1:0] states_1_flow_ingress_node; // @[InputUnit.scala 191:19]
  reg [1:0] states_1_flow_egress_node; // @[InputUnit.scala 191:19]
  reg [2:0] states_2_g; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_2_0; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_1_0; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_1_1; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_1_2; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_0_1; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_0_2; // @[InputUnit.scala 191:19]
  reg [1:0] states_2_flow_ingress_node; // @[InputUnit.scala 191:19]
  reg [1:0] states_2_flow_egress_node; // @[InputUnit.scala 191:19]
  reg [2:0] states_3_g; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_2_0; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_1_0; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_1_1; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_1_2; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_1_3; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_0_1; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_0_2; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_0_3; // @[InputUnit.scala 191:19]
  reg [1:0] states_3_flow_ingress_node; // @[InputUnit.scala 191:19]
  reg [1:0] states_3_flow_egress_node; // @[InputUnit.scala 191:19]
  wire  _T = io_in_flit_0_valid & io_in_flit_0_bits_head; // @[InputUnit.scala 194:32]
  wire  _T_3 = ~reset; // @[InputUnit.scala 196:13]
  wire [2:0] _GEN_1 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? states_1_g : states_0_g; // @[InputUnit.scala 197:{27,27}]
  wire [2:0] _GEN_2 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? states_2_g : _GEN_1; // @[InputUnit.scala 197:{27,27}]
  wire [2:0] _GEN_3 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? states_3_g : _GEN_2; // @[InputUnit.scala 197:{27,27}]
  wire  at_dest = io_in_flit_0_bits_flow_egress_node == 2'h2; // @[InputUnit.scala 198:57]
  wire [2:0] _states_g_T = at_dest ? 3'h2 : 3'h1; // @[InputUnit.scala 199:26]
  wire [2:0] _GEN_4 = 2'h0 == io_in_flit_0_bits_virt_channel_id ? _states_g_T : states_0_g; // @[InputUnit.scala 191:19 199:{20,20}]
  wire [2:0] _GEN_5 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? _states_g_T : states_1_g; // @[InputUnit.scala 191:19 199:{20,20}]
  wire [2:0] _GEN_6 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? _states_g_T : states_2_g; // @[InputUnit.scala 191:19 199:{20,20}]
  wire [2:0] _GEN_7 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? _states_g_T : states_3_g; // @[InputUnit.scala 191:19 199:{20,20}]
  wire  _GEN_8 = 2'h0 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_0_vc_sel_0_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_13 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_1_vc_sel_0_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_14 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_0_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_15 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_0_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_18 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_0_2; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_19 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_0_2; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_23 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_0_3; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_24 = 2'h0 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_0_vc_sel_1_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_25 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_1_vc_sel_1_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_26 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_1_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_27 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_1_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_29 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_1_vc_sel_1_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_30 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_1_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_31 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_1_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_34 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_1_2; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_35 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_1_2; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_39 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_1_3; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_40 = 2'h0 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_0_vc_sel_2_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_41 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_1_vc_sel_2_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_42 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_2_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_43 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_2_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_44 = 2'h0 == io_in_flit_0_bits_virt_channel_id | _GEN_40; // @[InputUnit.scala 203:{44,44}]
  wire  _GEN_45 = 2'h1 == io_in_flit_0_bits_virt_channel_id | _GEN_41; // @[InputUnit.scala 203:{44,44}]
  wire  _GEN_46 = 2'h2 == io_in_flit_0_bits_virt_channel_id | _GEN_42; // @[InputUnit.scala 203:{44,44}]
  wire  _GEN_47 = 2'h3 == io_in_flit_0_bits_virt_channel_id | _GEN_43; // @[InputUnit.scala 203:{44,44}]
  wire [2:0] _GEN_72 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_4 : states_0_g; // @[InputUnit.scala 191:19 194:60]
  wire [2:0] _GEN_73 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_5 : states_1_g; // @[InputUnit.scala 191:19 194:60]
  wire [2:0] _GEN_74 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_6 : states_2_g; // @[InputUnit.scala 191:19 194:60]
  wire [2:0] _GEN_75 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_7 : states_3_g; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_76 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_8 : states_0_vc_sel_0_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_81 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_13 : states_1_vc_sel_0_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_82 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_14 : states_2_vc_sel_0_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_83 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_15 : states_3_vc_sel_0_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_86 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_18 : states_2_vc_sel_0_2; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_87 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_19 : states_3_vc_sel_0_2; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_91 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_23 : states_3_vc_sel_0_3; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_92 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_24 : states_0_vc_sel_1_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_93 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_25 : states_1_vc_sel_1_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_94 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_26 : states_2_vc_sel_1_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_95 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_27 : states_3_vc_sel_1_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_97 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_29 : states_1_vc_sel_1_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_98 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_30 : states_2_vc_sel_1_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_99 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_31 : states_3_vc_sel_1_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_102 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_34 : states_2_vc_sel_1_2; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_103 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_35 : states_3_vc_sel_1_2; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_107 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_39 : states_3_vc_sel_1_3; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_108 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_44 : states_0_vc_sel_2_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_109 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_45 : states_1_vc_sel_2_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_110 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_46 : states_2_vc_sel_2_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_111 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_47 : states_3_vc_sel_2_0; // @[InputUnit.scala 191:19 194:60]
  wire  _T_10 = route_arbiter_io_in_0_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_132 = _T_10 ? 3'h2 : _GEN_72; // @[InputUnit.scala 215:{23,29}]
  wire  _T_11 = route_arbiter_io_in_1_ready & route_arbiter_io_in_1_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_133 = _T_11 ? 3'h2 : _GEN_73; // @[InputUnit.scala 215:{23,29}]
  wire  _T_12 = route_arbiter_io_in_2_ready & route_arbiter_io_in_2_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_134 = _T_12 ? 3'h2 : _GEN_74; // @[InputUnit.scala 215:{23,29}]
  wire  _T_13 = route_arbiter_io_in_3_ready & route_arbiter_io_in_3_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_135 = _T_13 ? 3'h2 : _GEN_75; // @[InputUnit.scala 215:{23,29}]
  wire [2:0] _GEN_137 = 2'h1 == io_router_req_bits_src_virt_id ? states_1_g : states_0_g; // @[InputUnit.scala 224:{25,25}]
  wire [2:0] _GEN_138 = 2'h2 == io_router_req_bits_src_virt_id ? states_2_g : _GEN_137; // @[InputUnit.scala 224:{25,25}]
  wire [2:0] _GEN_139 = 2'h3 == io_router_req_bits_src_virt_id ? states_3_g : _GEN_138; // @[InputUnit.scala 224:{25,25}]
  wire [2:0] _GEN_140 = 2'h0 == io_router_req_bits_src_virt_id ? 3'h2 : _GEN_132; // @[InputUnit.scala 225:{18,18}]
  wire [2:0] _GEN_141 = 2'h1 == io_router_req_bits_src_virt_id ? 3'h2 : _GEN_133; // @[InputUnit.scala 225:{18,18}]
  wire [2:0] _GEN_142 = 2'h2 == io_router_req_bits_src_virt_id ? 3'h2 : _GEN_134; // @[InputUnit.scala 225:{18,18}]
  wire [2:0] _GEN_143 = 2'h3 == io_router_req_bits_src_virt_id ? 3'h2 : _GEN_135; // @[InputUnit.scala 225:{18,18}]
  wire  _GEN_144 = 2'h0 == io_router_req_bits_src_virt_id ? 1'h0 : _GEN_108; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_145 = 2'h0 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_0 : _GEN_92; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_149 = 2'h0 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_0 : _GEN_76; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_153 = 2'h1 == io_router_req_bits_src_virt_id ? 1'h0 : _GEN_109; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_154 = 2'h1 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_0 : _GEN_93; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_155 = 2'h1 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_1 : _GEN_97; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_159 = 2'h1 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_1 : _GEN_81; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_162 = 2'h2 == io_router_req_bits_src_virt_id ? 1'h0 : _GEN_110; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_163 = 2'h2 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_0 : _GEN_94; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_164 = 2'h2 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_1 : _GEN_98; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_165 = 2'h2 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_2 : _GEN_102; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_168 = 2'h2 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_1 : _GEN_82; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_169 = 2'h2 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_2 : _GEN_86; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_171 = 2'h3 == io_router_req_bits_src_virt_id ? 1'h0 : _GEN_111; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_172 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_0 : _GEN_95; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_173 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_1 : _GEN_99; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_174 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_2 : _GEN_103; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_175 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_3 : _GEN_107; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_177 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_1 : _GEN_83; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_178 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_2 : _GEN_87; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_179 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_3 : _GEN_91; // @[InputUnit.scala 227:25 228:26]
  wire [2:0] _GEN_180 = io_router_req_valid ? _GEN_140 : _GEN_132; // @[InputUnit.scala 222:31]
  wire [2:0] _GEN_181 = io_router_req_valid ? _GEN_141 : _GEN_133; // @[InputUnit.scala 222:31]
  wire [2:0] _GEN_182 = io_router_req_valid ? _GEN_142 : _GEN_134; // @[InputUnit.scala 222:31]
  wire [2:0] _GEN_183 = io_router_req_valid ? _GEN_143 : _GEN_135; // @[InputUnit.scala 222:31]
  wire  _GEN_184 = io_router_req_valid ? _GEN_144 : _GEN_108; // @[InputUnit.scala 222:31]
  wire  _GEN_185 = io_router_req_valid ? _GEN_145 : _GEN_92; // @[InputUnit.scala 222:31]
  wire  _GEN_189 = io_router_req_valid ? _GEN_149 : _GEN_76; // @[InputUnit.scala 222:31]
  wire  _GEN_193 = io_router_req_valid ? _GEN_153 : _GEN_109; // @[InputUnit.scala 222:31]
  wire  _GEN_194 = io_router_req_valid ? _GEN_154 : _GEN_93; // @[InputUnit.scala 222:31]
  wire  _GEN_195 = io_router_req_valid ? _GEN_155 : _GEN_97; // @[InputUnit.scala 222:31]
  wire  _GEN_199 = io_router_req_valid ? _GEN_159 : _GEN_81; // @[InputUnit.scala 222:31]
  wire  _GEN_202 = io_router_req_valid ? _GEN_162 : _GEN_110; // @[InputUnit.scala 222:31]
  wire  _GEN_203 = io_router_req_valid ? _GEN_163 : _GEN_94; // @[InputUnit.scala 222:31]
  wire  _GEN_204 = io_router_req_valid ? _GEN_164 : _GEN_98; // @[InputUnit.scala 222:31]
  wire  _GEN_205 = io_router_req_valid ? _GEN_165 : _GEN_102; // @[InputUnit.scala 222:31]
  wire  _GEN_208 = io_router_req_valid ? _GEN_168 : _GEN_82; // @[InputUnit.scala 222:31]
  wire  _GEN_209 = io_router_req_valid ? _GEN_169 : _GEN_86; // @[InputUnit.scala 222:31]
  wire  _GEN_211 = io_router_req_valid ? _GEN_171 : _GEN_111; // @[InputUnit.scala 222:31]
  wire  _GEN_212 = io_router_req_valid ? _GEN_172 : _GEN_95; // @[InputUnit.scala 222:31]
  wire  _GEN_213 = io_router_req_valid ? _GEN_173 : _GEN_99; // @[InputUnit.scala 222:31]
  wire  _GEN_214 = io_router_req_valid ? _GEN_174 : _GEN_103; // @[InputUnit.scala 222:31]
  wire  _GEN_215 = io_router_req_valid ? _GEN_175 : _GEN_107; // @[InputUnit.scala 222:31]
  wire  _GEN_217 = io_router_req_valid ? _GEN_177 : _GEN_83; // @[InputUnit.scala 222:31]
  wire  _GEN_218 = io_router_req_valid ? _GEN_178 : _GEN_87; // @[InputUnit.scala 222:31]
  wire  _GEN_219 = io_router_req_valid ? _GEN_179 : _GEN_91; // @[InputUnit.scala 222:31]
  reg [3:0] mask; // @[InputUnit.scala 233:21]
  wire  vcalloc_vals_1 = states_1_g == 3'h2; // @[InputUnit.scala 249:32]
  wire  vcalloc_vals_0 = states_0_g == 3'h2; // @[InputUnit.scala 249:32]
  wire  vcalloc_vals_3 = states_3_g == 3'h2; // @[InputUnit.scala 249:32]
  wire  vcalloc_vals_2 = states_2_g == 3'h2; // @[InputUnit.scala 249:32]
  wire [3:0] _vcalloc_filter_T = {vcalloc_vals_3,vcalloc_vals_2,vcalloc_vals_1,vcalloc_vals_0}; // @[InputUnit.scala 236:59]
  wire [3:0] _vcalloc_filter_T_2 = ~mask; // @[InputUnit.scala 236:89]
  wire [3:0] _vcalloc_filter_T_3 = _vcalloc_filter_T & _vcalloc_filter_T_2; // @[InputUnit.scala 236:87]
  wire [7:0] _vcalloc_filter_T_4 = {vcalloc_vals_3,vcalloc_vals_2,vcalloc_vals_1,vcalloc_vals_0,_vcalloc_filter_T_3}; // @[Cat.scala 33:92]
  wire [7:0] _vcalloc_filter_T_13 = _vcalloc_filter_T_4[7] ? 8'h80 : 8'h0; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_14 = _vcalloc_filter_T_4[6] ? 8'h40 : _vcalloc_filter_T_13; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_15 = _vcalloc_filter_T_4[5] ? 8'h20 : _vcalloc_filter_T_14; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_16 = _vcalloc_filter_T_4[4] ? 8'h10 : _vcalloc_filter_T_15; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_17 = _vcalloc_filter_T_4[3] ? 8'h8 : _vcalloc_filter_T_16; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_18 = _vcalloc_filter_T_4[2] ? 8'h4 : _vcalloc_filter_T_17; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_19 = _vcalloc_filter_T_4[1] ? 8'h2 : _vcalloc_filter_T_18; // @[Mux.scala 47:70]
  wire [7:0] vcalloc_filter = _vcalloc_filter_T_4[0] ? 8'h1 : _vcalloc_filter_T_19; // @[Mux.scala 47:70]
  wire [3:0] vcalloc_sel = vcalloc_filter[3:0] | vcalloc_filter[7:4]; // @[InputUnit.scala 237:58]
  wire [3:0] _mask_T = 4'h1 << io_router_req_bits_src_virt_id; // @[InputUnit.scala 240:18]
  wire [3:0] _mask_T_2 = _mask_T - 4'h1; // @[InputUnit.scala 240:53]
  wire  _T_26 = vcalloc_vals_0 | vcalloc_vals_1 | vcalloc_vals_2 | vcalloc_vals_3; // @[package.scala 73:59]
  wire [1:0] _mask_T_12 = vcalloc_sel[1] ? 2'h3 : 2'h0; // @[Mux.scala 27:73]
  wire [2:0] _mask_T_13 = vcalloc_sel[2] ? 3'h7 : 3'h0; // @[Mux.scala 27:73]
  wire [3:0] _mask_T_14 = vcalloc_sel[3] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [1:0] _GEN_60 = {{1'd0}, vcalloc_sel[0]}; // @[Mux.scala 27:73]
  wire [1:0] _mask_T_15 = _GEN_60 | _mask_T_12; // @[Mux.scala 27:73]
  wire [2:0] _GEN_61 = {{1'd0}, _mask_T_15}; // @[Mux.scala 27:73]
  wire [2:0] _mask_T_16 = _GEN_61 | _mask_T_13; // @[Mux.scala 27:73]
  wire [3:0] _GEN_62 = {{1'd0}, _mask_T_16}; // @[Mux.scala 27:73]
  wire [3:0] _mask_T_17 = _GEN_62 | _mask_T_14; // @[Mux.scala 27:73]
  wire [2:0] _GEN_222 = vcalloc_vals_0 & vcalloc_sel[0] & io_vcalloc_req_ready ? 3'h3 : _GEN_180; // @[InputUnit.scala 253:{76,82}]
  wire [2:0] _GEN_223 = vcalloc_vals_1 & vcalloc_sel[1] & io_vcalloc_req_ready ? 3'h3 : _GEN_181; // @[InputUnit.scala 253:{76,82}]
  wire [2:0] _GEN_224 = vcalloc_vals_2 & vcalloc_sel[2] & io_vcalloc_req_ready ? 3'h3 : _GEN_182; // @[InputUnit.scala 253:{76,82}]
  wire [2:0] _GEN_225 = vcalloc_vals_3 & vcalloc_sel[3] & io_vcalloc_req_ready ? 3'h3 : _GEN_183; // @[InputUnit.scala 253:{76,82}]
  wire [1:0] _io_debug_va_stall_T = vcalloc_vals_0 + vcalloc_vals_1; // @[Bitwise.scala 51:90]
  wire [1:0] _io_debug_va_stall_T_2 = vcalloc_vals_2 + vcalloc_vals_3; // @[Bitwise.scala 51:90]
  wire [2:0] _io_debug_va_stall_T_4 = _io_debug_va_stall_T + _io_debug_va_stall_T_2; // @[Bitwise.scala 51:90]
  wire [2:0] _GEN_63 = {{2'd0}, io_vcalloc_req_ready}; // @[InputUnit.scala 266:47]
  wire [2:0] _io_debug_va_stall_T_7 = _io_debug_va_stall_T_4 - _GEN_63; // @[InputUnit.scala 266:47]
  wire  _T_39 = io_vcalloc_req_ready & io_vcalloc_req_valid; // @[Decoupled.scala 51:35]
  wire [8:0] _credit_available_T = {states_0_vc_sel_2_0,1'h0,1'h0,1'h0,states_0_vc_sel_1_0,2'h0,1'h0,states_0_vc_sel_0_0
    }; // @[InputUnit.scala 287:40]
  wire [8:0] _credit_available_T_1 = {io_out_credit_available_2_0,io_out_credit_available_1_3,
    io_out_credit_available_1_2,io_out_credit_available_1_1,io_out_credit_available_1_0,io_out_credit_available_0_3,
    io_out_credit_available_0_2,io_out_credit_available_0_1,io_out_credit_available_0_0}; // @[InputUnit.scala 287:73]
  wire [8:0] _credit_available_T_2 = _credit_available_T & _credit_available_T_1; // @[InputUnit.scala 287:47]
  wire  credit_available = _credit_available_T_2 != 9'h0; // @[InputUnit.scala 287:81]
  wire  _T_60 = salloc_arb_io_in_0_ready & salloc_arb_io_in_0_valid; // @[Decoupled.scala 51:35]
  wire [8:0] _credit_available_T_3 = {states_1_vc_sel_2_0,1'h0,1'h0,states_1_vc_sel_1_1,states_1_vc_sel_1_0,2'h0,
    states_1_vc_sel_0_1,1'h0}; // @[InputUnit.scala 287:40]
  wire [8:0] _credit_available_T_5 = _credit_available_T_3 & _credit_available_T_1; // @[InputUnit.scala 287:47]
  wire  credit_available_1 = _credit_available_T_5 != 9'h0; // @[InputUnit.scala 287:81]
  wire  _T_62 = salloc_arb_io_in_1_ready & salloc_arb_io_in_1_valid; // @[Decoupled.scala 51:35]
  wire [8:0] _credit_available_T_6 = {states_2_vc_sel_2_0,1'h0,states_2_vc_sel_1_2,states_2_vc_sel_1_1,
    states_2_vc_sel_1_0,1'h0,states_2_vc_sel_0_2,states_2_vc_sel_0_1,1'h0}; // @[InputUnit.scala 287:40]
  wire [8:0] _credit_available_T_8 = _credit_available_T_6 & _credit_available_T_1; // @[InputUnit.scala 287:47]
  wire  credit_available_2 = _credit_available_T_8 != 9'h0; // @[InputUnit.scala 287:81]
  wire  _T_64 = salloc_arb_io_in_2_ready & salloc_arb_io_in_2_valid; // @[Decoupled.scala 51:35]
  wire [8:0] _credit_available_T_9 = {states_3_vc_sel_2_0,states_3_vc_sel_1_3,states_3_vc_sel_1_2,states_3_vc_sel_1_1,
    states_3_vc_sel_1_0,states_3_vc_sel_0_3,states_3_vc_sel_0_2,states_3_vc_sel_0_1,1'h0}; // @[InputUnit.scala 287:40]
  wire [8:0] _credit_available_T_11 = _credit_available_T_9 & _credit_available_T_1; // @[InputUnit.scala 287:47]
  wire  credit_available_3 = _credit_available_T_11 != 9'h0; // @[InputUnit.scala 287:81]
  wire  _T_66 = salloc_arb_io_in_3_ready & salloc_arb_io_in_3_valid; // @[Decoupled.scala 51:35]
  wire  _io_debug_sa_stall_T_1 = salloc_arb_io_in_0_valid & ~salloc_arb_io_in_0_ready; // @[InputUnit.scala 301:67]
  wire  _io_debug_sa_stall_T_3 = salloc_arb_io_in_1_valid & ~salloc_arb_io_in_1_ready; // @[InputUnit.scala 301:67]
  wire  _io_debug_sa_stall_T_5 = salloc_arb_io_in_2_valid & ~salloc_arb_io_in_2_ready; // @[InputUnit.scala 301:67]
  wire  _io_debug_sa_stall_T_7 = salloc_arb_io_in_3_valid & ~salloc_arb_io_in_3_ready; // @[InputUnit.scala 301:67]
  wire [1:0] _io_debug_sa_stall_T_8 = _io_debug_sa_stall_T_1 + _io_debug_sa_stall_T_3; // @[Bitwise.scala 51:90]
  wire [1:0] _io_debug_sa_stall_T_10 = _io_debug_sa_stall_T_5 + _io_debug_sa_stall_T_7; // @[Bitwise.scala 51:90]
  wire [2:0] _io_debug_sa_stall_T_12 = _io_debug_sa_stall_T_8 + _io_debug_sa_stall_T_10; // @[Bitwise.scala 51:90]
  reg  salloc_outs_0_valid; // @[InputUnit.scala 318:8]
  reg [1:0] salloc_outs_0_out_vid; // @[InputUnit.scala 318:8]
  reg  salloc_outs_0_flit_head; // @[InputUnit.scala 318:8]
  reg  salloc_outs_0_flit_tail; // @[InputUnit.scala 318:8]
  reg [63:0] salloc_outs_0_flit_payload; // @[InputUnit.scala 318:8]
  reg [1:0] salloc_outs_0_flit_flow_ingress_node; // @[InputUnit.scala 318:8]
  reg [1:0] salloc_outs_0_flit_flow_egress_node; // @[InputUnit.scala 318:8]
  wire  _io_in_credit_return_T = salloc_arb_io_out_0_ready & salloc_arb_io_out_0_valid; // @[Decoupled.scala 51:35]
  wire  _io_in_vc_free_T_11 = salloc_arb_io_chosen_oh_0[0] & input_buffer_io_deq_0_bits_tail | salloc_arb_io_chosen_oh_0
    [1] & input_buffer_io_deq_1_bits_tail | salloc_arb_io_chosen_oh_0[2] & input_buffer_io_deq_2_bits_tail |
    salloc_arb_io_chosen_oh_0[3] & input_buffer_io_deq_3_bits_tail; // @[Mux.scala 27:73]
  wire  vc_sel_0_0 = salloc_arb_io_chosen_oh_0[0] & states_0_vc_sel_0_0; // @[Mux.scala 27:73]
  wire  vc_sel_0_1 = salloc_arb_io_chosen_oh_0[1] & states_1_vc_sel_0_1 | salloc_arb_io_chosen_oh_0[2] &
    states_2_vc_sel_0_1 | salloc_arb_io_chosen_oh_0[3] & states_3_vc_sel_0_1; // @[Mux.scala 27:73]
  wire  vc_sel_0_2 = salloc_arb_io_chosen_oh_0[2] & states_2_vc_sel_0_2 | salloc_arb_io_chosen_oh_0[3] &
    states_3_vc_sel_0_2; // @[Mux.scala 27:73]
  wire  vc_sel_0_3 = salloc_arb_io_chosen_oh_0[3] & states_3_vc_sel_0_3; // @[Mux.scala 27:73]
  wire  vc_sel_1_0 = salloc_arb_io_chosen_oh_0[0] & states_0_vc_sel_1_0 | salloc_arb_io_chosen_oh_0[1] &
    states_1_vc_sel_1_0 | salloc_arb_io_chosen_oh_0[2] & states_2_vc_sel_1_0 | salloc_arb_io_chosen_oh_0[3] &
    states_3_vc_sel_1_0; // @[Mux.scala 27:73]
  wire  vc_sel_1_1 = salloc_arb_io_chosen_oh_0[1] & states_1_vc_sel_1_1 | salloc_arb_io_chosen_oh_0[2] &
    states_2_vc_sel_1_1 | salloc_arb_io_chosen_oh_0[3] & states_3_vc_sel_1_1; // @[Mux.scala 27:73]
  wire  vc_sel_1_2 = salloc_arb_io_chosen_oh_0[2] & states_2_vc_sel_1_2 | salloc_arb_io_chosen_oh_0[3] &
    states_3_vc_sel_1_2; // @[Mux.scala 27:73]
  wire  vc_sel_1_3 = salloc_arb_io_chosen_oh_0[3] & states_3_vc_sel_1_3; // @[Mux.scala 27:73]
  wire  channel_oh_0 = vc_sel_0_0 | vc_sel_0_1 | vc_sel_0_2 | vc_sel_0_3; // @[InputUnit.scala 334:43]
  wire  channel_oh_1 = vc_sel_1_0 | vc_sel_1_1 | vc_sel_1_2 | vc_sel_1_3; // @[InputUnit.scala 334:43]
  wire [3:0] _virt_channel_T = {vc_sel_0_3,vc_sel_0_2,vc_sel_0_1,vc_sel_0_0}; // @[OneHot.scala 22:45]
  wire [1:0] virt_channel_hi_1 = _virt_channel_T[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] virt_channel_lo_1 = _virt_channel_T[1:0]; // @[OneHot.scala 31:18]
  wire  _virt_channel_T_1 = |virt_channel_hi_1; // @[OneHot.scala 32:14]
  wire [1:0] _virt_channel_T_2 = virt_channel_hi_1 | virt_channel_lo_1; // @[OneHot.scala 32:28]
  wire [1:0] _virt_channel_T_4 = {_virt_channel_T_1,_virt_channel_T_2[1]}; // @[Cat.scala 33:92]
  wire [3:0] _virt_channel_T_5 = {vc_sel_1_3,vc_sel_1_2,vc_sel_1_1,vc_sel_1_0}; // @[OneHot.scala 22:45]
  wire [1:0] virt_channel_hi_3 = _virt_channel_T_5[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] virt_channel_lo_3 = _virt_channel_T_5[1:0]; // @[OneHot.scala 31:18]
  wire  _virt_channel_T_6 = |virt_channel_hi_3; // @[OneHot.scala 32:14]
  wire [1:0] _virt_channel_T_7 = virt_channel_hi_3 | virt_channel_lo_3; // @[OneHot.scala 32:28]
  wire [1:0] _virt_channel_T_9 = {_virt_channel_T_6,_virt_channel_T_7[1]}; // @[Cat.scala 33:92]
  wire [1:0] _virt_channel_T_10 = channel_oh_0 ? _virt_channel_T_4 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _virt_channel_T_11 = channel_oh_1 ? _virt_channel_T_9 : 2'h0; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_4 = salloc_arb_io_chosen_oh_0[0] ? input_buffer_io_deq_0_bits_payload : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_5 = salloc_arb_io_chosen_oh_0[1] ? input_buffer_io_deq_1_bits_payload : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_6 = salloc_arb_io_chosen_oh_0[2] ? input_buffer_io_deq_2_bits_payload : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_7 = salloc_arb_io_chosen_oh_0[3] ? input_buffer_io_deq_3_bits_payload : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_8 = _salloc_outs_0_flit_payload_T_4 | _salloc_outs_0_flit_payload_T_5; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_9 = _salloc_outs_0_flit_payload_T_8 | _salloc_outs_0_flit_payload_T_6; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_11 = salloc_arb_io_chosen_oh_0[0] ? states_0_flow_egress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_12 = salloc_arb_io_chosen_oh_0[1] ? states_1_flow_egress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_13 = salloc_arb_io_chosen_oh_0[2] ? states_2_flow_egress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_14 = salloc_arb_io_chosen_oh_0[3] ? states_3_flow_egress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_15 = _salloc_outs_0_flit_flow_T_11 | _salloc_outs_0_flit_flow_T_12; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_16 = _salloc_outs_0_flit_flow_T_15 | _salloc_outs_0_flit_flow_T_13; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_25 = salloc_arb_io_chosen_oh_0[0] ? states_0_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_26 = salloc_arb_io_chosen_oh_0[1] ? states_1_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_27 = salloc_arb_io_chosen_oh_0[2] ? states_2_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_28 = salloc_arb_io_chosen_oh_0[3] ? states_3_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_29 = _salloc_outs_0_flit_flow_T_25 | _salloc_outs_0_flit_flow_T_26; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_30 = _salloc_outs_0_flit_flow_T_29 | _salloc_outs_0_flit_flow_T_27; // @[Mux.scala 27:73]
  InputBuffer input_buffer ( // @[InputUnit.scala 180:28]
    .clock(input_buffer_clock),
    .reset(input_buffer_reset),
    .io_enq_0_valid(input_buffer_io_enq_0_valid),
    .io_enq_0_bits_head(input_buffer_io_enq_0_bits_head),
    .io_enq_0_bits_tail(input_buffer_io_enq_0_bits_tail),
    .io_enq_0_bits_payload(input_buffer_io_enq_0_bits_payload),
    .io_enq_0_bits_virt_channel_id(input_buffer_io_enq_0_bits_virt_channel_id),
    .io_deq_0_ready(input_buffer_io_deq_0_ready),
    .io_deq_0_valid(input_buffer_io_deq_0_valid),
    .io_deq_0_bits_head(input_buffer_io_deq_0_bits_head),
    .io_deq_0_bits_tail(input_buffer_io_deq_0_bits_tail),
    .io_deq_0_bits_payload(input_buffer_io_deq_0_bits_payload),
    .io_deq_1_ready(input_buffer_io_deq_1_ready),
    .io_deq_1_valid(input_buffer_io_deq_1_valid),
    .io_deq_1_bits_head(input_buffer_io_deq_1_bits_head),
    .io_deq_1_bits_tail(input_buffer_io_deq_1_bits_tail),
    .io_deq_1_bits_payload(input_buffer_io_deq_1_bits_payload),
    .io_deq_2_ready(input_buffer_io_deq_2_ready),
    .io_deq_2_valid(input_buffer_io_deq_2_valid),
    .io_deq_2_bits_head(input_buffer_io_deq_2_bits_head),
    .io_deq_2_bits_tail(input_buffer_io_deq_2_bits_tail),
    .io_deq_2_bits_payload(input_buffer_io_deq_2_bits_payload),
    .io_deq_3_ready(input_buffer_io_deq_3_ready),
    .io_deq_3_valid(input_buffer_io_deq_3_valid),
    .io_deq_3_bits_head(input_buffer_io_deq_3_bits_head),
    .io_deq_3_bits_tail(input_buffer_io_deq_3_bits_tail),
    .io_deq_3_bits_payload(input_buffer_io_deq_3_bits_payload)
  );
  Arbiter route_arbiter ( // @[InputUnit.scala 186:29]
    .io_in_0_valid(route_arbiter_io_in_0_valid),
    .io_in_0_bits_flow_ingress_node(route_arbiter_io_in_0_bits_flow_ingress_node),
    .io_in_0_bits_flow_egress_node(route_arbiter_io_in_0_bits_flow_egress_node),
    .io_in_1_ready(route_arbiter_io_in_1_ready),
    .io_in_1_valid(route_arbiter_io_in_1_valid),
    .io_in_1_bits_flow_ingress_node(route_arbiter_io_in_1_bits_flow_ingress_node),
    .io_in_1_bits_flow_egress_node(route_arbiter_io_in_1_bits_flow_egress_node),
    .io_in_2_ready(route_arbiter_io_in_2_ready),
    .io_in_2_valid(route_arbiter_io_in_2_valid),
    .io_in_2_bits_flow_ingress_node(route_arbiter_io_in_2_bits_flow_ingress_node),
    .io_in_2_bits_flow_egress_node(route_arbiter_io_in_2_bits_flow_egress_node),
    .io_in_3_ready(route_arbiter_io_in_3_ready),
    .io_in_3_valid(route_arbiter_io_in_3_valid),
    .io_in_3_bits_flow_ingress_node(route_arbiter_io_in_3_bits_flow_ingress_node),
    .io_in_3_bits_flow_egress_node(route_arbiter_io_in_3_bits_flow_egress_node),
    .io_out_valid(route_arbiter_io_out_valid),
    .io_out_bits_src_virt_id(route_arbiter_io_out_bits_src_virt_id),
    .io_out_bits_flow_ingress_node(route_arbiter_io_out_bits_flow_ingress_node),
    .io_out_bits_flow_egress_node(route_arbiter_io_out_bits_flow_egress_node)
  );
  SwitchArbiter salloc_arb ( // @[InputUnit.scala 279:26]
    .clock(salloc_arb_clock),
    .reset(salloc_arb_reset),
    .io_in_0_ready(salloc_arb_io_in_0_ready),
    .io_in_0_valid(salloc_arb_io_in_0_valid),
    .io_in_0_bits_vc_sel_2_0(salloc_arb_io_in_0_bits_vc_sel_2_0),
    .io_in_0_bits_vc_sel_1_0(salloc_arb_io_in_0_bits_vc_sel_1_0),
    .io_in_0_bits_vc_sel_0_0(salloc_arb_io_in_0_bits_vc_sel_0_0),
    .io_in_0_bits_tail(salloc_arb_io_in_0_bits_tail),
    .io_in_1_ready(salloc_arb_io_in_1_ready),
    .io_in_1_valid(salloc_arb_io_in_1_valid),
    .io_in_1_bits_vc_sel_2_0(salloc_arb_io_in_1_bits_vc_sel_2_0),
    .io_in_1_bits_vc_sel_1_0(salloc_arb_io_in_1_bits_vc_sel_1_0),
    .io_in_1_bits_vc_sel_1_1(salloc_arb_io_in_1_bits_vc_sel_1_1),
    .io_in_1_bits_vc_sel_0_0(salloc_arb_io_in_1_bits_vc_sel_0_0),
    .io_in_1_bits_vc_sel_0_1(salloc_arb_io_in_1_bits_vc_sel_0_1),
    .io_in_1_bits_tail(salloc_arb_io_in_1_bits_tail),
    .io_in_2_ready(salloc_arb_io_in_2_ready),
    .io_in_2_valid(salloc_arb_io_in_2_valid),
    .io_in_2_bits_vc_sel_2_0(salloc_arb_io_in_2_bits_vc_sel_2_0),
    .io_in_2_bits_vc_sel_1_0(salloc_arb_io_in_2_bits_vc_sel_1_0),
    .io_in_2_bits_vc_sel_1_1(salloc_arb_io_in_2_bits_vc_sel_1_1),
    .io_in_2_bits_vc_sel_1_2(salloc_arb_io_in_2_bits_vc_sel_1_2),
    .io_in_2_bits_vc_sel_0_0(salloc_arb_io_in_2_bits_vc_sel_0_0),
    .io_in_2_bits_vc_sel_0_1(salloc_arb_io_in_2_bits_vc_sel_0_1),
    .io_in_2_bits_vc_sel_0_2(salloc_arb_io_in_2_bits_vc_sel_0_2),
    .io_in_2_bits_tail(salloc_arb_io_in_2_bits_tail),
    .io_in_3_ready(salloc_arb_io_in_3_ready),
    .io_in_3_valid(salloc_arb_io_in_3_valid),
    .io_in_3_bits_vc_sel_2_0(salloc_arb_io_in_3_bits_vc_sel_2_0),
    .io_in_3_bits_vc_sel_1_0(salloc_arb_io_in_3_bits_vc_sel_1_0),
    .io_in_3_bits_vc_sel_1_1(salloc_arb_io_in_3_bits_vc_sel_1_1),
    .io_in_3_bits_vc_sel_1_2(salloc_arb_io_in_3_bits_vc_sel_1_2),
    .io_in_3_bits_vc_sel_1_3(salloc_arb_io_in_3_bits_vc_sel_1_3),
    .io_in_3_bits_vc_sel_0_0(salloc_arb_io_in_3_bits_vc_sel_0_0),
    .io_in_3_bits_vc_sel_0_1(salloc_arb_io_in_3_bits_vc_sel_0_1),
    .io_in_3_bits_vc_sel_0_2(salloc_arb_io_in_3_bits_vc_sel_0_2),
    .io_in_3_bits_vc_sel_0_3(salloc_arb_io_in_3_bits_vc_sel_0_3),
    .io_in_3_bits_tail(salloc_arb_io_in_3_bits_tail),
    .io_out_0_ready(salloc_arb_io_out_0_ready),
    .io_out_0_valid(salloc_arb_io_out_0_valid),
    .io_out_0_bits_vc_sel_2_0(salloc_arb_io_out_0_bits_vc_sel_2_0),
    .io_out_0_bits_vc_sel_1_0(salloc_arb_io_out_0_bits_vc_sel_1_0),
    .io_out_0_bits_vc_sel_1_1(salloc_arb_io_out_0_bits_vc_sel_1_1),
    .io_out_0_bits_vc_sel_1_2(salloc_arb_io_out_0_bits_vc_sel_1_2),
    .io_out_0_bits_vc_sel_1_3(salloc_arb_io_out_0_bits_vc_sel_1_3),
    .io_out_0_bits_vc_sel_0_0(salloc_arb_io_out_0_bits_vc_sel_0_0),
    .io_out_0_bits_vc_sel_0_1(salloc_arb_io_out_0_bits_vc_sel_0_1),
    .io_out_0_bits_vc_sel_0_2(salloc_arb_io_out_0_bits_vc_sel_0_2),
    .io_out_0_bits_vc_sel_0_3(salloc_arb_io_out_0_bits_vc_sel_0_3),
    .io_out_0_bits_tail(salloc_arb_io_out_0_bits_tail),
    .io_chosen_oh_0(salloc_arb_io_chosen_oh_0)
  );
  assign io_router_req_valid = route_arbiter_io_out_valid; // @[InputUnit.scala 189:17]
  assign io_router_req_bits_src_virt_id = route_arbiter_io_out_bits_src_virt_id; // @[InputUnit.scala 189:17]
  assign io_router_req_bits_flow_ingress_node = route_arbiter_io_out_bits_flow_ingress_node; // @[InputUnit.scala 189:17]
  assign io_router_req_bits_flow_egress_node = route_arbiter_io_out_bits_flow_egress_node; // @[InputUnit.scala 189:17]
  assign io_vcalloc_req_valid = vcalloc_vals_0 | vcalloc_vals_1 | vcalloc_vals_2 | vcalloc_vals_3; // @[package.scala 73:59]
  assign io_vcalloc_req_bits_vc_sel_2_0 = vcalloc_sel[0] & states_0_vc_sel_2_0 | vcalloc_sel[1] & states_1_vc_sel_2_0 |
    vcalloc_sel[2] & states_2_vc_sel_2_0 | vcalloc_sel[3] & states_3_vc_sel_2_0; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_1_0 = vcalloc_sel[0] & states_0_vc_sel_1_0 | vcalloc_sel[1] & states_1_vc_sel_1_0 |
    vcalloc_sel[2] & states_2_vc_sel_1_0 | vcalloc_sel[3] & states_3_vc_sel_1_0; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_1_1 = vcalloc_sel[1] & states_1_vc_sel_1_1 | vcalloc_sel[2] & states_2_vc_sel_1_1 |
    vcalloc_sel[3] & states_3_vc_sel_1_1; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_1_2 = vcalloc_sel[2] & states_2_vc_sel_1_2 | vcalloc_sel[3] & states_3_vc_sel_1_2; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_1_3 = vcalloc_sel[3] & states_3_vc_sel_1_3; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_0_0 = vcalloc_sel[0] & states_0_vc_sel_0_0; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_0_1 = vcalloc_sel[1] & states_1_vc_sel_0_1 | vcalloc_sel[2] & states_2_vc_sel_0_1 |
    vcalloc_sel[3] & states_3_vc_sel_0_1; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_0_2 = vcalloc_sel[2] & states_2_vc_sel_0_2 | vcalloc_sel[3] & states_3_vc_sel_0_2; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_0_3 = vcalloc_sel[3] & states_3_vc_sel_0_3; // @[Mux.scala 27:73]
  assign io_salloc_req_0_valid = salloc_arb_io_out_0_valid; // @[InputUnit.scala 302:17 303:19 305:35]
  assign io_salloc_req_0_bits_vc_sel_2_0 = salloc_arb_io_out_0_bits_vc_sel_2_0; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_1_0 = salloc_arb_io_out_0_bits_vc_sel_1_0; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_1_1 = salloc_arb_io_out_0_bits_vc_sel_1_1; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_1_2 = salloc_arb_io_out_0_bits_vc_sel_1_2; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_1_3 = salloc_arb_io_out_0_bits_vc_sel_1_3; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_0_0 = salloc_arb_io_out_0_bits_vc_sel_0_0; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_0_1 = salloc_arb_io_out_0_bits_vc_sel_0_1; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_0_2 = salloc_arb_io_out_0_bits_vc_sel_0_2; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_0_3 = salloc_arb_io_out_0_bits_vc_sel_0_3; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_tail = salloc_arb_io_out_0_bits_tail; // @[InputUnit.scala 302:17]
  assign io_out_0_valid = salloc_outs_0_valid; // @[InputUnit.scala 349:21]
  assign io_out_0_bits_flit_head = salloc_outs_0_flit_head; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_flit_tail = salloc_outs_0_flit_tail; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_flit_payload = salloc_outs_0_flit_payload; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_flit_flow_ingress_node = salloc_outs_0_flit_flow_ingress_node; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_flit_flow_egress_node = salloc_outs_0_flit_flow_egress_node; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_out_virt_channel = salloc_outs_0_out_vid; // @[InputUnit.scala 351:37]
  assign io_debug_va_stall = _io_debug_va_stall_T_7[1:0]; // @[InputUnit.scala 266:21]
  assign io_debug_sa_stall = _io_debug_sa_stall_T_12[1:0]; // @[InputUnit.scala 301:21]
  assign io_in_credit_return = _io_in_credit_return_T ? salloc_arb_io_chosen_oh_0 : 4'h0; // @[InputUnit.scala 322:8]
  assign io_in_vc_free = _io_in_credit_return_T & _io_in_vc_free_T_11 ? salloc_arb_io_chosen_oh_0 : 4'h0; // @[InputUnit.scala 325:8]
  assign input_buffer_clock = clock;
  assign input_buffer_reset = reset;
  assign input_buffer_io_enq_0_valid = io_in_flit_0_valid; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_head = io_in_flit_0_bits_head; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_tail = io_in_flit_0_bits_tail; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_payload = io_in_flit_0_bits_payload; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_virt_channel_id = io_in_flit_0_bits_virt_channel_id; // @[InputUnit.scala 182:28]
  assign input_buffer_io_deq_0_ready = salloc_arb_io_in_0_ready; // @[InputUnit.scala 295:36]
  assign input_buffer_io_deq_1_ready = salloc_arb_io_in_1_ready; // @[InputUnit.scala 295:36]
  assign input_buffer_io_deq_2_ready = salloc_arb_io_in_2_ready; // @[InputUnit.scala 295:36]
  assign input_buffer_io_deq_3_ready = salloc_arb_io_in_3_ready; // @[InputUnit.scala 295:36]
  assign route_arbiter_io_in_0_valid = states_0_g == 3'h1; // @[InputUnit.scala 212:22]
  assign route_arbiter_io_in_0_bits_flow_ingress_node = states_0_flow_ingress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_0_bits_flow_egress_node = states_0_flow_egress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_1_valid = states_1_g == 3'h1; // @[InputUnit.scala 212:22]
  assign route_arbiter_io_in_1_bits_flow_ingress_node = states_1_flow_ingress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_1_bits_flow_egress_node = states_1_flow_egress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_2_valid = states_2_g == 3'h1; // @[InputUnit.scala 212:22]
  assign route_arbiter_io_in_2_bits_flow_ingress_node = states_2_flow_ingress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_2_bits_flow_egress_node = states_2_flow_egress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_3_valid = states_3_g == 3'h1; // @[InputUnit.scala 212:22]
  assign route_arbiter_io_in_3_bits_flow_ingress_node = states_3_flow_ingress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_3_bits_flow_egress_node = states_3_flow_egress_node; // @[InputUnit.scala 213:19]
  assign salloc_arb_clock = clock;
  assign salloc_arb_reset = reset;
  assign salloc_arb_io_in_0_valid = states_0_g == 3'h3 & credit_available & input_buffer_io_deq_0_valid; // @[InputUnit.scala 288:50]
  assign salloc_arb_io_in_0_bits_vc_sel_2_0 = states_0_vc_sel_2_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_0_bits_vc_sel_1_0 = states_0_vc_sel_1_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_0_bits_vc_sel_0_0 = states_0_vc_sel_0_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_0_bits_tail = input_buffer_io_deq_0_bits_tail; // @[InputUnit.scala 291:19]
  assign salloc_arb_io_in_1_valid = states_1_g == 3'h3 & credit_available_1 & input_buffer_io_deq_1_valid; // @[InputUnit.scala 288:50]
  assign salloc_arb_io_in_1_bits_vc_sel_2_0 = states_1_vc_sel_2_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_1_bits_vc_sel_1_0 = states_1_vc_sel_1_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_1_bits_vc_sel_1_1 = states_1_vc_sel_1_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_1_bits_vc_sel_0_0 = 1'h0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_1_bits_vc_sel_0_1 = states_1_vc_sel_0_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_1_bits_tail = input_buffer_io_deq_1_bits_tail; // @[InputUnit.scala 291:19]
  assign salloc_arb_io_in_2_valid = states_2_g == 3'h3 & credit_available_2 & input_buffer_io_deq_2_valid; // @[InputUnit.scala 288:50]
  assign salloc_arb_io_in_2_bits_vc_sel_2_0 = states_2_vc_sel_2_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_1_0 = states_2_vc_sel_1_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_1_1 = states_2_vc_sel_1_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_1_2 = states_2_vc_sel_1_2; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_0_0 = 1'h0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_0_1 = states_2_vc_sel_0_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_0_2 = states_2_vc_sel_0_2; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_tail = input_buffer_io_deq_2_bits_tail; // @[InputUnit.scala 291:19]
  assign salloc_arb_io_in_3_valid = states_3_g == 3'h3 & credit_available_3 & input_buffer_io_deq_3_valid; // @[InputUnit.scala 288:50]
  assign salloc_arb_io_in_3_bits_vc_sel_2_0 = states_3_vc_sel_2_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_1_0 = states_3_vc_sel_1_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_1_1 = states_3_vc_sel_1_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_1_2 = states_3_vc_sel_1_2; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_1_3 = states_3_vc_sel_1_3; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_0_0 = 1'h0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_0_1 = states_3_vc_sel_0_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_0_2 = states_3_vc_sel_0_2; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_0_3 = states_3_vc_sel_0_3; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_tail = input_buffer_io_deq_3_bits_tail; // @[InputUnit.scala 291:19]
  assign salloc_arb_io_out_0_ready = io_salloc_req_0_ready; // @[InputUnit.scala 302:17 303:19 304:39]
  always @(posedge clock) begin
    if (reset) begin // @[InputUnit.scala 377:23]
      states_0_g <= 3'h0; // @[InputUnit.scala 378:24]
    end else if (_T_60 & input_buffer_io_deq_0_bits_tail) begin // @[InputUnit.scala 292:35]
      states_0_g <= 3'h0; // @[InputUnit.scala 293:13]
    end else if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[0]) begin // @[InputUnit.scala 270:29]
        states_0_g <= 3'h3; // @[InputUnit.scala 272:21]
      end else begin
        states_0_g <= _GEN_222;
      end
    end else begin
      states_0_g <= _GEN_222;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[0]) begin // @[InputUnit.scala 270:29]
        states_0_vc_sel_2_0 <= io_vcalloc_resp_vc_sel_2_0; // @[InputUnit.scala 271:26]
      end else begin
        states_0_vc_sel_2_0 <= _GEN_184;
      end
    end else begin
      states_0_vc_sel_2_0 <= _GEN_184;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[0]) begin // @[InputUnit.scala 270:29]
        states_0_vc_sel_1_0 <= io_vcalloc_resp_vc_sel_1_0; // @[InputUnit.scala 271:26]
      end else begin
        states_0_vc_sel_1_0 <= _GEN_185;
      end
    end else begin
      states_0_vc_sel_1_0 <= _GEN_185;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[0]) begin // @[InputUnit.scala 270:29]
        states_0_vc_sel_0_0 <= io_vcalloc_resp_vc_sel_0_0; // @[InputUnit.scala 271:26]
      end else begin
        states_0_vc_sel_0_0 <= _GEN_189;
      end
    end else begin
      states_0_vc_sel_0_0 <= _GEN_189;
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h0 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_0_flow_ingress_node <= io_in_flit_0_bits_flow_ingress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h0 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_0_flow_egress_node <= io_in_flit_0_bits_flow_egress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (reset) begin // @[InputUnit.scala 377:23]
      states_1_g <= 3'h0; // @[InputUnit.scala 378:24]
    end else if (_T_62 & input_buffer_io_deq_1_bits_tail) begin // @[InputUnit.scala 292:35]
      states_1_g <= 3'h0; // @[InputUnit.scala 293:13]
    end else if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_g <= 3'h3; // @[InputUnit.scala 272:21]
      end else begin
        states_1_g <= _GEN_223;
      end
    end else begin
      states_1_g <= _GEN_223;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_vc_sel_2_0 <= io_vcalloc_resp_vc_sel_2_0; // @[InputUnit.scala 271:26]
      end else begin
        states_1_vc_sel_2_0 <= _GEN_193;
      end
    end else begin
      states_1_vc_sel_2_0 <= _GEN_193;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_vc_sel_1_0 <= io_vcalloc_resp_vc_sel_1_0; // @[InputUnit.scala 271:26]
      end else begin
        states_1_vc_sel_1_0 <= _GEN_194;
      end
    end else begin
      states_1_vc_sel_1_0 <= _GEN_194;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_vc_sel_1_1 <= io_vcalloc_resp_vc_sel_1_1; // @[InputUnit.scala 271:26]
      end else begin
        states_1_vc_sel_1_1 <= _GEN_195;
      end
    end else begin
      states_1_vc_sel_1_1 <= _GEN_195;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_vc_sel_0_1 <= io_vcalloc_resp_vc_sel_0_1; // @[InputUnit.scala 271:26]
      end else begin
        states_1_vc_sel_0_1 <= _GEN_199;
      end
    end else begin
      states_1_vc_sel_0_1 <= _GEN_199;
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h1 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_1_flow_ingress_node <= io_in_flit_0_bits_flow_ingress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h1 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_1_flow_egress_node <= io_in_flit_0_bits_flow_egress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (reset) begin // @[InputUnit.scala 377:23]
      states_2_g <= 3'h0; // @[InputUnit.scala 378:24]
    end else if (_T_64 & input_buffer_io_deq_2_bits_tail) begin // @[InputUnit.scala 292:35]
      states_2_g <= 3'h0; // @[InputUnit.scala 293:13]
    end else if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_g <= 3'h3; // @[InputUnit.scala 272:21]
      end else begin
        states_2_g <= _GEN_224;
      end
    end else begin
      states_2_g <= _GEN_224;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_2_0 <= io_vcalloc_resp_vc_sel_2_0; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_2_0 <= _GEN_202;
      end
    end else begin
      states_2_vc_sel_2_0 <= _GEN_202;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_1_0 <= io_vcalloc_resp_vc_sel_1_0; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_1_0 <= _GEN_203;
      end
    end else begin
      states_2_vc_sel_1_0 <= _GEN_203;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_1_1 <= io_vcalloc_resp_vc_sel_1_1; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_1_1 <= _GEN_204;
      end
    end else begin
      states_2_vc_sel_1_1 <= _GEN_204;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_1_2 <= io_vcalloc_resp_vc_sel_1_2; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_1_2 <= _GEN_205;
      end
    end else begin
      states_2_vc_sel_1_2 <= _GEN_205;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_0_1 <= io_vcalloc_resp_vc_sel_0_1; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_0_1 <= _GEN_208;
      end
    end else begin
      states_2_vc_sel_0_1 <= _GEN_208;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_0_2 <= io_vcalloc_resp_vc_sel_0_2; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_0_2 <= _GEN_209;
      end
    end else begin
      states_2_vc_sel_0_2 <= _GEN_209;
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h2 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_2_flow_ingress_node <= io_in_flit_0_bits_flow_ingress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h2 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_2_flow_egress_node <= io_in_flit_0_bits_flow_egress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (reset) begin // @[InputUnit.scala 377:23]
      states_3_g <= 3'h0; // @[InputUnit.scala 378:24]
    end else if (_T_66 & input_buffer_io_deq_3_bits_tail) begin // @[InputUnit.scala 292:35]
      states_3_g <= 3'h0; // @[InputUnit.scala 293:13]
    end else if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_g <= 3'h3; // @[InputUnit.scala 272:21]
      end else begin
        states_3_g <= _GEN_225;
      end
    end else begin
      states_3_g <= _GEN_225;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_2_0 <= io_vcalloc_resp_vc_sel_2_0; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_2_0 <= _GEN_211;
      end
    end else begin
      states_3_vc_sel_2_0 <= _GEN_211;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_1_0 <= io_vcalloc_resp_vc_sel_1_0; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_1_0 <= _GEN_212;
      end
    end else begin
      states_3_vc_sel_1_0 <= _GEN_212;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_1_1 <= io_vcalloc_resp_vc_sel_1_1; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_1_1 <= _GEN_213;
      end
    end else begin
      states_3_vc_sel_1_1 <= _GEN_213;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_1_2 <= io_vcalloc_resp_vc_sel_1_2; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_1_2 <= _GEN_214;
      end
    end else begin
      states_3_vc_sel_1_2 <= _GEN_214;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_1_3 <= io_vcalloc_resp_vc_sel_1_3; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_1_3 <= _GEN_215;
      end
    end else begin
      states_3_vc_sel_1_3 <= _GEN_215;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_0_1 <= io_vcalloc_resp_vc_sel_0_1; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_0_1 <= _GEN_217;
      end
    end else begin
      states_3_vc_sel_0_1 <= _GEN_217;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_0_2 <= io_vcalloc_resp_vc_sel_0_2; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_0_2 <= _GEN_218;
      end
    end else begin
      states_3_vc_sel_0_2 <= _GEN_218;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_0_3 <= io_vcalloc_resp_vc_sel_0_3; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_0_3 <= _GEN_219;
      end
    end else begin
      states_3_vc_sel_0_3 <= _GEN_219;
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h3 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_3_flow_ingress_node <= io_in_flit_0_bits_flow_ingress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h3 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_3_flow_egress_node <= io_in_flit_0_bits_flow_egress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (reset) begin // @[InputUnit.scala 233:21]
      mask <= 4'h0; // @[InputUnit.scala 233:21]
    end else if (io_router_req_valid) begin // @[InputUnit.scala 239:31]
      mask <= _mask_T_2; // @[InputUnit.scala 240:10]
    end else if (_T_26) begin // @[InputUnit.scala 241:34]
      mask <= _mask_T_17; // @[InputUnit.scala 242:10]
    end
    salloc_outs_0_valid <= salloc_arb_io_out_0_ready & salloc_arb_io_out_0_valid; // @[Decoupled.scala 51:35]
    salloc_outs_0_out_vid <= _virt_channel_T_10 | _virt_channel_T_11; // @[Mux.scala 27:73]
    salloc_outs_0_flit_head <= salloc_arb_io_chosen_oh_0[0] & input_buffer_io_deq_0_bits_head |
      salloc_arb_io_chosen_oh_0[1] & input_buffer_io_deq_1_bits_head | salloc_arb_io_chosen_oh_0[2] &
      input_buffer_io_deq_2_bits_head | salloc_arb_io_chosen_oh_0[3] & input_buffer_io_deq_3_bits_head; // @[Mux.scala 27:73]
    salloc_outs_0_flit_tail <= salloc_arb_io_chosen_oh_0[0] & input_buffer_io_deq_0_bits_tail |
      salloc_arb_io_chosen_oh_0[1] & input_buffer_io_deq_1_bits_tail | salloc_arb_io_chosen_oh_0[2] &
      input_buffer_io_deq_2_bits_tail | salloc_arb_io_chosen_oh_0[3] & input_buffer_io_deq_3_bits_tail; // @[Mux.scala 27:73]
    salloc_outs_0_flit_payload <= _salloc_outs_0_flit_payload_T_9 | _salloc_outs_0_flit_payload_T_7; // @[Mux.scala 27:73]
    salloc_outs_0_flit_flow_ingress_node <= _salloc_outs_0_flit_flow_T_30 | _salloc_outs_0_flit_flow_T_28; // @[Mux.scala 27:73]
    salloc_outs_0_flit_flow_egress_node <= _salloc_outs_0_flit_flow_T_16 | _salloc_outs_0_flit_flow_T_14; // @[Mux.scala 27:73]
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T & _T_3 & ~(_GEN_3 == 3'h0)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:197 assert(states(id).g === g_i)\n"); // @[InputUnit.scala 197:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_router_req_valid & _T_3 & ~(_GEN_139 == 3'h1)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:224 assert(states(id).g === g_r)\n"); // @[InputUnit.scala 224:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_39 & vcalloc_sel[0] & _T_3 & ~vcalloc_vals_0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:274 assert(states(i).g === g_v)\n"); // @[InputUnit.scala 274:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_39 & vcalloc_sel[1] & _T_3 & ~vcalloc_vals_1) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:274 assert(states(i).g === g_v)\n"); // @[InputUnit.scala 274:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_39 & vcalloc_sel[2] & _T_3 & ~vcalloc_vals_2) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:274 assert(states(i).g === g_v)\n"); // @[InputUnit.scala 274:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_39 & vcalloc_sel[3] & _T_3 & ~vcalloc_vals_3) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:274 assert(states(i).g === g_v)\n"); // @[InputUnit.scala 274:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  states_0_g = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  states_0_vc_sel_2_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  states_0_vc_sel_1_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  states_0_vc_sel_0_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  states_0_flow_ingress_node = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  states_0_flow_egress_node = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  states_1_g = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  states_1_vc_sel_2_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  states_1_vc_sel_1_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  states_1_vc_sel_1_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  states_1_vc_sel_0_1 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  states_1_flow_ingress_node = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  states_1_flow_egress_node = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  states_2_g = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  states_2_vc_sel_2_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  states_2_vc_sel_1_0 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  states_2_vc_sel_1_1 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  states_2_vc_sel_1_2 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  states_2_vc_sel_0_1 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  states_2_vc_sel_0_2 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  states_2_flow_ingress_node = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  states_2_flow_egress_node = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  states_3_g = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  states_3_vc_sel_2_0 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  states_3_vc_sel_1_0 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  states_3_vc_sel_1_1 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  states_3_vc_sel_1_2 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  states_3_vc_sel_1_3 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  states_3_vc_sel_0_1 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  states_3_vc_sel_0_2 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  states_3_vc_sel_0_3 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  states_3_flow_ingress_node = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  states_3_flow_egress_node = _RAND_32[1:0];
  _RAND_33 = {1{`RANDOM}};
  mask = _RAND_33[3:0];
  _RAND_34 = {1{`RANDOM}};
  salloc_outs_0_valid = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  salloc_outs_0_out_vid = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  salloc_outs_0_flit_head = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  salloc_outs_0_flit_tail = _RAND_37[0:0];
  _RAND_38 = {2{`RANDOM}};
  salloc_outs_0_flit_payload = _RAND_38[63:0];
  _RAND_39 = {1{`RANDOM}};
  salloc_outs_0_flit_flow_ingress_node = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  salloc_outs_0_flit_flow_egress_node = _RAND_40[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (_T & ~reset) begin
      assert(1'h1); // @[InputUnit.scala 196:13]
    end
    //
    if (_T & _T_3) begin
      assert(_GEN_3 == 3'h0); // @[InputUnit.scala 197:13]
    end
    //
    if (io_router_req_valid & _T_3) begin
      assert(_GEN_139 == 3'h1); // @[InputUnit.scala 224:11]
    end
    //
    if (_T_39 & vcalloc_sel[0] & _T_3) begin
      assert(vcalloc_vals_0); // @[InputUnit.scala 274:17]
    end
    //
    if (_T_39 & vcalloc_sel[1] & _T_3) begin
      assert(vcalloc_vals_1); // @[InputUnit.scala 274:17]
    end
    //
    if (_T_39 & vcalloc_sel[2] & _T_3) begin
      assert(vcalloc_vals_2); // @[InputUnit.scala 274:17]
    end
    //
    if (_T_39 & vcalloc_sel[3] & _T_3) begin
      assert(vcalloc_vals_3); // @[InputUnit.scala 274:17]
    end
  end
endmodule
module InputUnit_5(
  input         clock,
  input         reset,
  output        io_router_req_valid,
  output [1:0]  io_router_req_bits_src_virt_id,
  output [1:0]  io_router_req_bits_flow_ingress_node,
  output [1:0]  io_router_req_bits_flow_egress_node,
  input         io_router_resp_vc_sel_1_0,
  input         io_router_resp_vc_sel_1_1,
  input         io_router_resp_vc_sel_1_2,
  input         io_router_resp_vc_sel_1_3,
  input         io_router_resp_vc_sel_0_0,
  input         io_router_resp_vc_sel_0_1,
  input         io_router_resp_vc_sel_0_2,
  input         io_router_resp_vc_sel_0_3,
  input         io_vcalloc_req_ready,
  output        io_vcalloc_req_valid,
  output        io_vcalloc_req_bits_vc_sel_2_0,
  output        io_vcalloc_req_bits_vc_sel_1_0,
  output        io_vcalloc_req_bits_vc_sel_1_1,
  output        io_vcalloc_req_bits_vc_sel_1_2,
  output        io_vcalloc_req_bits_vc_sel_1_3,
  output        io_vcalloc_req_bits_vc_sel_0_0,
  output        io_vcalloc_req_bits_vc_sel_0_1,
  output        io_vcalloc_req_bits_vc_sel_0_2,
  output        io_vcalloc_req_bits_vc_sel_0_3,
  input         io_vcalloc_resp_vc_sel_2_0,
  input         io_vcalloc_resp_vc_sel_1_0,
  input         io_vcalloc_resp_vc_sel_1_1,
  input         io_vcalloc_resp_vc_sel_1_2,
  input         io_vcalloc_resp_vc_sel_1_3,
  input         io_vcalloc_resp_vc_sel_0_0,
  input         io_vcalloc_resp_vc_sel_0_1,
  input         io_vcalloc_resp_vc_sel_0_2,
  input         io_vcalloc_resp_vc_sel_0_3,
  input         io_out_credit_available_2_0,
  input         io_out_credit_available_1_0,
  input         io_out_credit_available_1_1,
  input         io_out_credit_available_1_2,
  input         io_out_credit_available_1_3,
  input         io_out_credit_available_0_0,
  input         io_out_credit_available_0_1,
  input         io_out_credit_available_0_2,
  input         io_out_credit_available_0_3,
  input         io_salloc_req_0_ready,
  output        io_salloc_req_0_valid,
  output        io_salloc_req_0_bits_vc_sel_2_0,
  output        io_salloc_req_0_bits_vc_sel_1_0,
  output        io_salloc_req_0_bits_vc_sel_1_1,
  output        io_salloc_req_0_bits_vc_sel_1_2,
  output        io_salloc_req_0_bits_vc_sel_1_3,
  output        io_salloc_req_0_bits_vc_sel_0_0,
  output        io_salloc_req_0_bits_vc_sel_0_1,
  output        io_salloc_req_0_bits_vc_sel_0_2,
  output        io_salloc_req_0_bits_vc_sel_0_3,
  output        io_salloc_req_0_bits_tail,
  output        io_out_0_valid,
  output        io_out_0_bits_flit_head,
  output        io_out_0_bits_flit_tail,
  output [63:0] io_out_0_bits_flit_payload,
  output [1:0]  io_out_0_bits_flit_flow_ingress_node,
  output [1:0]  io_out_0_bits_flit_flow_egress_node,
  output [1:0]  io_out_0_bits_out_virt_channel,
  output [1:0]  io_debug_va_stall,
  output [1:0]  io_debug_sa_stall,
  input         io_in_flit_0_valid,
  input         io_in_flit_0_bits_head,
  input         io_in_flit_0_bits_tail,
  input  [63:0] io_in_flit_0_bits_payload,
  input  [1:0]  io_in_flit_0_bits_flow_ingress_node,
  input  [1:0]  io_in_flit_0_bits_flow_egress_node,
  input  [1:0]  io_in_flit_0_bits_virt_channel_id,
  output [3:0]  io_in_credit_return,
  output [3:0]  io_in_vc_free
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
`endif // RANDOMIZE_REG_INIT
  wire  input_buffer_clock; // @[InputUnit.scala 180:28]
  wire  input_buffer_reset; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_enq_0_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_enq_0_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_enq_0_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_enq_0_bits_payload; // @[InputUnit.scala 180:28]
  wire [1:0] input_buffer_io_enq_0_bits_virt_channel_id; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_0_ready; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_0_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_0_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_0_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_deq_0_bits_payload; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_ready; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_deq_1_bits_payload; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_ready; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_deq_2_bits_payload; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_3_ready; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_3_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_3_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_3_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_deq_3_bits_payload; // @[InputUnit.scala 180:28]
  wire  route_arbiter_io_in_0_valid; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_0_bits_flow_ingress_node; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_0_bits_flow_egress_node; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_1_ready; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_1_valid; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_1_bits_flow_ingress_node; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_1_bits_flow_egress_node; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_2_ready; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_2_valid; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_2_bits_flow_ingress_node; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_2_bits_flow_egress_node; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_3_ready; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_3_valid; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_3_bits_flow_ingress_node; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_3_bits_flow_egress_node; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_out_valid; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_out_bits_src_virt_id; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_out_bits_flow_ingress_node; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_out_bits_flow_egress_node; // @[InputUnit.scala 186:29]
  wire  salloc_arb_clock; // @[InputUnit.scala 279:26]
  wire  salloc_arb_reset; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_bits_vc_sel_2_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_bits_vc_sel_1_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_bits_tail; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_vc_sel_2_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_vc_sel_1_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_vc_sel_1_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_vc_sel_0_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_tail; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_2_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_1_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_1_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_1_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_0_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_0_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_tail; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_2_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_1_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_1_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_1_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_1_3; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_0_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_0_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_0_3; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_tail; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_2_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_1_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_1_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_1_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_1_3; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_0_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_0_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_0_3; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_tail; // @[InputUnit.scala 279:26]
  wire [3:0] salloc_arb_io_chosen_oh_0; // @[InputUnit.scala 279:26]
  reg [2:0] states_0_g; // @[InputUnit.scala 191:19]
  reg  states_0_vc_sel_2_0; // @[InputUnit.scala 191:19]
  reg  states_0_vc_sel_1_0; // @[InputUnit.scala 191:19]
  reg  states_0_vc_sel_0_0; // @[InputUnit.scala 191:19]
  reg [1:0] states_0_flow_ingress_node; // @[InputUnit.scala 191:19]
  reg [1:0] states_0_flow_egress_node; // @[InputUnit.scala 191:19]
  reg [2:0] states_1_g; // @[InputUnit.scala 191:19]
  reg  states_1_vc_sel_2_0; // @[InputUnit.scala 191:19]
  reg  states_1_vc_sel_1_1; // @[InputUnit.scala 191:19]
  reg  states_1_vc_sel_0_0; // @[InputUnit.scala 191:19]
  reg  states_1_vc_sel_0_1; // @[InputUnit.scala 191:19]
  reg [1:0] states_1_flow_ingress_node; // @[InputUnit.scala 191:19]
  reg [1:0] states_1_flow_egress_node; // @[InputUnit.scala 191:19]
  reg [2:0] states_2_g; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_2_0; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_1_1; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_1_2; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_0_0; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_0_1; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_0_2; // @[InputUnit.scala 191:19]
  reg [1:0] states_2_flow_ingress_node; // @[InputUnit.scala 191:19]
  reg [1:0] states_2_flow_egress_node; // @[InputUnit.scala 191:19]
  reg [2:0] states_3_g; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_2_0; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_1_1; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_1_2; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_1_3; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_0_0; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_0_1; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_0_2; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_0_3; // @[InputUnit.scala 191:19]
  reg [1:0] states_3_flow_ingress_node; // @[InputUnit.scala 191:19]
  reg [1:0] states_3_flow_egress_node; // @[InputUnit.scala 191:19]
  wire  _T = io_in_flit_0_valid & io_in_flit_0_bits_head; // @[InputUnit.scala 194:32]
  wire  _T_3 = ~reset; // @[InputUnit.scala 196:13]
  wire [2:0] _GEN_1 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? states_1_g : states_0_g; // @[InputUnit.scala 197:{27,27}]
  wire [2:0] _GEN_2 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? states_2_g : _GEN_1; // @[InputUnit.scala 197:{27,27}]
  wire [2:0] _GEN_3 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? states_3_g : _GEN_2; // @[InputUnit.scala 197:{27,27}]
  wire  at_dest = io_in_flit_0_bits_flow_egress_node == 2'h2; // @[InputUnit.scala 198:57]
  wire [2:0] _states_g_T = at_dest ? 3'h2 : 3'h1; // @[InputUnit.scala 199:26]
  wire [2:0] _GEN_4 = 2'h0 == io_in_flit_0_bits_virt_channel_id ? _states_g_T : states_0_g; // @[InputUnit.scala 191:19 199:{20,20}]
  wire [2:0] _GEN_5 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? _states_g_T : states_1_g; // @[InputUnit.scala 191:19 199:{20,20}]
  wire [2:0] _GEN_6 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? _states_g_T : states_2_g; // @[InputUnit.scala 191:19 199:{20,20}]
  wire [2:0] _GEN_7 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? _states_g_T : states_3_g; // @[InputUnit.scala 191:19 199:{20,20}]
  wire  _GEN_8 = 2'h0 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_0_vc_sel_0_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_9 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_1_vc_sel_0_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_10 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_0_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_11 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_0_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_13 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_1_vc_sel_0_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_14 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_0_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_15 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_0_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_18 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_0_2; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_19 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_0_2; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_23 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_0_3; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_24 = 2'h0 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_0_vc_sel_1_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_29 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_1_vc_sel_1_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_30 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_1_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_31 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_1_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_34 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_1_2; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_35 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_1_2; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_39 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_1_3; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_40 = 2'h0 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_0_vc_sel_2_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_41 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_1_vc_sel_2_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_42 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_2_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_43 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_2_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_44 = 2'h0 == io_in_flit_0_bits_virt_channel_id | _GEN_40; // @[InputUnit.scala 203:{44,44}]
  wire  _GEN_45 = 2'h1 == io_in_flit_0_bits_virt_channel_id | _GEN_41; // @[InputUnit.scala 203:{44,44}]
  wire  _GEN_46 = 2'h2 == io_in_flit_0_bits_virt_channel_id | _GEN_42; // @[InputUnit.scala 203:{44,44}]
  wire  _GEN_47 = 2'h3 == io_in_flit_0_bits_virt_channel_id | _GEN_43; // @[InputUnit.scala 203:{44,44}]
  wire [2:0] _GEN_72 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_4 : states_0_g; // @[InputUnit.scala 191:19 194:60]
  wire [2:0] _GEN_73 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_5 : states_1_g; // @[InputUnit.scala 191:19 194:60]
  wire [2:0] _GEN_74 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_6 : states_2_g; // @[InputUnit.scala 191:19 194:60]
  wire [2:0] _GEN_75 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_7 : states_3_g; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_76 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_8 : states_0_vc_sel_0_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_77 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_9 : states_1_vc_sel_0_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_78 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_10 : states_2_vc_sel_0_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_79 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_11 : states_3_vc_sel_0_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_81 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_13 : states_1_vc_sel_0_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_82 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_14 : states_2_vc_sel_0_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_83 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_15 : states_3_vc_sel_0_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_86 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_18 : states_2_vc_sel_0_2; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_87 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_19 : states_3_vc_sel_0_2; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_91 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_23 : states_3_vc_sel_0_3; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_92 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_24 : states_0_vc_sel_1_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_97 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_29 : states_1_vc_sel_1_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_98 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_30 : states_2_vc_sel_1_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_99 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_31 : states_3_vc_sel_1_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_102 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_34 : states_2_vc_sel_1_2; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_103 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_35 : states_3_vc_sel_1_2; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_107 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_39 : states_3_vc_sel_1_3; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_108 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_44 : states_0_vc_sel_2_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_109 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_45 : states_1_vc_sel_2_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_110 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_46 : states_2_vc_sel_2_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_111 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_47 : states_3_vc_sel_2_0; // @[InputUnit.scala 191:19 194:60]
  wire  _T_10 = route_arbiter_io_in_0_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_132 = _T_10 ? 3'h2 : _GEN_72; // @[InputUnit.scala 215:{23,29}]
  wire  _T_11 = route_arbiter_io_in_1_ready & route_arbiter_io_in_1_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_133 = _T_11 ? 3'h2 : _GEN_73; // @[InputUnit.scala 215:{23,29}]
  wire  _T_12 = route_arbiter_io_in_2_ready & route_arbiter_io_in_2_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_134 = _T_12 ? 3'h2 : _GEN_74; // @[InputUnit.scala 215:{23,29}]
  wire  _T_13 = route_arbiter_io_in_3_ready & route_arbiter_io_in_3_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_135 = _T_13 ? 3'h2 : _GEN_75; // @[InputUnit.scala 215:{23,29}]
  wire [2:0] _GEN_137 = 2'h1 == io_router_req_bits_src_virt_id ? states_1_g : states_0_g; // @[InputUnit.scala 224:{25,25}]
  wire [2:0] _GEN_138 = 2'h2 == io_router_req_bits_src_virt_id ? states_2_g : _GEN_137; // @[InputUnit.scala 224:{25,25}]
  wire [2:0] _GEN_139 = 2'h3 == io_router_req_bits_src_virt_id ? states_3_g : _GEN_138; // @[InputUnit.scala 224:{25,25}]
  wire [2:0] _GEN_140 = 2'h0 == io_router_req_bits_src_virt_id ? 3'h2 : _GEN_132; // @[InputUnit.scala 225:{18,18}]
  wire [2:0] _GEN_141 = 2'h1 == io_router_req_bits_src_virt_id ? 3'h2 : _GEN_133; // @[InputUnit.scala 225:{18,18}]
  wire [2:0] _GEN_142 = 2'h2 == io_router_req_bits_src_virt_id ? 3'h2 : _GEN_134; // @[InputUnit.scala 225:{18,18}]
  wire [2:0] _GEN_143 = 2'h3 == io_router_req_bits_src_virt_id ? 3'h2 : _GEN_135; // @[InputUnit.scala 225:{18,18}]
  wire  _GEN_144 = 2'h0 == io_router_req_bits_src_virt_id ? 1'h0 : _GEN_108; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_145 = 2'h0 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_0 : _GEN_92; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_149 = 2'h0 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_0 : _GEN_76; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_153 = 2'h1 == io_router_req_bits_src_virt_id ? 1'h0 : _GEN_109; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_155 = 2'h1 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_1 : _GEN_97; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_158 = 2'h1 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_0 : _GEN_77; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_159 = 2'h1 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_1 : _GEN_81; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_162 = 2'h2 == io_router_req_bits_src_virt_id ? 1'h0 : _GEN_110; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_164 = 2'h2 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_1 : _GEN_98; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_165 = 2'h2 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_2 : _GEN_102; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_167 = 2'h2 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_0 : _GEN_78; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_168 = 2'h2 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_1 : _GEN_82; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_169 = 2'h2 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_2 : _GEN_86; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_171 = 2'h3 == io_router_req_bits_src_virt_id ? 1'h0 : _GEN_111; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_173 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_1 : _GEN_99; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_174 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_2 : _GEN_103; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_175 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_3 : _GEN_107; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_176 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_0 : _GEN_79; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_177 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_1 : _GEN_83; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_178 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_2 : _GEN_87; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_179 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_3 : _GEN_91; // @[InputUnit.scala 227:25 228:26]
  wire [2:0] _GEN_180 = io_router_req_valid ? _GEN_140 : _GEN_132; // @[InputUnit.scala 222:31]
  wire [2:0] _GEN_181 = io_router_req_valid ? _GEN_141 : _GEN_133; // @[InputUnit.scala 222:31]
  wire [2:0] _GEN_182 = io_router_req_valid ? _GEN_142 : _GEN_134; // @[InputUnit.scala 222:31]
  wire [2:0] _GEN_183 = io_router_req_valid ? _GEN_143 : _GEN_135; // @[InputUnit.scala 222:31]
  wire  _GEN_184 = io_router_req_valid ? _GEN_144 : _GEN_108; // @[InputUnit.scala 222:31]
  wire  _GEN_185 = io_router_req_valid ? _GEN_145 : _GEN_92; // @[InputUnit.scala 222:31]
  wire  _GEN_189 = io_router_req_valid ? _GEN_149 : _GEN_76; // @[InputUnit.scala 222:31]
  wire  _GEN_193 = io_router_req_valid ? _GEN_153 : _GEN_109; // @[InputUnit.scala 222:31]
  wire  _GEN_195 = io_router_req_valid ? _GEN_155 : _GEN_97; // @[InputUnit.scala 222:31]
  wire  _GEN_198 = io_router_req_valid ? _GEN_158 : _GEN_77; // @[InputUnit.scala 222:31]
  wire  _GEN_199 = io_router_req_valid ? _GEN_159 : _GEN_81; // @[InputUnit.scala 222:31]
  wire  _GEN_202 = io_router_req_valid ? _GEN_162 : _GEN_110; // @[InputUnit.scala 222:31]
  wire  _GEN_204 = io_router_req_valid ? _GEN_164 : _GEN_98; // @[InputUnit.scala 222:31]
  wire  _GEN_205 = io_router_req_valid ? _GEN_165 : _GEN_102; // @[InputUnit.scala 222:31]
  wire  _GEN_207 = io_router_req_valid ? _GEN_167 : _GEN_78; // @[InputUnit.scala 222:31]
  wire  _GEN_208 = io_router_req_valid ? _GEN_168 : _GEN_82; // @[InputUnit.scala 222:31]
  wire  _GEN_209 = io_router_req_valid ? _GEN_169 : _GEN_86; // @[InputUnit.scala 222:31]
  wire  _GEN_211 = io_router_req_valid ? _GEN_171 : _GEN_111; // @[InputUnit.scala 222:31]
  wire  _GEN_213 = io_router_req_valid ? _GEN_173 : _GEN_99; // @[InputUnit.scala 222:31]
  wire  _GEN_214 = io_router_req_valid ? _GEN_174 : _GEN_103; // @[InputUnit.scala 222:31]
  wire  _GEN_215 = io_router_req_valid ? _GEN_175 : _GEN_107; // @[InputUnit.scala 222:31]
  wire  _GEN_216 = io_router_req_valid ? _GEN_176 : _GEN_79; // @[InputUnit.scala 222:31]
  wire  _GEN_217 = io_router_req_valid ? _GEN_177 : _GEN_83; // @[InputUnit.scala 222:31]
  wire  _GEN_218 = io_router_req_valid ? _GEN_178 : _GEN_87; // @[InputUnit.scala 222:31]
  wire  _GEN_219 = io_router_req_valid ? _GEN_179 : _GEN_91; // @[InputUnit.scala 222:31]
  reg [3:0] mask; // @[InputUnit.scala 233:21]
  wire  vcalloc_vals_1 = states_1_g == 3'h2; // @[InputUnit.scala 249:32]
  wire  vcalloc_vals_0 = states_0_g == 3'h2; // @[InputUnit.scala 249:32]
  wire  vcalloc_vals_3 = states_3_g == 3'h2; // @[InputUnit.scala 249:32]
  wire  vcalloc_vals_2 = states_2_g == 3'h2; // @[InputUnit.scala 249:32]
  wire [3:0] _vcalloc_filter_T = {vcalloc_vals_3,vcalloc_vals_2,vcalloc_vals_1,vcalloc_vals_0}; // @[InputUnit.scala 236:59]
  wire [3:0] _vcalloc_filter_T_2 = ~mask; // @[InputUnit.scala 236:89]
  wire [3:0] _vcalloc_filter_T_3 = _vcalloc_filter_T & _vcalloc_filter_T_2; // @[InputUnit.scala 236:87]
  wire [7:0] _vcalloc_filter_T_4 = {vcalloc_vals_3,vcalloc_vals_2,vcalloc_vals_1,vcalloc_vals_0,_vcalloc_filter_T_3}; // @[Cat.scala 33:92]
  wire [7:0] _vcalloc_filter_T_13 = _vcalloc_filter_T_4[7] ? 8'h80 : 8'h0; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_14 = _vcalloc_filter_T_4[6] ? 8'h40 : _vcalloc_filter_T_13; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_15 = _vcalloc_filter_T_4[5] ? 8'h20 : _vcalloc_filter_T_14; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_16 = _vcalloc_filter_T_4[4] ? 8'h10 : _vcalloc_filter_T_15; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_17 = _vcalloc_filter_T_4[3] ? 8'h8 : _vcalloc_filter_T_16; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_18 = _vcalloc_filter_T_4[2] ? 8'h4 : _vcalloc_filter_T_17; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_19 = _vcalloc_filter_T_4[1] ? 8'h2 : _vcalloc_filter_T_18; // @[Mux.scala 47:70]
  wire [7:0] vcalloc_filter = _vcalloc_filter_T_4[0] ? 8'h1 : _vcalloc_filter_T_19; // @[Mux.scala 47:70]
  wire [3:0] vcalloc_sel = vcalloc_filter[3:0] | vcalloc_filter[7:4]; // @[InputUnit.scala 237:58]
  wire [3:0] _mask_T = 4'h1 << io_router_req_bits_src_virt_id; // @[InputUnit.scala 240:18]
  wire [3:0] _mask_T_2 = _mask_T - 4'h1; // @[InputUnit.scala 240:53]
  wire  _T_26 = vcalloc_vals_0 | vcalloc_vals_1 | vcalloc_vals_2 | vcalloc_vals_3; // @[package.scala 73:59]
  wire [1:0] _mask_T_12 = vcalloc_sel[1] ? 2'h3 : 2'h0; // @[Mux.scala 27:73]
  wire [2:0] _mask_T_13 = vcalloc_sel[2] ? 3'h7 : 3'h0; // @[Mux.scala 27:73]
  wire [3:0] _mask_T_14 = vcalloc_sel[3] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [1:0] _GEN_60 = {{1'd0}, vcalloc_sel[0]}; // @[Mux.scala 27:73]
  wire [1:0] _mask_T_15 = _GEN_60 | _mask_T_12; // @[Mux.scala 27:73]
  wire [2:0] _GEN_61 = {{1'd0}, _mask_T_15}; // @[Mux.scala 27:73]
  wire [2:0] _mask_T_16 = _GEN_61 | _mask_T_13; // @[Mux.scala 27:73]
  wire [3:0] _GEN_62 = {{1'd0}, _mask_T_16}; // @[Mux.scala 27:73]
  wire [3:0] _mask_T_17 = _GEN_62 | _mask_T_14; // @[Mux.scala 27:73]
  wire [2:0] _GEN_222 = vcalloc_vals_0 & vcalloc_sel[0] & io_vcalloc_req_ready ? 3'h3 : _GEN_180; // @[InputUnit.scala 253:{76,82}]
  wire [2:0] _GEN_223 = vcalloc_vals_1 & vcalloc_sel[1] & io_vcalloc_req_ready ? 3'h3 : _GEN_181; // @[InputUnit.scala 253:{76,82}]
  wire [2:0] _GEN_224 = vcalloc_vals_2 & vcalloc_sel[2] & io_vcalloc_req_ready ? 3'h3 : _GEN_182; // @[InputUnit.scala 253:{76,82}]
  wire [2:0] _GEN_225 = vcalloc_vals_3 & vcalloc_sel[3] & io_vcalloc_req_ready ? 3'h3 : _GEN_183; // @[InputUnit.scala 253:{76,82}]
  wire [1:0] _io_debug_va_stall_T = vcalloc_vals_0 + vcalloc_vals_1; // @[Bitwise.scala 51:90]
  wire [1:0] _io_debug_va_stall_T_2 = vcalloc_vals_2 + vcalloc_vals_3; // @[Bitwise.scala 51:90]
  wire [2:0] _io_debug_va_stall_T_4 = _io_debug_va_stall_T + _io_debug_va_stall_T_2; // @[Bitwise.scala 51:90]
  wire [2:0] _GEN_63 = {{2'd0}, io_vcalloc_req_ready}; // @[InputUnit.scala 266:47]
  wire [2:0] _io_debug_va_stall_T_7 = _io_debug_va_stall_T_4 - _GEN_63; // @[InputUnit.scala 266:47]
  wire  _T_39 = io_vcalloc_req_ready & io_vcalloc_req_valid; // @[Decoupled.scala 51:35]
  wire [8:0] _credit_available_T = {states_0_vc_sel_2_0,1'h0,1'h0,1'h0,states_0_vc_sel_1_0,2'h0,1'h0,states_0_vc_sel_0_0
    }; // @[InputUnit.scala 287:40]
  wire [8:0] _credit_available_T_1 = {io_out_credit_available_2_0,io_out_credit_available_1_3,
    io_out_credit_available_1_2,io_out_credit_available_1_1,io_out_credit_available_1_0,io_out_credit_available_0_3,
    io_out_credit_available_0_2,io_out_credit_available_0_1,io_out_credit_available_0_0}; // @[InputUnit.scala 287:73]
  wire [8:0] _credit_available_T_2 = _credit_available_T & _credit_available_T_1; // @[InputUnit.scala 287:47]
  wire  credit_available = _credit_available_T_2 != 9'h0; // @[InputUnit.scala 287:81]
  wire  _T_60 = salloc_arb_io_in_0_ready & salloc_arb_io_in_0_valid; // @[Decoupled.scala 51:35]
  wire [8:0] _credit_available_T_3 = {states_1_vc_sel_2_0,1'h0,1'h0,states_1_vc_sel_1_1,1'h0,2'h0,states_1_vc_sel_0_1,
    states_1_vc_sel_0_0}; // @[InputUnit.scala 287:40]
  wire [8:0] _credit_available_T_5 = _credit_available_T_3 & _credit_available_T_1; // @[InputUnit.scala 287:47]
  wire  credit_available_1 = _credit_available_T_5 != 9'h0; // @[InputUnit.scala 287:81]
  wire  _T_62 = salloc_arb_io_in_1_ready & salloc_arb_io_in_1_valid; // @[Decoupled.scala 51:35]
  wire [8:0] _credit_available_T_6 = {states_2_vc_sel_2_0,1'h0,states_2_vc_sel_1_2,states_2_vc_sel_1_1,1'h0,1'h0,
    states_2_vc_sel_0_2,states_2_vc_sel_0_1,states_2_vc_sel_0_0}; // @[InputUnit.scala 287:40]
  wire [8:0] _credit_available_T_8 = _credit_available_T_6 & _credit_available_T_1; // @[InputUnit.scala 287:47]
  wire  credit_available_2 = _credit_available_T_8 != 9'h0; // @[InputUnit.scala 287:81]
  wire  _T_64 = salloc_arb_io_in_2_ready & salloc_arb_io_in_2_valid; // @[Decoupled.scala 51:35]
  wire [8:0] _credit_available_T_9 = {states_3_vc_sel_2_0,states_3_vc_sel_1_3,states_3_vc_sel_1_2,states_3_vc_sel_1_1,1'h0
    ,states_3_vc_sel_0_3,states_3_vc_sel_0_2,states_3_vc_sel_0_1,states_3_vc_sel_0_0}; // @[InputUnit.scala 287:40]
  wire [8:0] _credit_available_T_11 = _credit_available_T_9 & _credit_available_T_1; // @[InputUnit.scala 287:47]
  wire  credit_available_3 = _credit_available_T_11 != 9'h0; // @[InputUnit.scala 287:81]
  wire  _T_66 = salloc_arb_io_in_3_ready & salloc_arb_io_in_3_valid; // @[Decoupled.scala 51:35]
  wire  _io_debug_sa_stall_T_1 = salloc_arb_io_in_0_valid & ~salloc_arb_io_in_0_ready; // @[InputUnit.scala 301:67]
  wire  _io_debug_sa_stall_T_3 = salloc_arb_io_in_1_valid & ~salloc_arb_io_in_1_ready; // @[InputUnit.scala 301:67]
  wire  _io_debug_sa_stall_T_5 = salloc_arb_io_in_2_valid & ~salloc_arb_io_in_2_ready; // @[InputUnit.scala 301:67]
  wire  _io_debug_sa_stall_T_7 = salloc_arb_io_in_3_valid & ~salloc_arb_io_in_3_ready; // @[InputUnit.scala 301:67]
  wire [1:0] _io_debug_sa_stall_T_8 = _io_debug_sa_stall_T_1 + _io_debug_sa_stall_T_3; // @[Bitwise.scala 51:90]
  wire [1:0] _io_debug_sa_stall_T_10 = _io_debug_sa_stall_T_5 + _io_debug_sa_stall_T_7; // @[Bitwise.scala 51:90]
  wire [2:0] _io_debug_sa_stall_T_12 = _io_debug_sa_stall_T_8 + _io_debug_sa_stall_T_10; // @[Bitwise.scala 51:90]
  reg  salloc_outs_0_valid; // @[InputUnit.scala 318:8]
  reg [1:0] salloc_outs_0_out_vid; // @[InputUnit.scala 318:8]
  reg  salloc_outs_0_flit_head; // @[InputUnit.scala 318:8]
  reg  salloc_outs_0_flit_tail; // @[InputUnit.scala 318:8]
  reg [63:0] salloc_outs_0_flit_payload; // @[InputUnit.scala 318:8]
  reg [1:0] salloc_outs_0_flit_flow_ingress_node; // @[InputUnit.scala 318:8]
  reg [1:0] salloc_outs_0_flit_flow_egress_node; // @[InputUnit.scala 318:8]
  wire  _io_in_credit_return_T = salloc_arb_io_out_0_ready & salloc_arb_io_out_0_valid; // @[Decoupled.scala 51:35]
  wire  _io_in_vc_free_T_11 = salloc_arb_io_chosen_oh_0[0] & input_buffer_io_deq_0_bits_tail | salloc_arb_io_chosen_oh_0
    [1] & input_buffer_io_deq_1_bits_tail | salloc_arb_io_chosen_oh_0[2] & input_buffer_io_deq_2_bits_tail |
    salloc_arb_io_chosen_oh_0[3] & input_buffer_io_deq_3_bits_tail; // @[Mux.scala 27:73]
  wire  vc_sel_0_0 = salloc_arb_io_chosen_oh_0[0] & states_0_vc_sel_0_0 | salloc_arb_io_chosen_oh_0[1] &
    states_1_vc_sel_0_0 | salloc_arb_io_chosen_oh_0[2] & states_2_vc_sel_0_0 | salloc_arb_io_chosen_oh_0[3] &
    states_3_vc_sel_0_0; // @[Mux.scala 27:73]
  wire  vc_sel_0_1 = salloc_arb_io_chosen_oh_0[1] & states_1_vc_sel_0_1 | salloc_arb_io_chosen_oh_0[2] &
    states_2_vc_sel_0_1 | salloc_arb_io_chosen_oh_0[3] & states_3_vc_sel_0_1; // @[Mux.scala 27:73]
  wire  vc_sel_0_2 = salloc_arb_io_chosen_oh_0[2] & states_2_vc_sel_0_2 | salloc_arb_io_chosen_oh_0[3] &
    states_3_vc_sel_0_2; // @[Mux.scala 27:73]
  wire  vc_sel_0_3 = salloc_arb_io_chosen_oh_0[3] & states_3_vc_sel_0_3; // @[Mux.scala 27:73]
  wire  vc_sel_1_0 = salloc_arb_io_chosen_oh_0[0] & states_0_vc_sel_1_0; // @[Mux.scala 27:73]
  wire  vc_sel_1_1 = salloc_arb_io_chosen_oh_0[1] & states_1_vc_sel_1_1 | salloc_arb_io_chosen_oh_0[2] &
    states_2_vc_sel_1_1 | salloc_arb_io_chosen_oh_0[3] & states_3_vc_sel_1_1; // @[Mux.scala 27:73]
  wire  vc_sel_1_2 = salloc_arb_io_chosen_oh_0[2] & states_2_vc_sel_1_2 | salloc_arb_io_chosen_oh_0[3] &
    states_3_vc_sel_1_2; // @[Mux.scala 27:73]
  wire  vc_sel_1_3 = salloc_arb_io_chosen_oh_0[3] & states_3_vc_sel_1_3; // @[Mux.scala 27:73]
  wire  channel_oh_0 = vc_sel_0_0 | vc_sel_0_1 | vc_sel_0_2 | vc_sel_0_3; // @[InputUnit.scala 334:43]
  wire  channel_oh_1 = vc_sel_1_0 | vc_sel_1_1 | vc_sel_1_2 | vc_sel_1_3; // @[InputUnit.scala 334:43]
  wire [3:0] _virt_channel_T = {vc_sel_0_3,vc_sel_0_2,vc_sel_0_1,vc_sel_0_0}; // @[OneHot.scala 22:45]
  wire [1:0] virt_channel_hi_1 = _virt_channel_T[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] virt_channel_lo_1 = _virt_channel_T[1:0]; // @[OneHot.scala 31:18]
  wire  _virt_channel_T_1 = |virt_channel_hi_1; // @[OneHot.scala 32:14]
  wire [1:0] _virt_channel_T_2 = virt_channel_hi_1 | virt_channel_lo_1; // @[OneHot.scala 32:28]
  wire [1:0] _virt_channel_T_4 = {_virt_channel_T_1,_virt_channel_T_2[1]}; // @[Cat.scala 33:92]
  wire [3:0] _virt_channel_T_5 = {vc_sel_1_3,vc_sel_1_2,vc_sel_1_1,vc_sel_1_0}; // @[OneHot.scala 22:45]
  wire [1:0] virt_channel_hi_3 = _virt_channel_T_5[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] virt_channel_lo_3 = _virt_channel_T_5[1:0]; // @[OneHot.scala 31:18]
  wire  _virt_channel_T_6 = |virt_channel_hi_3; // @[OneHot.scala 32:14]
  wire [1:0] _virt_channel_T_7 = virt_channel_hi_3 | virt_channel_lo_3; // @[OneHot.scala 32:28]
  wire [1:0] _virt_channel_T_9 = {_virt_channel_T_6,_virt_channel_T_7[1]}; // @[Cat.scala 33:92]
  wire [1:0] _virt_channel_T_10 = channel_oh_0 ? _virt_channel_T_4 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _virt_channel_T_11 = channel_oh_1 ? _virt_channel_T_9 : 2'h0; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_4 = salloc_arb_io_chosen_oh_0[0] ? input_buffer_io_deq_0_bits_payload : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_5 = salloc_arb_io_chosen_oh_0[1] ? input_buffer_io_deq_1_bits_payload : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_6 = salloc_arb_io_chosen_oh_0[2] ? input_buffer_io_deq_2_bits_payload : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_7 = salloc_arb_io_chosen_oh_0[3] ? input_buffer_io_deq_3_bits_payload : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_8 = _salloc_outs_0_flit_payload_T_4 | _salloc_outs_0_flit_payload_T_5; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_9 = _salloc_outs_0_flit_payload_T_8 | _salloc_outs_0_flit_payload_T_6; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_11 = salloc_arb_io_chosen_oh_0[0] ? states_0_flow_egress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_12 = salloc_arb_io_chosen_oh_0[1] ? states_1_flow_egress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_13 = salloc_arb_io_chosen_oh_0[2] ? states_2_flow_egress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_14 = salloc_arb_io_chosen_oh_0[3] ? states_3_flow_egress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_15 = _salloc_outs_0_flit_flow_T_11 | _salloc_outs_0_flit_flow_T_12; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_16 = _salloc_outs_0_flit_flow_T_15 | _salloc_outs_0_flit_flow_T_13; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_25 = salloc_arb_io_chosen_oh_0[0] ? states_0_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_26 = salloc_arb_io_chosen_oh_0[1] ? states_1_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_27 = salloc_arb_io_chosen_oh_0[2] ? states_2_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_28 = salloc_arb_io_chosen_oh_0[3] ? states_3_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_29 = _salloc_outs_0_flit_flow_T_25 | _salloc_outs_0_flit_flow_T_26; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_30 = _salloc_outs_0_flit_flow_T_29 | _salloc_outs_0_flit_flow_T_27; // @[Mux.scala 27:73]
  InputBuffer input_buffer ( // @[InputUnit.scala 180:28]
    .clock(input_buffer_clock),
    .reset(input_buffer_reset),
    .io_enq_0_valid(input_buffer_io_enq_0_valid),
    .io_enq_0_bits_head(input_buffer_io_enq_0_bits_head),
    .io_enq_0_bits_tail(input_buffer_io_enq_0_bits_tail),
    .io_enq_0_bits_payload(input_buffer_io_enq_0_bits_payload),
    .io_enq_0_bits_virt_channel_id(input_buffer_io_enq_0_bits_virt_channel_id),
    .io_deq_0_ready(input_buffer_io_deq_0_ready),
    .io_deq_0_valid(input_buffer_io_deq_0_valid),
    .io_deq_0_bits_head(input_buffer_io_deq_0_bits_head),
    .io_deq_0_bits_tail(input_buffer_io_deq_0_bits_tail),
    .io_deq_0_bits_payload(input_buffer_io_deq_0_bits_payload),
    .io_deq_1_ready(input_buffer_io_deq_1_ready),
    .io_deq_1_valid(input_buffer_io_deq_1_valid),
    .io_deq_1_bits_head(input_buffer_io_deq_1_bits_head),
    .io_deq_1_bits_tail(input_buffer_io_deq_1_bits_tail),
    .io_deq_1_bits_payload(input_buffer_io_deq_1_bits_payload),
    .io_deq_2_ready(input_buffer_io_deq_2_ready),
    .io_deq_2_valid(input_buffer_io_deq_2_valid),
    .io_deq_2_bits_head(input_buffer_io_deq_2_bits_head),
    .io_deq_2_bits_tail(input_buffer_io_deq_2_bits_tail),
    .io_deq_2_bits_payload(input_buffer_io_deq_2_bits_payload),
    .io_deq_3_ready(input_buffer_io_deq_3_ready),
    .io_deq_3_valid(input_buffer_io_deq_3_valid),
    .io_deq_3_bits_head(input_buffer_io_deq_3_bits_head),
    .io_deq_3_bits_tail(input_buffer_io_deq_3_bits_tail),
    .io_deq_3_bits_payload(input_buffer_io_deq_3_bits_payload)
  );
  Arbiter route_arbiter ( // @[InputUnit.scala 186:29]
    .io_in_0_valid(route_arbiter_io_in_0_valid),
    .io_in_0_bits_flow_ingress_node(route_arbiter_io_in_0_bits_flow_ingress_node),
    .io_in_0_bits_flow_egress_node(route_arbiter_io_in_0_bits_flow_egress_node),
    .io_in_1_ready(route_arbiter_io_in_1_ready),
    .io_in_1_valid(route_arbiter_io_in_1_valid),
    .io_in_1_bits_flow_ingress_node(route_arbiter_io_in_1_bits_flow_ingress_node),
    .io_in_1_bits_flow_egress_node(route_arbiter_io_in_1_bits_flow_egress_node),
    .io_in_2_ready(route_arbiter_io_in_2_ready),
    .io_in_2_valid(route_arbiter_io_in_2_valid),
    .io_in_2_bits_flow_ingress_node(route_arbiter_io_in_2_bits_flow_ingress_node),
    .io_in_2_bits_flow_egress_node(route_arbiter_io_in_2_bits_flow_egress_node),
    .io_in_3_ready(route_arbiter_io_in_3_ready),
    .io_in_3_valid(route_arbiter_io_in_3_valid),
    .io_in_3_bits_flow_ingress_node(route_arbiter_io_in_3_bits_flow_ingress_node),
    .io_in_3_bits_flow_egress_node(route_arbiter_io_in_3_bits_flow_egress_node),
    .io_out_valid(route_arbiter_io_out_valid),
    .io_out_bits_src_virt_id(route_arbiter_io_out_bits_src_virt_id),
    .io_out_bits_flow_ingress_node(route_arbiter_io_out_bits_flow_ingress_node),
    .io_out_bits_flow_egress_node(route_arbiter_io_out_bits_flow_egress_node)
  );
  SwitchArbiter salloc_arb ( // @[InputUnit.scala 279:26]
    .clock(salloc_arb_clock),
    .reset(salloc_arb_reset),
    .io_in_0_ready(salloc_arb_io_in_0_ready),
    .io_in_0_valid(salloc_arb_io_in_0_valid),
    .io_in_0_bits_vc_sel_2_0(salloc_arb_io_in_0_bits_vc_sel_2_0),
    .io_in_0_bits_vc_sel_1_0(salloc_arb_io_in_0_bits_vc_sel_1_0),
    .io_in_0_bits_vc_sel_0_0(salloc_arb_io_in_0_bits_vc_sel_0_0),
    .io_in_0_bits_tail(salloc_arb_io_in_0_bits_tail),
    .io_in_1_ready(salloc_arb_io_in_1_ready),
    .io_in_1_valid(salloc_arb_io_in_1_valid),
    .io_in_1_bits_vc_sel_2_0(salloc_arb_io_in_1_bits_vc_sel_2_0),
    .io_in_1_bits_vc_sel_1_0(salloc_arb_io_in_1_bits_vc_sel_1_0),
    .io_in_1_bits_vc_sel_1_1(salloc_arb_io_in_1_bits_vc_sel_1_1),
    .io_in_1_bits_vc_sel_0_0(salloc_arb_io_in_1_bits_vc_sel_0_0),
    .io_in_1_bits_vc_sel_0_1(salloc_arb_io_in_1_bits_vc_sel_0_1),
    .io_in_1_bits_tail(salloc_arb_io_in_1_bits_tail),
    .io_in_2_ready(salloc_arb_io_in_2_ready),
    .io_in_2_valid(salloc_arb_io_in_2_valid),
    .io_in_2_bits_vc_sel_2_0(salloc_arb_io_in_2_bits_vc_sel_2_0),
    .io_in_2_bits_vc_sel_1_0(salloc_arb_io_in_2_bits_vc_sel_1_0),
    .io_in_2_bits_vc_sel_1_1(salloc_arb_io_in_2_bits_vc_sel_1_1),
    .io_in_2_bits_vc_sel_1_2(salloc_arb_io_in_2_bits_vc_sel_1_2),
    .io_in_2_bits_vc_sel_0_0(salloc_arb_io_in_2_bits_vc_sel_0_0),
    .io_in_2_bits_vc_sel_0_1(salloc_arb_io_in_2_bits_vc_sel_0_1),
    .io_in_2_bits_vc_sel_0_2(salloc_arb_io_in_2_bits_vc_sel_0_2),
    .io_in_2_bits_tail(salloc_arb_io_in_2_bits_tail),
    .io_in_3_ready(salloc_arb_io_in_3_ready),
    .io_in_3_valid(salloc_arb_io_in_3_valid),
    .io_in_3_bits_vc_sel_2_0(salloc_arb_io_in_3_bits_vc_sel_2_0),
    .io_in_3_bits_vc_sel_1_0(salloc_arb_io_in_3_bits_vc_sel_1_0),
    .io_in_3_bits_vc_sel_1_1(salloc_arb_io_in_3_bits_vc_sel_1_1),
    .io_in_3_bits_vc_sel_1_2(salloc_arb_io_in_3_bits_vc_sel_1_2),
    .io_in_3_bits_vc_sel_1_3(salloc_arb_io_in_3_bits_vc_sel_1_3),
    .io_in_3_bits_vc_sel_0_0(salloc_arb_io_in_3_bits_vc_sel_0_0),
    .io_in_3_bits_vc_sel_0_1(salloc_arb_io_in_3_bits_vc_sel_0_1),
    .io_in_3_bits_vc_sel_0_2(salloc_arb_io_in_3_bits_vc_sel_0_2),
    .io_in_3_bits_vc_sel_0_3(salloc_arb_io_in_3_bits_vc_sel_0_3),
    .io_in_3_bits_tail(salloc_arb_io_in_3_bits_tail),
    .io_out_0_ready(salloc_arb_io_out_0_ready),
    .io_out_0_valid(salloc_arb_io_out_0_valid),
    .io_out_0_bits_vc_sel_2_0(salloc_arb_io_out_0_bits_vc_sel_2_0),
    .io_out_0_bits_vc_sel_1_0(salloc_arb_io_out_0_bits_vc_sel_1_0),
    .io_out_0_bits_vc_sel_1_1(salloc_arb_io_out_0_bits_vc_sel_1_1),
    .io_out_0_bits_vc_sel_1_2(salloc_arb_io_out_0_bits_vc_sel_1_2),
    .io_out_0_bits_vc_sel_1_3(salloc_arb_io_out_0_bits_vc_sel_1_3),
    .io_out_0_bits_vc_sel_0_0(salloc_arb_io_out_0_bits_vc_sel_0_0),
    .io_out_0_bits_vc_sel_0_1(salloc_arb_io_out_0_bits_vc_sel_0_1),
    .io_out_0_bits_vc_sel_0_2(salloc_arb_io_out_0_bits_vc_sel_0_2),
    .io_out_0_bits_vc_sel_0_3(salloc_arb_io_out_0_bits_vc_sel_0_3),
    .io_out_0_bits_tail(salloc_arb_io_out_0_bits_tail),
    .io_chosen_oh_0(salloc_arb_io_chosen_oh_0)
  );
  assign io_router_req_valid = route_arbiter_io_out_valid; // @[InputUnit.scala 189:17]
  assign io_router_req_bits_src_virt_id = route_arbiter_io_out_bits_src_virt_id; // @[InputUnit.scala 189:17]
  assign io_router_req_bits_flow_ingress_node = route_arbiter_io_out_bits_flow_ingress_node; // @[InputUnit.scala 189:17]
  assign io_router_req_bits_flow_egress_node = route_arbiter_io_out_bits_flow_egress_node; // @[InputUnit.scala 189:17]
  assign io_vcalloc_req_valid = vcalloc_vals_0 | vcalloc_vals_1 | vcalloc_vals_2 | vcalloc_vals_3; // @[package.scala 73:59]
  assign io_vcalloc_req_bits_vc_sel_2_0 = vcalloc_sel[0] & states_0_vc_sel_2_0 | vcalloc_sel[1] & states_1_vc_sel_2_0 |
    vcalloc_sel[2] & states_2_vc_sel_2_0 | vcalloc_sel[3] & states_3_vc_sel_2_0; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_1_0 = vcalloc_sel[0] & states_0_vc_sel_1_0; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_1_1 = vcalloc_sel[1] & states_1_vc_sel_1_1 | vcalloc_sel[2] & states_2_vc_sel_1_1 |
    vcalloc_sel[3] & states_3_vc_sel_1_1; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_1_2 = vcalloc_sel[2] & states_2_vc_sel_1_2 | vcalloc_sel[3] & states_3_vc_sel_1_2; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_1_3 = vcalloc_sel[3] & states_3_vc_sel_1_3; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_0_0 = vcalloc_sel[0] & states_0_vc_sel_0_0 | vcalloc_sel[1] & states_1_vc_sel_0_0 |
    vcalloc_sel[2] & states_2_vc_sel_0_0 | vcalloc_sel[3] & states_3_vc_sel_0_0; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_0_1 = vcalloc_sel[1] & states_1_vc_sel_0_1 | vcalloc_sel[2] & states_2_vc_sel_0_1 |
    vcalloc_sel[3] & states_3_vc_sel_0_1; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_0_2 = vcalloc_sel[2] & states_2_vc_sel_0_2 | vcalloc_sel[3] & states_3_vc_sel_0_2; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_0_3 = vcalloc_sel[3] & states_3_vc_sel_0_3; // @[Mux.scala 27:73]
  assign io_salloc_req_0_valid = salloc_arb_io_out_0_valid; // @[InputUnit.scala 302:17 303:19 305:35]
  assign io_salloc_req_0_bits_vc_sel_2_0 = salloc_arb_io_out_0_bits_vc_sel_2_0; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_1_0 = salloc_arb_io_out_0_bits_vc_sel_1_0; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_1_1 = salloc_arb_io_out_0_bits_vc_sel_1_1; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_1_2 = salloc_arb_io_out_0_bits_vc_sel_1_2; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_1_3 = salloc_arb_io_out_0_bits_vc_sel_1_3; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_0_0 = salloc_arb_io_out_0_bits_vc_sel_0_0; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_0_1 = salloc_arb_io_out_0_bits_vc_sel_0_1; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_0_2 = salloc_arb_io_out_0_bits_vc_sel_0_2; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_0_3 = salloc_arb_io_out_0_bits_vc_sel_0_3; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_tail = salloc_arb_io_out_0_bits_tail; // @[InputUnit.scala 302:17]
  assign io_out_0_valid = salloc_outs_0_valid; // @[InputUnit.scala 349:21]
  assign io_out_0_bits_flit_head = salloc_outs_0_flit_head; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_flit_tail = salloc_outs_0_flit_tail; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_flit_payload = salloc_outs_0_flit_payload; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_flit_flow_ingress_node = salloc_outs_0_flit_flow_ingress_node; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_flit_flow_egress_node = salloc_outs_0_flit_flow_egress_node; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_out_virt_channel = salloc_outs_0_out_vid; // @[InputUnit.scala 351:37]
  assign io_debug_va_stall = _io_debug_va_stall_T_7[1:0]; // @[InputUnit.scala 266:21]
  assign io_debug_sa_stall = _io_debug_sa_stall_T_12[1:0]; // @[InputUnit.scala 301:21]
  assign io_in_credit_return = _io_in_credit_return_T ? salloc_arb_io_chosen_oh_0 : 4'h0; // @[InputUnit.scala 322:8]
  assign io_in_vc_free = _io_in_credit_return_T & _io_in_vc_free_T_11 ? salloc_arb_io_chosen_oh_0 : 4'h0; // @[InputUnit.scala 325:8]
  assign input_buffer_clock = clock;
  assign input_buffer_reset = reset;
  assign input_buffer_io_enq_0_valid = io_in_flit_0_valid; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_head = io_in_flit_0_bits_head; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_tail = io_in_flit_0_bits_tail; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_payload = io_in_flit_0_bits_payload; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_virt_channel_id = io_in_flit_0_bits_virt_channel_id; // @[InputUnit.scala 182:28]
  assign input_buffer_io_deq_0_ready = salloc_arb_io_in_0_ready; // @[InputUnit.scala 295:36]
  assign input_buffer_io_deq_1_ready = salloc_arb_io_in_1_ready; // @[InputUnit.scala 295:36]
  assign input_buffer_io_deq_2_ready = salloc_arb_io_in_2_ready; // @[InputUnit.scala 295:36]
  assign input_buffer_io_deq_3_ready = salloc_arb_io_in_3_ready; // @[InputUnit.scala 295:36]
  assign route_arbiter_io_in_0_valid = states_0_g == 3'h1; // @[InputUnit.scala 212:22]
  assign route_arbiter_io_in_0_bits_flow_ingress_node = states_0_flow_ingress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_0_bits_flow_egress_node = states_0_flow_egress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_1_valid = states_1_g == 3'h1; // @[InputUnit.scala 212:22]
  assign route_arbiter_io_in_1_bits_flow_ingress_node = states_1_flow_ingress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_1_bits_flow_egress_node = states_1_flow_egress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_2_valid = states_2_g == 3'h1; // @[InputUnit.scala 212:22]
  assign route_arbiter_io_in_2_bits_flow_ingress_node = states_2_flow_ingress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_2_bits_flow_egress_node = states_2_flow_egress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_3_valid = states_3_g == 3'h1; // @[InputUnit.scala 212:22]
  assign route_arbiter_io_in_3_bits_flow_ingress_node = states_3_flow_ingress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_3_bits_flow_egress_node = states_3_flow_egress_node; // @[InputUnit.scala 213:19]
  assign salloc_arb_clock = clock;
  assign salloc_arb_reset = reset;
  assign salloc_arb_io_in_0_valid = states_0_g == 3'h3 & credit_available & input_buffer_io_deq_0_valid; // @[InputUnit.scala 288:50]
  assign salloc_arb_io_in_0_bits_vc_sel_2_0 = states_0_vc_sel_2_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_0_bits_vc_sel_1_0 = states_0_vc_sel_1_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_0_bits_vc_sel_0_0 = states_0_vc_sel_0_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_0_bits_tail = input_buffer_io_deq_0_bits_tail; // @[InputUnit.scala 291:19]
  assign salloc_arb_io_in_1_valid = states_1_g == 3'h3 & credit_available_1 & input_buffer_io_deq_1_valid; // @[InputUnit.scala 288:50]
  assign salloc_arb_io_in_1_bits_vc_sel_2_0 = states_1_vc_sel_2_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_1_bits_vc_sel_1_0 = 1'h0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_1_bits_vc_sel_1_1 = states_1_vc_sel_1_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_1_bits_vc_sel_0_0 = states_1_vc_sel_0_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_1_bits_vc_sel_0_1 = states_1_vc_sel_0_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_1_bits_tail = input_buffer_io_deq_1_bits_tail; // @[InputUnit.scala 291:19]
  assign salloc_arb_io_in_2_valid = states_2_g == 3'h3 & credit_available_2 & input_buffer_io_deq_2_valid; // @[InputUnit.scala 288:50]
  assign salloc_arb_io_in_2_bits_vc_sel_2_0 = states_2_vc_sel_2_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_1_0 = 1'h0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_1_1 = states_2_vc_sel_1_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_1_2 = states_2_vc_sel_1_2; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_0_0 = states_2_vc_sel_0_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_0_1 = states_2_vc_sel_0_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_0_2 = states_2_vc_sel_0_2; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_tail = input_buffer_io_deq_2_bits_tail; // @[InputUnit.scala 291:19]
  assign salloc_arb_io_in_3_valid = states_3_g == 3'h3 & credit_available_3 & input_buffer_io_deq_3_valid; // @[InputUnit.scala 288:50]
  assign salloc_arb_io_in_3_bits_vc_sel_2_0 = states_3_vc_sel_2_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_1_0 = 1'h0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_1_1 = states_3_vc_sel_1_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_1_2 = states_3_vc_sel_1_2; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_1_3 = states_3_vc_sel_1_3; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_0_0 = states_3_vc_sel_0_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_0_1 = states_3_vc_sel_0_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_0_2 = states_3_vc_sel_0_2; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_0_3 = states_3_vc_sel_0_3; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_tail = input_buffer_io_deq_3_bits_tail; // @[InputUnit.scala 291:19]
  assign salloc_arb_io_out_0_ready = io_salloc_req_0_ready; // @[InputUnit.scala 302:17 303:19 304:39]
  always @(posedge clock) begin
    if (reset) begin // @[InputUnit.scala 377:23]
      states_0_g <= 3'h0; // @[InputUnit.scala 378:24]
    end else if (_T_60 & input_buffer_io_deq_0_bits_tail) begin // @[InputUnit.scala 292:35]
      states_0_g <= 3'h0; // @[InputUnit.scala 293:13]
    end else if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[0]) begin // @[InputUnit.scala 270:29]
        states_0_g <= 3'h3; // @[InputUnit.scala 272:21]
      end else begin
        states_0_g <= _GEN_222;
      end
    end else begin
      states_0_g <= _GEN_222;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[0]) begin // @[InputUnit.scala 270:29]
        states_0_vc_sel_2_0 <= io_vcalloc_resp_vc_sel_2_0; // @[InputUnit.scala 271:26]
      end else begin
        states_0_vc_sel_2_0 <= _GEN_184;
      end
    end else begin
      states_0_vc_sel_2_0 <= _GEN_184;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[0]) begin // @[InputUnit.scala 270:29]
        states_0_vc_sel_1_0 <= io_vcalloc_resp_vc_sel_1_0; // @[InputUnit.scala 271:26]
      end else begin
        states_0_vc_sel_1_0 <= _GEN_185;
      end
    end else begin
      states_0_vc_sel_1_0 <= _GEN_185;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[0]) begin // @[InputUnit.scala 270:29]
        states_0_vc_sel_0_0 <= io_vcalloc_resp_vc_sel_0_0; // @[InputUnit.scala 271:26]
      end else begin
        states_0_vc_sel_0_0 <= _GEN_189;
      end
    end else begin
      states_0_vc_sel_0_0 <= _GEN_189;
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h0 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_0_flow_ingress_node <= io_in_flit_0_bits_flow_ingress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h0 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_0_flow_egress_node <= io_in_flit_0_bits_flow_egress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (reset) begin // @[InputUnit.scala 377:23]
      states_1_g <= 3'h0; // @[InputUnit.scala 378:24]
    end else if (_T_62 & input_buffer_io_deq_1_bits_tail) begin // @[InputUnit.scala 292:35]
      states_1_g <= 3'h0; // @[InputUnit.scala 293:13]
    end else if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_g <= 3'h3; // @[InputUnit.scala 272:21]
      end else begin
        states_1_g <= _GEN_223;
      end
    end else begin
      states_1_g <= _GEN_223;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_vc_sel_2_0 <= io_vcalloc_resp_vc_sel_2_0; // @[InputUnit.scala 271:26]
      end else begin
        states_1_vc_sel_2_0 <= _GEN_193;
      end
    end else begin
      states_1_vc_sel_2_0 <= _GEN_193;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_vc_sel_1_1 <= io_vcalloc_resp_vc_sel_1_1; // @[InputUnit.scala 271:26]
      end else begin
        states_1_vc_sel_1_1 <= _GEN_195;
      end
    end else begin
      states_1_vc_sel_1_1 <= _GEN_195;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_vc_sel_0_0 <= io_vcalloc_resp_vc_sel_0_0; // @[InputUnit.scala 271:26]
      end else begin
        states_1_vc_sel_0_0 <= _GEN_198;
      end
    end else begin
      states_1_vc_sel_0_0 <= _GEN_198;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_vc_sel_0_1 <= io_vcalloc_resp_vc_sel_0_1; // @[InputUnit.scala 271:26]
      end else begin
        states_1_vc_sel_0_1 <= _GEN_199;
      end
    end else begin
      states_1_vc_sel_0_1 <= _GEN_199;
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h1 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_1_flow_ingress_node <= io_in_flit_0_bits_flow_ingress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h1 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_1_flow_egress_node <= io_in_flit_0_bits_flow_egress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (reset) begin // @[InputUnit.scala 377:23]
      states_2_g <= 3'h0; // @[InputUnit.scala 378:24]
    end else if (_T_64 & input_buffer_io_deq_2_bits_tail) begin // @[InputUnit.scala 292:35]
      states_2_g <= 3'h0; // @[InputUnit.scala 293:13]
    end else if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_g <= 3'h3; // @[InputUnit.scala 272:21]
      end else begin
        states_2_g <= _GEN_224;
      end
    end else begin
      states_2_g <= _GEN_224;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_2_0 <= io_vcalloc_resp_vc_sel_2_0; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_2_0 <= _GEN_202;
      end
    end else begin
      states_2_vc_sel_2_0 <= _GEN_202;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_1_1 <= io_vcalloc_resp_vc_sel_1_1; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_1_1 <= _GEN_204;
      end
    end else begin
      states_2_vc_sel_1_1 <= _GEN_204;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_1_2 <= io_vcalloc_resp_vc_sel_1_2; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_1_2 <= _GEN_205;
      end
    end else begin
      states_2_vc_sel_1_2 <= _GEN_205;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_0_0 <= io_vcalloc_resp_vc_sel_0_0; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_0_0 <= _GEN_207;
      end
    end else begin
      states_2_vc_sel_0_0 <= _GEN_207;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_0_1 <= io_vcalloc_resp_vc_sel_0_1; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_0_1 <= _GEN_208;
      end
    end else begin
      states_2_vc_sel_0_1 <= _GEN_208;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_0_2 <= io_vcalloc_resp_vc_sel_0_2; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_0_2 <= _GEN_209;
      end
    end else begin
      states_2_vc_sel_0_2 <= _GEN_209;
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h2 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_2_flow_ingress_node <= io_in_flit_0_bits_flow_ingress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h2 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_2_flow_egress_node <= io_in_flit_0_bits_flow_egress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (reset) begin // @[InputUnit.scala 377:23]
      states_3_g <= 3'h0; // @[InputUnit.scala 378:24]
    end else if (_T_66 & input_buffer_io_deq_3_bits_tail) begin // @[InputUnit.scala 292:35]
      states_3_g <= 3'h0; // @[InputUnit.scala 293:13]
    end else if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_g <= 3'h3; // @[InputUnit.scala 272:21]
      end else begin
        states_3_g <= _GEN_225;
      end
    end else begin
      states_3_g <= _GEN_225;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_2_0 <= io_vcalloc_resp_vc_sel_2_0; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_2_0 <= _GEN_211;
      end
    end else begin
      states_3_vc_sel_2_0 <= _GEN_211;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_1_1 <= io_vcalloc_resp_vc_sel_1_1; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_1_1 <= _GEN_213;
      end
    end else begin
      states_3_vc_sel_1_1 <= _GEN_213;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_1_2 <= io_vcalloc_resp_vc_sel_1_2; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_1_2 <= _GEN_214;
      end
    end else begin
      states_3_vc_sel_1_2 <= _GEN_214;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_1_3 <= io_vcalloc_resp_vc_sel_1_3; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_1_3 <= _GEN_215;
      end
    end else begin
      states_3_vc_sel_1_3 <= _GEN_215;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_0_0 <= io_vcalloc_resp_vc_sel_0_0; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_0_0 <= _GEN_216;
      end
    end else begin
      states_3_vc_sel_0_0 <= _GEN_216;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_0_1 <= io_vcalloc_resp_vc_sel_0_1; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_0_1 <= _GEN_217;
      end
    end else begin
      states_3_vc_sel_0_1 <= _GEN_217;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_0_2 <= io_vcalloc_resp_vc_sel_0_2; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_0_2 <= _GEN_218;
      end
    end else begin
      states_3_vc_sel_0_2 <= _GEN_218;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_0_3 <= io_vcalloc_resp_vc_sel_0_3; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_0_3 <= _GEN_219;
      end
    end else begin
      states_3_vc_sel_0_3 <= _GEN_219;
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h3 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_3_flow_ingress_node <= io_in_flit_0_bits_flow_ingress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h3 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_3_flow_egress_node <= io_in_flit_0_bits_flow_egress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (reset) begin // @[InputUnit.scala 233:21]
      mask <= 4'h0; // @[InputUnit.scala 233:21]
    end else if (io_router_req_valid) begin // @[InputUnit.scala 239:31]
      mask <= _mask_T_2; // @[InputUnit.scala 240:10]
    end else if (_T_26) begin // @[InputUnit.scala 241:34]
      mask <= _mask_T_17; // @[InputUnit.scala 242:10]
    end
    salloc_outs_0_valid <= salloc_arb_io_out_0_ready & salloc_arb_io_out_0_valid; // @[Decoupled.scala 51:35]
    salloc_outs_0_out_vid <= _virt_channel_T_10 | _virt_channel_T_11; // @[Mux.scala 27:73]
    salloc_outs_0_flit_head <= salloc_arb_io_chosen_oh_0[0] & input_buffer_io_deq_0_bits_head |
      salloc_arb_io_chosen_oh_0[1] & input_buffer_io_deq_1_bits_head | salloc_arb_io_chosen_oh_0[2] &
      input_buffer_io_deq_2_bits_head | salloc_arb_io_chosen_oh_0[3] & input_buffer_io_deq_3_bits_head; // @[Mux.scala 27:73]
    salloc_outs_0_flit_tail <= salloc_arb_io_chosen_oh_0[0] & input_buffer_io_deq_0_bits_tail |
      salloc_arb_io_chosen_oh_0[1] & input_buffer_io_deq_1_bits_tail | salloc_arb_io_chosen_oh_0[2] &
      input_buffer_io_deq_2_bits_tail | salloc_arb_io_chosen_oh_0[3] & input_buffer_io_deq_3_bits_tail; // @[Mux.scala 27:73]
    salloc_outs_0_flit_payload <= _salloc_outs_0_flit_payload_T_9 | _salloc_outs_0_flit_payload_T_7; // @[Mux.scala 27:73]
    salloc_outs_0_flit_flow_ingress_node <= _salloc_outs_0_flit_flow_T_30 | _salloc_outs_0_flit_flow_T_28; // @[Mux.scala 27:73]
    salloc_outs_0_flit_flow_egress_node <= _salloc_outs_0_flit_flow_T_16 | _salloc_outs_0_flit_flow_T_14; // @[Mux.scala 27:73]
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T & _T_3 & ~(_GEN_3 == 3'h0)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:197 assert(states(id).g === g_i)\n"); // @[InputUnit.scala 197:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_router_req_valid & _T_3 & ~(_GEN_139 == 3'h1)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:224 assert(states(id).g === g_r)\n"); // @[InputUnit.scala 224:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_39 & vcalloc_sel[0] & _T_3 & ~vcalloc_vals_0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:274 assert(states(i).g === g_v)\n"); // @[InputUnit.scala 274:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_39 & vcalloc_sel[1] & _T_3 & ~vcalloc_vals_1) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:274 assert(states(i).g === g_v)\n"); // @[InputUnit.scala 274:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_39 & vcalloc_sel[2] & _T_3 & ~vcalloc_vals_2) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:274 assert(states(i).g === g_v)\n"); // @[InputUnit.scala 274:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_39 & vcalloc_sel[3] & _T_3 & ~vcalloc_vals_3) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:274 assert(states(i).g === g_v)\n"); // @[InputUnit.scala 274:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  states_0_g = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  states_0_vc_sel_2_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  states_0_vc_sel_1_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  states_0_vc_sel_0_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  states_0_flow_ingress_node = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  states_0_flow_egress_node = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  states_1_g = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  states_1_vc_sel_2_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  states_1_vc_sel_1_1 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  states_1_vc_sel_0_0 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  states_1_vc_sel_0_1 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  states_1_flow_ingress_node = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  states_1_flow_egress_node = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  states_2_g = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  states_2_vc_sel_2_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  states_2_vc_sel_1_1 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  states_2_vc_sel_1_2 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  states_2_vc_sel_0_0 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  states_2_vc_sel_0_1 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  states_2_vc_sel_0_2 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  states_2_flow_ingress_node = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  states_2_flow_egress_node = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  states_3_g = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  states_3_vc_sel_2_0 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  states_3_vc_sel_1_1 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  states_3_vc_sel_1_2 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  states_3_vc_sel_1_3 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  states_3_vc_sel_0_0 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  states_3_vc_sel_0_1 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  states_3_vc_sel_0_2 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  states_3_vc_sel_0_3 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  states_3_flow_ingress_node = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  states_3_flow_egress_node = _RAND_32[1:0];
  _RAND_33 = {1{`RANDOM}};
  mask = _RAND_33[3:0];
  _RAND_34 = {1{`RANDOM}};
  salloc_outs_0_valid = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  salloc_outs_0_out_vid = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  salloc_outs_0_flit_head = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  salloc_outs_0_flit_tail = _RAND_37[0:0];
  _RAND_38 = {2{`RANDOM}};
  salloc_outs_0_flit_payload = _RAND_38[63:0];
  _RAND_39 = {1{`RANDOM}};
  salloc_outs_0_flit_flow_ingress_node = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  salloc_outs_0_flit_flow_egress_node = _RAND_40[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (_T & ~reset) begin
      assert(1'h1); // @[InputUnit.scala 196:13]
    end
    //
    if (_T & _T_3) begin
      assert(_GEN_3 == 3'h0); // @[InputUnit.scala 197:13]
    end
    //
    if (io_router_req_valid & _T_3) begin
      assert(_GEN_139 == 3'h1); // @[InputUnit.scala 224:11]
    end
    //
    if (_T_39 & vcalloc_sel[0] & _T_3) begin
      assert(vcalloc_vals_0); // @[InputUnit.scala 274:17]
    end
    //
    if (_T_39 & vcalloc_sel[1] & _T_3) begin
      assert(vcalloc_vals_1); // @[InputUnit.scala 274:17]
    end
    //
    if (_T_39 & vcalloc_sel[2] & _T_3) begin
      assert(vcalloc_vals_2); // @[InputUnit.scala 274:17]
    end
    //
    if (_T_39 & vcalloc_sel[3] & _T_3) begin
      assert(vcalloc_vals_3); // @[InputUnit.scala 274:17]
    end
  end
endmodule
module IngressUnit_2(
  input         clock,
  input         reset,
  output        io_router_req_valid,
  output [1:0]  io_router_req_bits_flow_ingress_node,
  output [1:0]  io_router_req_bits_flow_egress_node,
  input         io_router_resp_vc_sel_1_0,
  input         io_router_resp_vc_sel_1_1,
  input         io_router_resp_vc_sel_1_2,
  input         io_router_resp_vc_sel_1_3,
  input         io_router_resp_vc_sel_0_0,
  input         io_router_resp_vc_sel_0_1,
  input         io_router_resp_vc_sel_0_2,
  input         io_router_resp_vc_sel_0_3,
  input         io_vcalloc_req_ready,
  output        io_vcalloc_req_valid,
  output        io_vcalloc_req_bits_vc_sel_2_0,
  output        io_vcalloc_req_bits_vc_sel_1_0,
  output        io_vcalloc_req_bits_vc_sel_1_1,
  output        io_vcalloc_req_bits_vc_sel_1_2,
  output        io_vcalloc_req_bits_vc_sel_1_3,
  output        io_vcalloc_req_bits_vc_sel_0_0,
  output        io_vcalloc_req_bits_vc_sel_0_1,
  output        io_vcalloc_req_bits_vc_sel_0_2,
  output        io_vcalloc_req_bits_vc_sel_0_3,
  input         io_vcalloc_resp_vc_sel_2_0,
  input         io_vcalloc_resp_vc_sel_1_0,
  input         io_vcalloc_resp_vc_sel_1_1,
  input         io_vcalloc_resp_vc_sel_1_2,
  input         io_vcalloc_resp_vc_sel_1_3,
  input         io_vcalloc_resp_vc_sel_0_0,
  input         io_vcalloc_resp_vc_sel_0_1,
  input         io_vcalloc_resp_vc_sel_0_2,
  input         io_vcalloc_resp_vc_sel_0_3,
  input         io_out_credit_available_2_0,
  input         io_out_credit_available_1_0,
  input         io_out_credit_available_1_1,
  input         io_out_credit_available_1_2,
  input         io_out_credit_available_1_3,
  input         io_out_credit_available_0_0,
  input         io_out_credit_available_0_1,
  input         io_out_credit_available_0_2,
  input         io_out_credit_available_0_3,
  input         io_salloc_req_0_ready,
  output        io_salloc_req_0_valid,
  output        io_salloc_req_0_bits_vc_sel_2_0,
  output        io_salloc_req_0_bits_vc_sel_1_0,
  output        io_salloc_req_0_bits_vc_sel_1_1,
  output        io_salloc_req_0_bits_vc_sel_1_2,
  output        io_salloc_req_0_bits_vc_sel_1_3,
  output        io_salloc_req_0_bits_vc_sel_0_0,
  output        io_salloc_req_0_bits_vc_sel_0_1,
  output        io_salloc_req_0_bits_vc_sel_0_2,
  output        io_salloc_req_0_bits_vc_sel_0_3,
  output        io_salloc_req_0_bits_tail,
  output        io_out_0_valid,
  output        io_out_0_bits_flit_head,
  output        io_out_0_bits_flit_tail,
  output [63:0] io_out_0_bits_flit_payload,
  output [1:0]  io_out_0_bits_flit_flow_ingress_node,
  output [1:0]  io_out_0_bits_flit_flow_egress_node,
  output [1:0]  io_out_0_bits_out_virt_channel,
  output        io_in_ready,
  input         io_in_valid,
  input         io_in_bits_head,
  input         io_in_bits_tail,
  input  [63:0] io_in_bits_payload,
  input  [1:0]  io_in_bits_egress_id
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  route_buffer_clock; // @[IngressUnit.scala 26:28]
  wire  route_buffer_reset; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_enq_ready; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_enq_valid; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_enq_bits_head; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_enq_bits_tail; // @[IngressUnit.scala 26:28]
  wire [63:0] route_buffer_io_enq_bits_payload; // @[IngressUnit.scala 26:28]
  wire [1:0] route_buffer_io_enq_bits_flow_ingress_node; // @[IngressUnit.scala 26:28]
  wire [1:0] route_buffer_io_enq_bits_flow_egress_node; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_deq_ready; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_deq_valid; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_deq_bits_head; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_deq_bits_tail; // @[IngressUnit.scala 26:28]
  wire [63:0] route_buffer_io_deq_bits_payload; // @[IngressUnit.scala 26:28]
  wire [1:0] route_buffer_io_deq_bits_flow_ingress_node; // @[IngressUnit.scala 26:28]
  wire [1:0] route_buffer_io_deq_bits_flow_egress_node; // @[IngressUnit.scala 26:28]
  wire  route_q_clock; // @[IngressUnit.scala 27:23]
  wire  route_q_reset; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_ready; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_valid; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_2_0; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_1_0; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_1_1; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_1_2; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_1_3; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_0_0; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_0_1; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_0_2; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_0_3; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_ready; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_valid; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_2_0; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_1_0; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_1_1; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_1_2; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_1_3; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_0_0; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_0_1; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_0_2; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_0_3; // @[IngressUnit.scala 27:23]
  wire  vcalloc_buffer_clock; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_reset; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_enq_ready; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_enq_valid; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_enq_bits_head; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_enq_bits_tail; // @[IngressUnit.scala 75:30]
  wire [63:0] vcalloc_buffer_io_enq_bits_payload; // @[IngressUnit.scala 75:30]
  wire [1:0] vcalloc_buffer_io_enq_bits_flow_ingress_node; // @[IngressUnit.scala 75:30]
  wire [1:0] vcalloc_buffer_io_enq_bits_flow_egress_node; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_deq_ready; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_deq_valid; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_deq_bits_head; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_deq_bits_tail; // @[IngressUnit.scala 75:30]
  wire [63:0] vcalloc_buffer_io_deq_bits_payload; // @[IngressUnit.scala 75:30]
  wire [1:0] vcalloc_buffer_io_deq_bits_flow_ingress_node; // @[IngressUnit.scala 75:30]
  wire [1:0] vcalloc_buffer_io_deq_bits_flow_egress_node; // @[IngressUnit.scala 75:30]
  wire  vcalloc_q_clock; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_reset; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_ready; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_valid; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_2_0; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_1_0; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_1_1; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_1_2; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_1_3; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_0_0; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_0_1; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_0_2; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_0_3; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_ready; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_valid; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_2_0; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_1_0; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_1_1; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_1_2; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_1_3; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_0_0; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_0_1; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_0_2; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_0_3; // @[IngressUnit.scala 76:25]
  wire  _T = 2'h0 == io_in_bits_egress_id; // @[IngressUnit.scala 30:72]
  wire  _T_1 = 2'h1 == io_in_bits_egress_id; // @[IngressUnit.scala 30:72]
  wire  _T_2 = 2'h2 == io_in_bits_egress_id; // @[IngressUnit.scala 30:72]
  wire  _T_3 = 2'h3 == io_in_bits_egress_id; // @[IngressUnit.scala 30:72]
  wire  _T_6 = _T | _T_1 | _T_2 | _T_3; // @[package.scala 73:59]
  wire  _T_11 = ~reset; // @[IngressUnit.scala 30:9]
  wire [1:0] _route_buffer_io_enq_bits_flow_egress_node_T_6 = _T_2 ? 2'h2 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _route_buffer_io_enq_bits_flow_egress_node_T_7 = _T_3 ? 2'h3 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _GEN_11 = {{1'd0}, _T_1}; // @[Mux.scala 27:73]
  wire [1:0] _route_buffer_io_enq_bits_flow_egress_node_T_9 = _GEN_11 | _route_buffer_io_enq_bits_flow_egress_node_T_6; // @[Mux.scala 27:73]
  wire  at_dest = route_buffer_io_enq_bits_flow_egress_node == 2'h2; // @[IngressUnit.scala 55:59]
  wire  _T_13 = io_in_ready & io_in_valid; // @[Decoupled.scala 51:35]
  wire  _vcalloc_buffer_io_enq_valid_T = ~route_buffer_io_deq_bits_head; // @[IngressUnit.scala 88:30]
  wire  _vcalloc_buffer_io_enq_valid_T_1 = route_q_io_deq_valid | ~route_buffer_io_deq_bits_head; // @[IngressUnit.scala 88:27]
  wire  _vcalloc_buffer_io_enq_valid_T_2 = route_buffer_io_deq_valid & _vcalloc_buffer_io_enq_valid_T_1; // @[IngressUnit.scala 87:61]
  wire  _vcalloc_buffer_io_enq_valid_T_4 = io_vcalloc_req_ready | _vcalloc_buffer_io_enq_valid_T; // @[IngressUnit.scala 89:27]
  wire  _io_vcalloc_req_valid_T_1 = route_buffer_io_deq_valid & route_q_io_deq_valid & route_buffer_io_deq_bits_head; // @[IngressUnit.scala 91:78]
  wire  _route_buffer_io_deq_ready_T_2 = vcalloc_buffer_io_enq_ready & _vcalloc_buffer_io_enq_valid_T_1; // @[IngressUnit.scala 93:61]
  wire  _route_buffer_io_deq_ready_T_5 = _route_buffer_io_deq_ready_T_2 & _vcalloc_buffer_io_enq_valid_T_4; // @[IngressUnit.scala 94:37]
  wire  _route_buffer_io_deq_ready_T_7 = vcalloc_q_io_enq_ready | _vcalloc_buffer_io_enq_valid_T; // @[IngressUnit.scala 96:29]
  wire  _route_q_io_deq_ready_T = route_buffer_io_deq_ready & route_buffer_io_deq_valid; // @[Decoupled.scala 51:35]
  wire [3:0] c_lo = {vcalloc_q_io_deq_bits_vc_sel_0_3,vcalloc_q_io_deq_bits_vc_sel_0_2,vcalloc_q_io_deq_bits_vc_sel_0_1,
    vcalloc_q_io_deq_bits_vc_sel_0_0}; // @[IngressUnit.scala 107:41]
  wire [8:0] _c_T = {vcalloc_q_io_deq_bits_vc_sel_2_0,vcalloc_q_io_deq_bits_vc_sel_1_3,vcalloc_q_io_deq_bits_vc_sel_1_2,
    vcalloc_q_io_deq_bits_vc_sel_1_1,vcalloc_q_io_deq_bits_vc_sel_1_0,vcalloc_q_io_deq_bits_vc_sel_0_3,
    vcalloc_q_io_deq_bits_vc_sel_0_2,vcalloc_q_io_deq_bits_vc_sel_0_1,vcalloc_q_io_deq_bits_vc_sel_0_0}; // @[IngressUnit.scala 107:41]
  wire [8:0] _c_T_1 = {io_out_credit_available_2_0,io_out_credit_available_1_3,io_out_credit_available_1_2,
    io_out_credit_available_1_1,io_out_credit_available_1_0,io_out_credit_available_0_3,io_out_credit_available_0_2,
    io_out_credit_available_0_1,io_out_credit_available_0_0}; // @[IngressUnit.scala 107:74]
  wire [8:0] _c_T_2 = _c_T & _c_T_1; // @[IngressUnit.scala 107:48]
  wire  c = _c_T_2 != 9'h0; // @[IngressUnit.scala 107:82]
  wire  _vcalloc_q_io_deq_ready_T = vcalloc_buffer_io_deq_ready & vcalloc_buffer_io_deq_valid; // @[Decoupled.scala 51:35]
  reg  out_bundle_valid; // @[IngressUnit.scala 116:8]
  reg  out_bundle_bits_flit_head; // @[IngressUnit.scala 116:8]
  reg  out_bundle_bits_flit_tail; // @[IngressUnit.scala 116:8]
  reg [63:0] out_bundle_bits_flit_payload; // @[IngressUnit.scala 116:8]
  reg [1:0] out_bundle_bits_flit_flow_ingress_node; // @[IngressUnit.scala 116:8]
  reg [1:0] out_bundle_bits_flit_flow_egress_node; // @[IngressUnit.scala 116:8]
  reg [1:0] out_bundle_bits_out_virt_channel; // @[IngressUnit.scala 116:8]
  wire  out_channel_oh_0 = vcalloc_q_io_deq_bits_vc_sel_0_0 | vcalloc_q_io_deq_bits_vc_sel_0_1 |
    vcalloc_q_io_deq_bits_vc_sel_0_2 | vcalloc_q_io_deq_bits_vc_sel_0_3; // @[IngressUnit.scala 123:67]
  wire  out_channel_oh_1 = vcalloc_q_io_deq_bits_vc_sel_1_0 | vcalloc_q_io_deq_bits_vc_sel_1_1 |
    vcalloc_q_io_deq_bits_vc_sel_1_2 | vcalloc_q_io_deq_bits_vc_sel_1_3; // @[IngressUnit.scala 123:67]
  wire [1:0] out_bundle_bits_out_virt_channel_hi_1 = c_lo[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] out_bundle_bits_out_virt_channel_lo_1 = c_lo[1:0]; // @[OneHot.scala 31:18]
  wire  _out_bundle_bits_out_virt_channel_T_1 = |out_bundle_bits_out_virt_channel_hi_1; // @[OneHot.scala 32:14]
  wire [1:0] _out_bundle_bits_out_virt_channel_T_2 = out_bundle_bits_out_virt_channel_hi_1 |
    out_bundle_bits_out_virt_channel_lo_1; // @[OneHot.scala 32:28]
  wire [1:0] _out_bundle_bits_out_virt_channel_T_4 = {_out_bundle_bits_out_virt_channel_T_1,
    _out_bundle_bits_out_virt_channel_T_2[1]}; // @[Cat.scala 33:92]
  wire [3:0] _out_bundle_bits_out_virt_channel_T_5 = {vcalloc_q_io_deq_bits_vc_sel_1_3,vcalloc_q_io_deq_bits_vc_sel_1_2,
    vcalloc_q_io_deq_bits_vc_sel_1_1,vcalloc_q_io_deq_bits_vc_sel_1_0}; // @[OneHot.scala 22:45]
  wire [1:0] out_bundle_bits_out_virt_channel_hi_3 = _out_bundle_bits_out_virt_channel_T_5[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] out_bundle_bits_out_virt_channel_lo_3 = _out_bundle_bits_out_virt_channel_T_5[1:0]; // @[OneHot.scala 31:18]
  wire  _out_bundle_bits_out_virt_channel_T_6 = |out_bundle_bits_out_virt_channel_hi_3; // @[OneHot.scala 32:14]
  wire [1:0] _out_bundle_bits_out_virt_channel_T_7 = out_bundle_bits_out_virt_channel_hi_3 |
    out_bundle_bits_out_virt_channel_lo_3; // @[OneHot.scala 32:28]
  wire [1:0] _out_bundle_bits_out_virt_channel_T_9 = {_out_bundle_bits_out_virt_channel_T_6,
    _out_bundle_bits_out_virt_channel_T_7[1]}; // @[Cat.scala 33:92]
  wire [1:0] _out_bundle_bits_out_virt_channel_T_10 = out_channel_oh_0 ? _out_bundle_bits_out_virt_channel_T_4 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _out_bundle_bits_out_virt_channel_T_11 = out_channel_oh_1 ? _out_bundle_bits_out_virt_channel_T_9 : 2'h0; // @[Mux.scala 27:73]
  Queue_8 route_buffer ( // @[IngressUnit.scala 26:28]
    .clock(route_buffer_clock),
    .reset(route_buffer_reset),
    .io_enq_ready(route_buffer_io_enq_ready),
    .io_enq_valid(route_buffer_io_enq_valid),
    .io_enq_bits_head(route_buffer_io_enq_bits_head),
    .io_enq_bits_tail(route_buffer_io_enq_bits_tail),
    .io_enq_bits_payload(route_buffer_io_enq_bits_payload),
    .io_enq_bits_flow_ingress_node(route_buffer_io_enq_bits_flow_ingress_node),
    .io_enq_bits_flow_egress_node(route_buffer_io_enq_bits_flow_egress_node),
    .io_deq_ready(route_buffer_io_deq_ready),
    .io_deq_valid(route_buffer_io_deq_valid),
    .io_deq_bits_head(route_buffer_io_deq_bits_head),
    .io_deq_bits_tail(route_buffer_io_deq_bits_tail),
    .io_deq_bits_payload(route_buffer_io_deq_bits_payload),
    .io_deq_bits_flow_ingress_node(route_buffer_io_deq_bits_flow_ingress_node),
    .io_deq_bits_flow_egress_node(route_buffer_io_deq_bits_flow_egress_node)
  );
  Queue_9 route_q ( // @[IngressUnit.scala 27:23]
    .clock(route_q_clock),
    .reset(route_q_reset),
    .io_enq_ready(route_q_io_enq_ready),
    .io_enq_valid(route_q_io_enq_valid),
    .io_enq_bits_vc_sel_2_0(route_q_io_enq_bits_vc_sel_2_0),
    .io_enq_bits_vc_sel_1_0(route_q_io_enq_bits_vc_sel_1_0),
    .io_enq_bits_vc_sel_1_1(route_q_io_enq_bits_vc_sel_1_1),
    .io_enq_bits_vc_sel_1_2(route_q_io_enq_bits_vc_sel_1_2),
    .io_enq_bits_vc_sel_1_3(route_q_io_enq_bits_vc_sel_1_3),
    .io_enq_bits_vc_sel_0_0(route_q_io_enq_bits_vc_sel_0_0),
    .io_enq_bits_vc_sel_0_1(route_q_io_enq_bits_vc_sel_0_1),
    .io_enq_bits_vc_sel_0_2(route_q_io_enq_bits_vc_sel_0_2),
    .io_enq_bits_vc_sel_0_3(route_q_io_enq_bits_vc_sel_0_3),
    .io_deq_ready(route_q_io_deq_ready),
    .io_deq_valid(route_q_io_deq_valid),
    .io_deq_bits_vc_sel_2_0(route_q_io_deq_bits_vc_sel_2_0),
    .io_deq_bits_vc_sel_1_0(route_q_io_deq_bits_vc_sel_1_0),
    .io_deq_bits_vc_sel_1_1(route_q_io_deq_bits_vc_sel_1_1),
    .io_deq_bits_vc_sel_1_2(route_q_io_deq_bits_vc_sel_1_2),
    .io_deq_bits_vc_sel_1_3(route_q_io_deq_bits_vc_sel_1_3),
    .io_deq_bits_vc_sel_0_0(route_q_io_deq_bits_vc_sel_0_0),
    .io_deq_bits_vc_sel_0_1(route_q_io_deq_bits_vc_sel_0_1),
    .io_deq_bits_vc_sel_0_2(route_q_io_deq_bits_vc_sel_0_2),
    .io_deq_bits_vc_sel_0_3(route_q_io_deq_bits_vc_sel_0_3)
  );
  Queue_8 vcalloc_buffer ( // @[IngressUnit.scala 75:30]
    .clock(vcalloc_buffer_clock),
    .reset(vcalloc_buffer_reset),
    .io_enq_ready(vcalloc_buffer_io_enq_ready),
    .io_enq_valid(vcalloc_buffer_io_enq_valid),
    .io_enq_bits_head(vcalloc_buffer_io_enq_bits_head),
    .io_enq_bits_tail(vcalloc_buffer_io_enq_bits_tail),
    .io_enq_bits_payload(vcalloc_buffer_io_enq_bits_payload),
    .io_enq_bits_flow_ingress_node(vcalloc_buffer_io_enq_bits_flow_ingress_node),
    .io_enq_bits_flow_egress_node(vcalloc_buffer_io_enq_bits_flow_egress_node),
    .io_deq_ready(vcalloc_buffer_io_deq_ready),
    .io_deq_valid(vcalloc_buffer_io_deq_valid),
    .io_deq_bits_head(vcalloc_buffer_io_deq_bits_head),
    .io_deq_bits_tail(vcalloc_buffer_io_deq_bits_tail),
    .io_deq_bits_payload(vcalloc_buffer_io_deq_bits_payload),
    .io_deq_bits_flow_ingress_node(vcalloc_buffer_io_deq_bits_flow_ingress_node),
    .io_deq_bits_flow_egress_node(vcalloc_buffer_io_deq_bits_flow_egress_node)
  );
  Queue_11 vcalloc_q ( // @[IngressUnit.scala 76:25]
    .clock(vcalloc_q_clock),
    .reset(vcalloc_q_reset),
    .io_enq_ready(vcalloc_q_io_enq_ready),
    .io_enq_valid(vcalloc_q_io_enq_valid),
    .io_enq_bits_vc_sel_2_0(vcalloc_q_io_enq_bits_vc_sel_2_0),
    .io_enq_bits_vc_sel_1_0(vcalloc_q_io_enq_bits_vc_sel_1_0),
    .io_enq_bits_vc_sel_1_1(vcalloc_q_io_enq_bits_vc_sel_1_1),
    .io_enq_bits_vc_sel_1_2(vcalloc_q_io_enq_bits_vc_sel_1_2),
    .io_enq_bits_vc_sel_1_3(vcalloc_q_io_enq_bits_vc_sel_1_3),
    .io_enq_bits_vc_sel_0_0(vcalloc_q_io_enq_bits_vc_sel_0_0),
    .io_enq_bits_vc_sel_0_1(vcalloc_q_io_enq_bits_vc_sel_0_1),
    .io_enq_bits_vc_sel_0_2(vcalloc_q_io_enq_bits_vc_sel_0_2),
    .io_enq_bits_vc_sel_0_3(vcalloc_q_io_enq_bits_vc_sel_0_3),
    .io_deq_ready(vcalloc_q_io_deq_ready),
    .io_deq_valid(vcalloc_q_io_deq_valid),
    .io_deq_bits_vc_sel_2_0(vcalloc_q_io_deq_bits_vc_sel_2_0),
    .io_deq_bits_vc_sel_1_0(vcalloc_q_io_deq_bits_vc_sel_1_0),
    .io_deq_bits_vc_sel_1_1(vcalloc_q_io_deq_bits_vc_sel_1_1),
    .io_deq_bits_vc_sel_1_2(vcalloc_q_io_deq_bits_vc_sel_1_2),
    .io_deq_bits_vc_sel_1_3(vcalloc_q_io_deq_bits_vc_sel_1_3),
    .io_deq_bits_vc_sel_0_0(vcalloc_q_io_deq_bits_vc_sel_0_0),
    .io_deq_bits_vc_sel_0_1(vcalloc_q_io_deq_bits_vc_sel_0_1),
    .io_deq_bits_vc_sel_0_2(vcalloc_q_io_deq_bits_vc_sel_0_2),
    .io_deq_bits_vc_sel_0_3(vcalloc_q_io_deq_bits_vc_sel_0_3)
  );
  assign io_router_req_valid = io_in_valid & route_buffer_io_enq_ready & io_in_bits_head & ~at_dest; // @[IngressUnit.scala 58:86]
  assign io_router_req_bits_flow_ingress_node = route_buffer_io_enq_bits_flow_ingress_node; // @[IngressUnit.scala 53:27]
  assign io_router_req_bits_flow_egress_node = route_buffer_io_enq_bits_flow_egress_node; // @[IngressUnit.scala 53:27]
  assign io_vcalloc_req_valid = _io_vcalloc_req_valid_T_1 & vcalloc_buffer_io_enq_ready & vcalloc_q_io_enq_ready; // @[IngressUnit.scala 92:41]
  assign io_vcalloc_req_bits_vc_sel_2_0 = route_q_io_deq_bits_vc_sel_2_0; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_1_0 = route_q_io_deq_bits_vc_sel_1_0; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_1_1 = route_q_io_deq_bits_vc_sel_1_1; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_1_2 = route_q_io_deq_bits_vc_sel_1_2; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_1_3 = route_q_io_deq_bits_vc_sel_1_3; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_0_0 = route_q_io_deq_bits_vc_sel_0_0; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_0_1 = route_q_io_deq_bits_vc_sel_0_1; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_0_2 = route_q_io_deq_bits_vc_sel_0_2; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_0_3 = route_q_io_deq_bits_vc_sel_0_3; // @[IngressUnit.scala 81:30]
  assign io_salloc_req_0_valid = vcalloc_buffer_io_deq_valid & vcalloc_q_io_deq_valid & c; // @[IngressUnit.scala 109:83]
  assign io_salloc_req_0_bits_vc_sel_2_0 = vcalloc_q_io_deq_bits_vc_sel_2_0; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_1_0 = vcalloc_q_io_deq_bits_vc_sel_1_0; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_1_1 = vcalloc_q_io_deq_bits_vc_sel_1_1; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_1_2 = vcalloc_q_io_deq_bits_vc_sel_1_2; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_1_3 = vcalloc_q_io_deq_bits_vc_sel_1_3; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_0_0 = vcalloc_q_io_deq_bits_vc_sel_0_0; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_0_1 = vcalloc_q_io_deq_bits_vc_sel_0_1; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_0_2 = vcalloc_q_io_deq_bits_vc_sel_0_2; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_0_3 = vcalloc_q_io_deq_bits_vc_sel_0_3; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_tail = vcalloc_buffer_io_deq_bits_tail; // @[IngressUnit.scala 105:30]
  assign io_out_0_valid = out_bundle_valid; // @[IngressUnit.scala 118:13]
  assign io_out_0_bits_flit_head = out_bundle_bits_flit_head; // @[IngressUnit.scala 118:13]
  assign io_out_0_bits_flit_tail = out_bundle_bits_flit_tail; // @[IngressUnit.scala 118:13]
  assign io_out_0_bits_flit_payload = out_bundle_bits_flit_payload; // @[IngressUnit.scala 118:13]
  assign io_out_0_bits_flit_flow_ingress_node = out_bundle_bits_flit_flow_ingress_node; // @[IngressUnit.scala 118:13]
  assign io_out_0_bits_flit_flow_egress_node = out_bundle_bits_flit_flow_egress_node; // @[IngressUnit.scala 118:13]
  assign io_out_0_bits_out_virt_channel = out_bundle_bits_out_virt_channel; // @[IngressUnit.scala 118:13]
  assign io_in_ready = route_buffer_io_enq_ready; // @[IngressUnit.scala 59:44]
  assign route_buffer_clock = clock;
  assign route_buffer_reset = reset;
  assign route_buffer_io_enq_valid = io_in_valid; // @[IngressUnit.scala 56:44]
  assign route_buffer_io_enq_bits_head = io_in_bits_head; // @[IngressUnit.scala 32:33]
  assign route_buffer_io_enq_bits_tail = io_in_bits_tail; // @[IngressUnit.scala 33:33]
  assign route_buffer_io_enq_bits_payload = io_in_bits_payload; // @[IngressUnit.scala 50:36]
  assign route_buffer_io_enq_bits_flow_ingress_node = 2'h2; // @[IngressUnit.scala 38:51]
  assign route_buffer_io_enq_bits_flow_egress_node = _route_buffer_io_enq_bits_flow_egress_node_T_9 |
    _route_buffer_io_enq_bits_flow_egress_node_T_7; // @[Mux.scala 27:73]
  assign route_buffer_io_deq_ready = _route_buffer_io_deq_ready_T_5 & _route_buffer_io_deq_ready_T_7; // @[IngressUnit.scala 95:37]
  assign route_q_clock = clock;
  assign route_q_reset = reset;
  assign route_q_io_enq_valid = _T_13 & io_in_bits_head & at_dest | io_router_req_valid; // @[IngressUnit.scala 62:24 64:53 65:26]
  assign route_q_io_enq_bits_vc_sel_2_0 = _T_13 & io_in_bits_head & at_dest & _T_2; // @[IngressUnit.scala 63:23 64:53]
  assign route_q_io_enq_bits_vc_sel_1_0 = _T_13 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_1_0; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_1_1 = _T_13 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_1_1; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_1_2 = _T_13 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_1_2; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_1_3 = _T_13 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_1_3; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_0_0 = _T_13 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_0_0; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_0_1 = _T_13 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_0_1; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_0_2 = _T_13 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_0_2; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_0_3 = _T_13 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_0_3; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_deq_ready = _route_q_io_deq_ready_T & route_buffer_io_deq_bits_tail; // @[IngressUnit.scala 97:55]
  assign vcalloc_buffer_clock = clock;
  assign vcalloc_buffer_reset = reset;
  assign vcalloc_buffer_io_enq_valid = _vcalloc_buffer_io_enq_valid_T_2 & _vcalloc_buffer_io_enq_valid_T_4; // @[IngressUnit.scala 88:37]
  assign vcalloc_buffer_io_enq_bits_head = route_buffer_io_deq_bits_head; // @[IngressUnit.scala 79:30]
  assign vcalloc_buffer_io_enq_bits_tail = route_buffer_io_deq_bits_tail; // @[IngressUnit.scala 79:30]
  assign vcalloc_buffer_io_enq_bits_payload = route_buffer_io_deq_bits_payload; // @[IngressUnit.scala 79:30]
  assign vcalloc_buffer_io_enq_bits_flow_ingress_node = route_buffer_io_deq_bits_flow_ingress_node; // @[IngressUnit.scala 79:30]
  assign vcalloc_buffer_io_enq_bits_flow_egress_node = route_buffer_io_deq_bits_flow_egress_node; // @[IngressUnit.scala 79:30]
  assign vcalloc_buffer_io_deq_ready = io_salloc_req_0_ready & vcalloc_q_io_deq_valid & c; // @[IngressUnit.scala 110:83]
  assign vcalloc_q_clock = clock;
  assign vcalloc_q_reset = reset;
  assign vcalloc_q_io_enq_valid = io_vcalloc_req_ready & io_vcalloc_req_valid; // @[Decoupled.scala 51:35]
  assign vcalloc_q_io_enq_bits_vc_sel_2_0 = io_vcalloc_resp_vc_sel_2_0; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_1_0 = io_vcalloc_resp_vc_sel_1_0; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_1_1 = io_vcalloc_resp_vc_sel_1_1; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_1_2 = io_vcalloc_resp_vc_sel_1_2; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_1_3 = io_vcalloc_resp_vc_sel_1_3; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_0_0 = io_vcalloc_resp_vc_sel_0_0; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_0_1 = io_vcalloc_resp_vc_sel_0_1; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_0_2 = io_vcalloc_resp_vc_sel_0_2; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_0_3 = io_vcalloc_resp_vc_sel_0_3; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_deq_ready = vcalloc_buffer_io_deq_bits_tail & _vcalloc_q_io_deq_ready_T; // @[IngressUnit.scala 111:42]
  always @(posedge clock) begin
    out_bundle_valid <= vcalloc_buffer_io_deq_ready & vcalloc_buffer_io_deq_valid; // @[Decoupled.scala 51:35]
    out_bundle_bits_flit_head <= vcalloc_buffer_io_deq_bits_head; // @[IngressUnit.scala 121:24]
    out_bundle_bits_flit_tail <= vcalloc_buffer_io_deq_bits_tail; // @[IngressUnit.scala 121:24]
    out_bundle_bits_flit_payload <= vcalloc_buffer_io_deq_bits_payload; // @[IngressUnit.scala 121:24]
    out_bundle_bits_flit_flow_ingress_node <= vcalloc_buffer_io_deq_bits_flow_ingress_node; // @[IngressUnit.scala 121:24]
    out_bundle_bits_flit_flow_egress_node <= vcalloc_buffer_io_deq_bits_flow_egress_node; // @[IngressUnit.scala 121:24]
    out_bundle_bits_out_virt_channel <= _out_bundle_bits_out_virt_channel_T_10 | _out_bundle_bits_out_virt_channel_T_11; // @[Mux.scala 27:73]
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~(io_in_valid & ~_T_6))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at IngressUnit.scala:30 assert(!(io.in.valid && !cParam.possibleFlows.toSeq.map(_.egressId.U === io.in.bits.egress_id).orR))\n"
            ); // @[IngressUnit.scala 30:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_11 & ~(~(route_q_io_enq_valid & ~route_q_io_enq_ready))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at IngressUnit.scala:73 assert(!(route_q.io.enq.valid && !route_q.io.enq.ready))\n"); // @[IngressUnit.scala 73:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_11 & ~(~(vcalloc_q_io_enq_valid & ~vcalloc_q_io_enq_ready))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at IngressUnit.scala:102 assert(!(vcalloc_q.io.enq.valid && !vcalloc_q.io.enq.ready))\n"
            ); // @[IngressUnit.scala 102:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  out_bundle_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  out_bundle_bits_flit_head = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  out_bundle_bits_flit_tail = _RAND_2[0:0];
  _RAND_3 = {2{`RANDOM}};
  out_bundle_bits_flit_payload = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  out_bundle_bits_flit_flow_ingress_node = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  out_bundle_bits_flit_flow_egress_node = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  out_bundle_bits_out_virt_channel = _RAND_6[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(~(io_in_valid & ~_T_6)); // @[IngressUnit.scala 30:9]
    end
    //
    if (_T_11) begin
      assert(~(route_q_io_enq_valid & ~route_q_io_enq_ready)); // @[IngressUnit.scala 73:9]
    end
    //
    if (_T_11) begin
      assert(~(vcalloc_q_io_enq_valid & ~vcalloc_q_io_enq_ready)); // @[IngressUnit.scala 102:9]
    end
  end
endmodule
module RouteComputer_2(
  input  [1:0] io_req_2_bits_flow_ingress_node,
  input  [1:0] io_req_2_bits_flow_egress_node,
  input  [1:0] io_req_1_bits_src_virt_id,
  input  [1:0] io_req_1_bits_flow_ingress_node,
  input  [1:0] io_req_1_bits_flow_egress_node,
  input  [1:0] io_req_0_bits_src_virt_id,
  input  [1:0] io_req_0_bits_flow_ingress_node,
  input  [1:0] io_req_0_bits_flow_egress_node,
  output       io_resp_2_vc_sel_1_0,
  output       io_resp_2_vc_sel_1_1,
  output       io_resp_2_vc_sel_1_2,
  output       io_resp_2_vc_sel_1_3,
  output       io_resp_2_vc_sel_0_0,
  output       io_resp_2_vc_sel_0_1,
  output       io_resp_2_vc_sel_0_2,
  output       io_resp_2_vc_sel_0_3,
  output       io_resp_1_vc_sel_1_0,
  output       io_resp_1_vc_sel_1_1,
  output       io_resp_1_vc_sel_1_2,
  output       io_resp_1_vc_sel_1_3,
  output       io_resp_1_vc_sel_0_0,
  output       io_resp_1_vc_sel_0_1,
  output       io_resp_1_vc_sel_0_2,
  output       io_resp_1_vc_sel_0_3,
  output       io_resp_0_vc_sel_1_0,
  output       io_resp_0_vc_sel_1_1,
  output       io_resp_0_vc_sel_1_2,
  output       io_resp_0_vc_sel_1_3,
  output       io_resp_0_vc_sel_0_0,
  output       io_resp_0_vc_sel_0_1,
  output       io_resp_0_vc_sel_0_2,
  output       io_resp_0_vc_sel_0_3
);
  wire [5:0] addr = {io_req_0_bits_src_virt_id,io_req_0_bits_flow_ingress_node,io_req_0_bits_flow_egress_node}; // @[RouteComputer.scala 74:27]
  wire [5:0] decoded_invInputs = ~addr; // @[pla.scala 78:21]
  wire  decoded_andMatrixInput_0 = decoded_invInputs[4]; // @[pla.scala 91:29]
  wire  decoded_andMatrixInput_1 = decoded_invInputs[5]; // @[pla.scala 91:29]
  wire [1:0] _decoded_T = {decoded_andMatrixInput_0,decoded_andMatrixInput_1}; // @[Cat.scala 33:92]
  wire  _decoded_T_1 = &_decoded_T; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_0_1 = decoded_invInputs[0]; // @[pla.scala 91:29]
  wire  decoded_andMatrixInput_1_1 = decoded_invInputs[3]; // @[pla.scala 91:29]
  wire [3:0] _decoded_T_2 = {decoded_andMatrixInput_0_1,decoded_andMatrixInput_1_1,decoded_andMatrixInput_0,
    decoded_andMatrixInput_1}; // @[Cat.scala 33:92]
  wire  _decoded_T_3 = &_decoded_T_2; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_0_2 = addr[0]; // @[pla.scala 90:45]
  wire  decoded_andMatrixInput_1_2 = addr[1]; // @[pla.scala 90:45]
  wire [1:0] _decoded_T_4 = {decoded_andMatrixInput_0_2,decoded_andMatrixInput_1_2}; // @[Cat.scala 33:92]
  wire  _decoded_T_5 = &_decoded_T_4; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_1_3 = addr[4]; // @[pla.scala 90:45]
  wire [1:0] _decoded_T_6 = {decoded_andMatrixInput_1_2,decoded_andMatrixInput_1_3}; // @[Cat.scala 33:92]
  wire  _decoded_T_7 = &_decoded_T_6; // @[pla.scala 98:74]
  wire [3:0] _decoded_T_8 = {decoded_andMatrixInput_0_1,decoded_andMatrixInput_1_2,decoded_andMatrixInput_1_1,
    decoded_andMatrixInput_1_3}; // @[Cat.scala 33:92]
  wire  _decoded_T_9 = &_decoded_T_8; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_1_5 = addr[5]; // @[pla.scala 90:45]
  wire [1:0] _decoded_T_10 = {decoded_andMatrixInput_1_2,decoded_andMatrixInput_1_5}; // @[Cat.scala 33:92]
  wire  _decoded_T_11 = &_decoded_T_10; // @[pla.scala 98:74]
  wire [3:0] _decoded_T_12 = {decoded_andMatrixInput_0_1,decoded_andMatrixInput_1_2,decoded_andMatrixInput_1_1,
    decoded_andMatrixInput_1_5}; // @[Cat.scala 33:92]
  wire  _decoded_T_13 = &_decoded_T_12; // @[pla.scala 98:74]
  wire [1:0] _decoded_T_14 = {decoded_andMatrixInput_1_3,decoded_andMatrixInput_1_5}; // @[Cat.scala 33:92]
  wire  _decoded_T_15 = &_decoded_T_14; // @[pla.scala 98:74]
  wire [3:0] _decoded_T_16 = {decoded_andMatrixInput_0_1,decoded_andMatrixInput_1_1,decoded_andMatrixInput_1_3,
    decoded_andMatrixInput_1_5}; // @[Cat.scala 33:92]
  wire  _decoded_T_17 = &_decoded_T_16; // @[pla.scala 98:74]
  wire  _decoded_orMatrixOutputs_T = |_decoded_T_15; // @[pla.scala 114:39]
  wire  _decoded_orMatrixOutputs_T_1 = |_decoded_T_11; // @[pla.scala 114:39]
  wire [1:0] _decoded_orMatrixOutputs_T_2 = {_decoded_T_7,_decoded_T_11}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_3 = |_decoded_orMatrixOutputs_T_2; // @[pla.scala 114:39]
  wire [1:0] _decoded_orMatrixOutputs_T_4 = {_decoded_T_1,_decoded_T_5}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_5 = |_decoded_orMatrixOutputs_T_4; // @[pla.scala 114:39]
  wire  _decoded_orMatrixOutputs_T_6 = |_decoded_T_17; // @[pla.scala 114:39]
  wire  _decoded_orMatrixOutputs_T_7 = |_decoded_T_13; // @[pla.scala 114:39]
  wire [1:0] _decoded_orMatrixOutputs_T_8 = {_decoded_T_9,_decoded_T_13}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_9 = |_decoded_orMatrixOutputs_T_8; // @[pla.scala 114:39]
  wire  _decoded_orMatrixOutputs_T_10 = |_decoded_T_3; // @[pla.scala 114:39]
  wire [7:0] decoded_orMatrixOutputs = {_decoded_orMatrixOutputs_T_10,_decoded_orMatrixOutputs_T_9,
    _decoded_orMatrixOutputs_T_7,_decoded_orMatrixOutputs_T_6,_decoded_orMatrixOutputs_T_5,_decoded_orMatrixOutputs_T_3,
    _decoded_orMatrixOutputs_T_1,_decoded_orMatrixOutputs_T}; // @[Cat.scala 33:92]
  wire [7:0] decoded_invMatrixOutputs = {decoded_orMatrixOutputs[7],decoded_orMatrixOutputs[6],decoded_orMatrixOutputs[5
    ],decoded_orMatrixOutputs[4],decoded_orMatrixOutputs[3],decoded_orMatrixOutputs[2],decoded_orMatrixOutputs[1],
    decoded_orMatrixOutputs[0]}; // @[Cat.scala 33:92]
  wire [7:0] _GEN_0 = {{4'd0}, decoded_invMatrixOutputs[7:4]}; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_21 = _GEN_0 & 8'hf; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_23 = {decoded_invMatrixOutputs[3:0], 4'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _decoded_T_25 = _decoded_T_23 & 8'hf0; // @[Bitwise.scala 108:80]
  wire [7:0] _decoded_T_26 = _decoded_T_21 | _decoded_T_25; // @[Bitwise.scala 108:39]
  wire [7:0] _GEN_1 = {{2'd0}, _decoded_T_26[7:2]}; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_31 = _GEN_1 & 8'h33; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_33 = {_decoded_T_26[5:0], 2'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _decoded_T_35 = _decoded_T_33 & 8'hcc; // @[Bitwise.scala 108:80]
  wire [7:0] _decoded_T_36 = _decoded_T_31 | _decoded_T_35; // @[Bitwise.scala 108:39]
  wire [7:0] _GEN_2 = {{1'd0}, _decoded_T_36[7:1]}; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_41 = _GEN_2 & 8'h55; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_43 = {_decoded_T_36[6:0], 1'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _decoded_T_45 = _decoded_T_43 & 8'haa; // @[Bitwise.scala 108:80]
  wire [7:0] decoded = _decoded_T_41 | _decoded_T_45; // @[Bitwise.scala 108:39]
  wire [5:0] addr_1 = {io_req_1_bits_src_virt_id,io_req_1_bits_flow_ingress_node,io_req_1_bits_flow_egress_node}; // @[RouteComputer.scala 74:27]
  wire [5:0] decoded_invInputs_1 = ~addr_1; // @[pla.scala 78:21]
  wire  decoded_andMatrixInput_0_9 = decoded_invInputs_1[4]; // @[pla.scala 91:29]
  wire  decoded_andMatrixInput_1_9 = decoded_invInputs_1[5]; // @[pla.scala 91:29]
  wire [1:0] _decoded_T_46 = {decoded_andMatrixInput_0_9,decoded_andMatrixInput_1_9}; // @[Cat.scala 33:92]
  wire  _decoded_T_47 = &_decoded_T_46; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_0_10 = decoded_invInputs_1[3]; // @[pla.scala 91:29]
  wire [2:0] _decoded_T_48 = {decoded_andMatrixInput_0_10,decoded_andMatrixInput_0_9,decoded_andMatrixInput_1_9}; // @[Cat.scala 33:92]
  wire  _decoded_T_49 = &_decoded_T_48; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_0_11 = addr_1[0]; // @[pla.scala 90:45]
  wire  decoded_andMatrixInput_1_11 = decoded_invInputs_1[1]; // @[pla.scala 91:29]
  wire [1:0] _decoded_T_50 = {decoded_andMatrixInput_0_11,decoded_andMatrixInput_1_11}; // @[Cat.scala 33:92]
  wire  _decoded_T_51 = &_decoded_T_50; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_0_12 = addr_1[1]; // @[pla.scala 90:45]
  wire  decoded_andMatrixInput_1_12 = addr_1[2]; // @[pla.scala 90:45]
  wire  decoded_andMatrixInput_2_5 = addr_1[3]; // @[pla.scala 90:45]
  wire [4:0] _decoded_T_52 = {decoded_andMatrixInput_0_12,decoded_andMatrixInput_1_12,decoded_andMatrixInput_2_5,
    decoded_andMatrixInput_0_9,decoded_andMatrixInput_1_9}; // @[Cat.scala 33:92]
  wire  _decoded_T_53 = &_decoded_T_52; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_0_13 = decoded_invInputs_1[0]; // @[pla.scala 91:29]
  wire  decoded_andMatrixInput_1_13 = addr_1[4]; // @[pla.scala 90:45]
  wire [1:0] _decoded_T_54 = {decoded_andMatrixInput_0_13,decoded_andMatrixInput_1_13}; // @[Cat.scala 33:92]
  wire  _decoded_T_55 = &_decoded_T_54; // @[pla.scala 98:74]
  wire [1:0] _decoded_T_56 = {decoded_andMatrixInput_1_12,decoded_andMatrixInput_1_13}; // @[Cat.scala 33:92]
  wire  _decoded_T_57 = &_decoded_T_56; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_1_15 = addr_1[5]; // @[pla.scala 90:45]
  wire [1:0] _decoded_T_58 = {decoded_andMatrixInput_0_13,decoded_andMatrixInput_1_15}; // @[Cat.scala 33:92]
  wire  _decoded_T_59 = &_decoded_T_58; // @[pla.scala 98:74]
  wire [1:0] _decoded_T_60 = {decoded_andMatrixInput_1_12,decoded_andMatrixInput_1_15}; // @[Cat.scala 33:92]
  wire  _decoded_T_61 = &_decoded_T_60; // @[pla.scala 98:74]
  wire [1:0] _decoded_T_62 = {decoded_andMatrixInput_1_13,decoded_andMatrixInput_1_15}; // @[Cat.scala 33:92]
  wire  _decoded_T_63 = &_decoded_T_62; // @[pla.scala 98:74]
  wire [2:0] _decoded_T_64 = {decoded_andMatrixInput_0_10,decoded_andMatrixInput_1_13,decoded_andMatrixInput_1_15}; // @[Cat.scala 33:92]
  wire  _decoded_T_65 = &_decoded_T_64; // @[pla.scala 98:74]
  wire [4:0] _decoded_T_66 = {decoded_andMatrixInput_0_12,decoded_andMatrixInput_1_12,decoded_andMatrixInput_2_5,
    decoded_andMatrixInput_1_13,decoded_andMatrixInput_1_15}; // @[Cat.scala 33:92]
  wire  _decoded_T_67 = &_decoded_T_66; // @[pla.scala 98:74]
  wire [1:0] _decoded_orMatrixOutputs_T_11 = {_decoded_T_65,_decoded_T_67}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_12 = |_decoded_orMatrixOutputs_T_11; // @[pla.scala 114:39]
  wire  _decoded_orMatrixOutputs_T_13 = |_decoded_T_59; // @[pla.scala 114:39]
  wire [1:0] _decoded_orMatrixOutputs_T_14 = {_decoded_T_55,_decoded_T_59}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_15 = |_decoded_orMatrixOutputs_T_14; // @[pla.scala 114:39]
  wire [1:0] _decoded_orMatrixOutputs_T_16 = {_decoded_T_49,_decoded_T_53}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_17 = |_decoded_orMatrixOutputs_T_16; // @[pla.scala 114:39]
  wire  _decoded_orMatrixOutputs_T_18 = |_decoded_T_63; // @[pla.scala 114:39]
  wire [1:0] _decoded_orMatrixOutputs_T_19 = {_decoded_T_59,_decoded_T_61}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_20 = |_decoded_orMatrixOutputs_T_19; // @[pla.scala 114:39]
  wire [3:0] _decoded_orMatrixOutputs_T_21 = {_decoded_T_55,_decoded_T_57,_decoded_T_59,_decoded_T_61}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_22 = |_decoded_orMatrixOutputs_T_21; // @[pla.scala 114:39]
  wire [1:0] _decoded_orMatrixOutputs_T_23 = {_decoded_T_47,_decoded_T_51}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_24 = |_decoded_orMatrixOutputs_T_23; // @[pla.scala 114:39]
  wire [7:0] decoded_orMatrixOutputs_1 = {_decoded_orMatrixOutputs_T_24,_decoded_orMatrixOutputs_T_22,
    _decoded_orMatrixOutputs_T_20,_decoded_orMatrixOutputs_T_18,_decoded_orMatrixOutputs_T_17,
    _decoded_orMatrixOutputs_T_15,_decoded_orMatrixOutputs_T_13,_decoded_orMatrixOutputs_T_12}; // @[Cat.scala 33:92]
  wire [7:0] decoded_invMatrixOutputs_1 = {decoded_orMatrixOutputs_1[7],decoded_orMatrixOutputs_1[6],
    decoded_orMatrixOutputs_1[5],decoded_orMatrixOutputs_1[4],decoded_orMatrixOutputs_1[3],decoded_orMatrixOutputs_1[2],
    decoded_orMatrixOutputs_1[1],decoded_orMatrixOutputs_1[0]}; // @[Cat.scala 33:92]
  wire [7:0] _GEN_3 = {{4'd0}, decoded_invMatrixOutputs_1[7:4]}; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_71 = _GEN_3 & 8'hf; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_73 = {decoded_invMatrixOutputs_1[3:0], 4'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _decoded_T_75 = _decoded_T_73 & 8'hf0; // @[Bitwise.scala 108:80]
  wire [7:0] _decoded_T_76 = _decoded_T_71 | _decoded_T_75; // @[Bitwise.scala 108:39]
  wire [7:0] _GEN_4 = {{2'd0}, _decoded_T_76[7:2]}; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_81 = _GEN_4 & 8'h33; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_83 = {_decoded_T_76[5:0], 2'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _decoded_T_85 = _decoded_T_83 & 8'hcc; // @[Bitwise.scala 108:80]
  wire [7:0] _decoded_T_86 = _decoded_T_81 | _decoded_T_85; // @[Bitwise.scala 108:39]
  wire [7:0] _GEN_5 = {{1'd0}, _decoded_T_86[7:1]}; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_91 = _GEN_5 & 8'h55; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_93 = {_decoded_T_86[6:0], 1'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _decoded_T_95 = _decoded_T_93 & 8'haa; // @[Bitwise.scala 108:80]
  wire [7:0] decoded_1 = _decoded_T_91 | _decoded_T_95; // @[Bitwise.scala 108:39]
  wire [5:0] addr_2 = {2'h0,io_req_2_bits_flow_ingress_node,io_req_2_bits_flow_egress_node}; // @[RouteComputer.scala 74:27]
  wire [5:0] decoded_invInputs_2 = ~addr_2; // @[pla.scala 78:21]
  wire  decoded_andMatrixInput_0_20 = decoded_invInputs_2[0]; // @[pla.scala 91:29]
  wire  decoded_andMatrixInput_1_20 = decoded_invInputs_2[2]; // @[pla.scala 91:29]
  wire  decoded_andMatrixInput_2_8 = addr_2[3]; // @[pla.scala 90:45]
  wire  decoded_andMatrixInput_3_6 = decoded_invInputs_2[4]; // @[pla.scala 91:29]
  wire  decoded_andMatrixInput_4_2 = decoded_invInputs_2[5]; // @[pla.scala 91:29]
  wire [4:0] _decoded_T_96 = {decoded_andMatrixInput_0_20,decoded_andMatrixInput_1_20,decoded_andMatrixInput_2_8,
    decoded_andMatrixInput_3_6,decoded_andMatrixInput_4_2}; // @[Cat.scala 33:92]
  wire  _decoded_T_97 = &_decoded_T_96; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_0_21 = decoded_invInputs_2[1]; // @[pla.scala 91:29]
  wire [4:0] _decoded_T_98 = {decoded_andMatrixInput_0_21,decoded_andMatrixInput_1_20,decoded_andMatrixInput_2_8,
    decoded_andMatrixInput_3_6,decoded_andMatrixInput_4_2}; // @[Cat.scala 33:92]
  wire  _decoded_T_99 = &_decoded_T_98; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_0_22 = addr_2[1]; // @[pla.scala 90:45]
  wire [4:0] _decoded_T_100 = {decoded_andMatrixInput_0_22,decoded_andMatrixInput_1_20,decoded_andMatrixInput_2_8,
    decoded_andMatrixInput_3_6,decoded_andMatrixInput_4_2}; // @[Cat.scala 33:92]
  wire  _decoded_T_101 = &_decoded_T_100; // @[pla.scala 98:74]
  wire [1:0] _decoded_orMatrixOutputs_T_25 = {_decoded_T_97,_decoded_T_101}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_26 = |_decoded_orMatrixOutputs_T_25; // @[pla.scala 114:39]
  wire [1:0] _decoded_orMatrixOutputs_T_31 = {_decoded_T_97,_decoded_T_99}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_32 = |_decoded_orMatrixOutputs_T_31; // @[pla.scala 114:39]
  wire [7:0] decoded_orMatrixOutputs_2 = {1'h0,_decoded_orMatrixOutputs_T_32,_decoded_orMatrixOutputs_T_32,
    _decoded_orMatrixOutputs_T_32,1'h0,_decoded_orMatrixOutputs_T_26,_decoded_orMatrixOutputs_T_26,
    _decoded_orMatrixOutputs_T_26}; // @[Cat.scala 33:92]
  wire [7:0] decoded_invMatrixOutputs_2 = {decoded_orMatrixOutputs_2[7],decoded_orMatrixOutputs_2[6],
    decoded_orMatrixOutputs_2[5],decoded_orMatrixOutputs_2[4],decoded_orMatrixOutputs_2[3],decoded_orMatrixOutputs_2[2],
    decoded_orMatrixOutputs_2[1],decoded_orMatrixOutputs_2[0]}; // @[Cat.scala 33:92]
  wire [7:0] _GEN_6 = {{4'd0}, decoded_invMatrixOutputs_2[7:4]}; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_105 = _GEN_6 & 8'hf; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_107 = {decoded_invMatrixOutputs_2[3:0], 4'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _decoded_T_109 = _decoded_T_107 & 8'hf0; // @[Bitwise.scala 108:80]
  wire [7:0] _decoded_T_110 = _decoded_T_105 | _decoded_T_109; // @[Bitwise.scala 108:39]
  wire [7:0] _GEN_7 = {{2'd0}, _decoded_T_110[7:2]}; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_115 = _GEN_7 & 8'h33; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_117 = {_decoded_T_110[5:0], 2'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _decoded_T_119 = _decoded_T_117 & 8'hcc; // @[Bitwise.scala 108:80]
  wire [7:0] _decoded_T_120 = _decoded_T_115 | _decoded_T_119; // @[Bitwise.scala 108:39]
  wire [7:0] _GEN_8 = {{1'd0}, _decoded_T_120[7:1]}; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_125 = _GEN_8 & 8'h55; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_127 = {_decoded_T_120[6:0], 1'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _decoded_T_129 = _decoded_T_127 & 8'haa; // @[Bitwise.scala 108:80]
  wire [7:0] decoded_2 = _decoded_T_125 | _decoded_T_129; // @[Bitwise.scala 108:39]
  assign io_resp_2_vc_sel_1_0 = decoded_2[4]; // @[RouteComputer.scala 90:46]
  assign io_resp_2_vc_sel_1_1 = decoded_2[5]; // @[RouteComputer.scala 90:46]
  assign io_resp_2_vc_sel_1_2 = decoded_2[6]; // @[RouteComputer.scala 90:46]
  assign io_resp_2_vc_sel_1_3 = decoded_2[7]; // @[RouteComputer.scala 90:46]
  assign io_resp_2_vc_sel_0_0 = decoded_2[0]; // @[RouteComputer.scala 90:46]
  assign io_resp_2_vc_sel_0_1 = decoded_2[1]; // @[RouteComputer.scala 90:46]
  assign io_resp_2_vc_sel_0_2 = decoded_2[2]; // @[RouteComputer.scala 90:46]
  assign io_resp_2_vc_sel_0_3 = decoded_2[3]; // @[RouteComputer.scala 90:46]
  assign io_resp_1_vc_sel_1_0 = decoded_1[4]; // @[RouteComputer.scala 90:46]
  assign io_resp_1_vc_sel_1_1 = decoded_1[5]; // @[RouteComputer.scala 90:46]
  assign io_resp_1_vc_sel_1_2 = decoded_1[6]; // @[RouteComputer.scala 90:46]
  assign io_resp_1_vc_sel_1_3 = decoded_1[7]; // @[RouteComputer.scala 90:46]
  assign io_resp_1_vc_sel_0_0 = decoded_1[0]; // @[RouteComputer.scala 90:46]
  assign io_resp_1_vc_sel_0_1 = decoded_1[1]; // @[RouteComputer.scala 90:46]
  assign io_resp_1_vc_sel_0_2 = decoded_1[2]; // @[RouteComputer.scala 90:46]
  assign io_resp_1_vc_sel_0_3 = decoded_1[3]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_1_0 = decoded[4]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_1_1 = decoded[5]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_1_2 = decoded[6]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_1_3 = decoded[7]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_0_0 = decoded[0]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_0_1 = decoded[1]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_0_2 = decoded[2]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_0_3 = decoded[3]; // @[RouteComputer.scala 90:46]
endmodule
module Router_2(
  input         clock,
  input         reset,
  output [1:0]  auto_debug_out_va_stall_0,
  output [1:0]  auto_debug_out_va_stall_1,
  output [1:0]  auto_debug_out_sa_stall_0,
  output [1:0]  auto_debug_out_sa_stall_1,
  output        auto_egress_nodes_out_flit_valid,
  output        auto_egress_nodes_out_flit_bits_head,
  output        auto_egress_nodes_out_flit_bits_tail,
  output [63:0] auto_egress_nodes_out_flit_bits_payload,
  output [1:0]  auto_egress_nodes_out_flit_bits_ingress_id,
  output        auto_ingress_nodes_in_flit_ready,
  input         auto_ingress_nodes_in_flit_valid,
  input         auto_ingress_nodes_in_flit_bits_head,
  input         auto_ingress_nodes_in_flit_bits_tail,
  input  [63:0] auto_ingress_nodes_in_flit_bits_payload,
  input  [1:0]  auto_ingress_nodes_in_flit_bits_egress_id,
  output        auto_source_nodes_out_1_flit_0_valid,
  output        auto_source_nodes_out_1_flit_0_bits_head,
  output        auto_source_nodes_out_1_flit_0_bits_tail,
  output [63:0] auto_source_nodes_out_1_flit_0_bits_payload,
  output [1:0]  auto_source_nodes_out_1_flit_0_bits_flow_ingress_node,
  output [1:0]  auto_source_nodes_out_1_flit_0_bits_flow_egress_node,
  output [1:0]  auto_source_nodes_out_1_flit_0_bits_virt_channel_id,
  input  [3:0]  auto_source_nodes_out_1_credit_return,
  input  [3:0]  auto_source_nodes_out_1_vc_free,
  output        auto_source_nodes_out_0_flit_0_valid,
  output        auto_source_nodes_out_0_flit_0_bits_head,
  output        auto_source_nodes_out_0_flit_0_bits_tail,
  output [63:0] auto_source_nodes_out_0_flit_0_bits_payload,
  output [1:0]  auto_source_nodes_out_0_flit_0_bits_flow_ingress_node,
  output [1:0]  auto_source_nodes_out_0_flit_0_bits_flow_egress_node,
  output [1:0]  auto_source_nodes_out_0_flit_0_bits_virt_channel_id,
  input  [3:0]  auto_source_nodes_out_0_credit_return,
  input  [3:0]  auto_source_nodes_out_0_vc_free,
  input         auto_dest_nodes_in_1_flit_0_valid,
  input         auto_dest_nodes_in_1_flit_0_bits_head,
  input         auto_dest_nodes_in_1_flit_0_bits_tail,
  input  [63:0] auto_dest_nodes_in_1_flit_0_bits_payload,
  input  [1:0]  auto_dest_nodes_in_1_flit_0_bits_flow_ingress_node,
  input  [1:0]  auto_dest_nodes_in_1_flit_0_bits_flow_egress_node,
  input  [1:0]  auto_dest_nodes_in_1_flit_0_bits_virt_channel_id,
  output [3:0]  auto_dest_nodes_in_1_credit_return,
  output [3:0]  auto_dest_nodes_in_1_vc_free,
  input         auto_dest_nodes_in_0_flit_0_valid,
  input         auto_dest_nodes_in_0_flit_0_bits_head,
  input         auto_dest_nodes_in_0_flit_0_bits_tail,
  input  [63:0] auto_dest_nodes_in_0_flit_0_bits_payload,
  input  [1:0]  auto_dest_nodes_in_0_flit_0_bits_flow_ingress_node,
  input  [1:0]  auto_dest_nodes_in_0_flit_0_bits_flow_egress_node,
  input  [1:0]  auto_dest_nodes_in_0_flit_0_bits_virt_channel_id,
  output [3:0]  auto_dest_nodes_in_0_credit_return,
  output [3:0]  auto_dest_nodes_in_0_vc_free
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_REG_INIT
  wire  monitor_clock; // @[Nodes.scala 24:25]
  wire  monitor_reset; // @[Nodes.scala 24:25]
  wire  monitor_io_in_flit_0_valid; // @[Nodes.scala 24:25]
  wire  monitor_io_in_flit_0_bits_head; // @[Nodes.scala 24:25]
  wire  monitor_io_in_flit_0_bits_tail; // @[Nodes.scala 24:25]
  wire [1:0] monitor_io_in_flit_0_bits_flow_ingress_node; // @[Nodes.scala 24:25]
  wire [1:0] monitor_io_in_flit_0_bits_flow_egress_node; // @[Nodes.scala 24:25]
  wire [1:0] monitor_io_in_flit_0_bits_virt_channel_id; // @[Nodes.scala 24:25]
  wire  monitor_1_clock; // @[Nodes.scala 24:25]
  wire  monitor_1_reset; // @[Nodes.scala 24:25]
  wire  monitor_1_io_in_flit_0_valid; // @[Nodes.scala 24:25]
  wire  monitor_1_io_in_flit_0_bits_head; // @[Nodes.scala 24:25]
  wire  monitor_1_io_in_flit_0_bits_tail; // @[Nodes.scala 24:25]
  wire [1:0] monitor_1_io_in_flit_0_bits_flow_ingress_node; // @[Nodes.scala 24:25]
  wire [1:0] monitor_1_io_in_flit_0_bits_flow_egress_node; // @[Nodes.scala 24:25]
  wire [1:0] monitor_1_io_in_flit_0_bits_virt_channel_id; // @[Nodes.scala 24:25]
  wire  input_unit_0_from_1_clock; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_reset; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_router_req_valid; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_1_io_router_req_bits_src_virt_id; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_1_io_router_req_bits_flow_ingress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_1_io_router_req_bits_flow_egress_node; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_router_resp_vc_sel_1_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_router_resp_vc_sel_1_1; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_router_resp_vc_sel_1_2; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_router_resp_vc_sel_1_3; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_router_resp_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_router_resp_vc_sel_0_1; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_router_resp_vc_sel_0_2; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_router_resp_vc_sel_0_3; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_vcalloc_req_ready; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_vcalloc_req_valid; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_2_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_1_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_1_1; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_1_2; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_1_3; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_0_1; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_0_2; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_0_3; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_vcalloc_resp_vc_sel_2_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_vcalloc_resp_vc_sel_1_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_vcalloc_resp_vc_sel_1_1; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_vcalloc_resp_vc_sel_1_2; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_vcalloc_resp_vc_sel_1_3; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_vcalloc_resp_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_vcalloc_resp_vc_sel_0_1; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_vcalloc_resp_vc_sel_0_2; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_vcalloc_resp_vc_sel_0_3; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_out_credit_available_2_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_out_credit_available_1_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_out_credit_available_1_1; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_out_credit_available_1_2; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_out_credit_available_1_3; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_out_credit_available_0_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_out_credit_available_0_1; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_out_credit_available_0_2; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_out_credit_available_0_3; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_salloc_req_0_ready; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_salloc_req_0_valid; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_2_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_1_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_1_1; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_1_2; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_1_3; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_0_1; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_0_2; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_0_3; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_salloc_req_0_bits_tail; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_out_0_valid; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_out_0_bits_flit_head; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_out_0_bits_flit_tail; // @[Router.scala 112:13]
  wire [63:0] input_unit_0_from_1_io_out_0_bits_flit_payload; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_1_io_out_0_bits_flit_flow_ingress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_1_io_out_0_bits_flit_flow_egress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_1_io_out_0_bits_out_virt_channel; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_1_io_debug_va_stall; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_1_io_debug_sa_stall; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_in_flit_0_valid; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_in_flit_0_bits_head; // @[Router.scala 112:13]
  wire  input_unit_0_from_1_io_in_flit_0_bits_tail; // @[Router.scala 112:13]
  wire [63:0] input_unit_0_from_1_io_in_flit_0_bits_payload; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_1_io_in_flit_0_bits_flow_ingress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_1_io_in_flit_0_bits_flow_egress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_1_io_in_flit_0_bits_virt_channel_id; // @[Router.scala 112:13]
  wire [3:0] input_unit_0_from_1_io_in_credit_return; // @[Router.scala 112:13]
  wire [3:0] input_unit_0_from_1_io_in_vc_free; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_clock; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_reset; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_router_req_valid; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_3_io_router_req_bits_src_virt_id; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_3_io_router_req_bits_flow_ingress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_3_io_router_req_bits_flow_egress_node; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_router_resp_vc_sel_1_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_router_resp_vc_sel_1_1; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_router_resp_vc_sel_1_2; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_router_resp_vc_sel_1_3; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_router_resp_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_router_resp_vc_sel_0_1; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_router_resp_vc_sel_0_2; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_router_resp_vc_sel_0_3; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_vcalloc_req_ready; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_vcalloc_req_valid; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_2_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_1_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_1_1; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_1_2; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_1_3; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_0_1; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_0_2; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_0_3; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_vcalloc_resp_vc_sel_2_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_vcalloc_resp_vc_sel_1_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_vcalloc_resp_vc_sel_1_1; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_vcalloc_resp_vc_sel_1_2; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_vcalloc_resp_vc_sel_1_3; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_vcalloc_resp_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_vcalloc_resp_vc_sel_0_1; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_vcalloc_resp_vc_sel_0_2; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_vcalloc_resp_vc_sel_0_3; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_out_credit_available_2_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_out_credit_available_1_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_out_credit_available_1_1; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_out_credit_available_1_2; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_out_credit_available_1_3; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_out_credit_available_0_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_out_credit_available_0_1; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_out_credit_available_0_2; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_out_credit_available_0_3; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_salloc_req_0_ready; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_salloc_req_0_valid; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_2_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_1_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_1_1; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_1_2; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_1_3; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_0_1; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_0_2; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_0_3; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_salloc_req_0_bits_tail; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_out_0_valid; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_out_0_bits_flit_head; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_out_0_bits_flit_tail; // @[Router.scala 112:13]
  wire [63:0] input_unit_1_from_3_io_out_0_bits_flit_payload; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_3_io_out_0_bits_flit_flow_ingress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_3_io_out_0_bits_flit_flow_egress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_3_io_out_0_bits_out_virt_channel; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_3_io_debug_va_stall; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_3_io_debug_sa_stall; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_in_flit_0_valid; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_in_flit_0_bits_head; // @[Router.scala 112:13]
  wire  input_unit_1_from_3_io_in_flit_0_bits_tail; // @[Router.scala 112:13]
  wire [63:0] input_unit_1_from_3_io_in_flit_0_bits_payload; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_3_io_in_flit_0_bits_flow_ingress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_3_io_in_flit_0_bits_flow_egress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_3_io_in_flit_0_bits_virt_channel_id; // @[Router.scala 112:13]
  wire [3:0] input_unit_1_from_3_io_in_credit_return; // @[Router.scala 112:13]
  wire [3:0] input_unit_1_from_3_io_in_vc_free; // @[Router.scala 112:13]
  wire  ingress_unit_2_from_2_clock; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_reset; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_router_req_valid; // @[Router.scala 116:13]
  wire [1:0] ingress_unit_2_from_2_io_router_req_bits_flow_ingress_node; // @[Router.scala 116:13]
  wire [1:0] ingress_unit_2_from_2_io_router_req_bits_flow_egress_node; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_router_resp_vc_sel_1_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_router_resp_vc_sel_1_1; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_router_resp_vc_sel_1_2; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_router_resp_vc_sel_1_3; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_router_resp_vc_sel_0_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_router_resp_vc_sel_0_1; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_router_resp_vc_sel_0_2; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_router_resp_vc_sel_0_3; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_vcalloc_req_ready; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_vcalloc_req_valid; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_vcalloc_req_bits_vc_sel_2_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_vcalloc_req_bits_vc_sel_1_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_vcalloc_req_bits_vc_sel_1_1; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_vcalloc_req_bits_vc_sel_1_2; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_vcalloc_req_bits_vc_sel_1_3; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_vcalloc_req_bits_vc_sel_0_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_vcalloc_req_bits_vc_sel_0_1; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_vcalloc_req_bits_vc_sel_0_2; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_vcalloc_req_bits_vc_sel_0_3; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_vcalloc_resp_vc_sel_2_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_vcalloc_resp_vc_sel_1_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_vcalloc_resp_vc_sel_1_1; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_vcalloc_resp_vc_sel_1_2; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_vcalloc_resp_vc_sel_1_3; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_vcalloc_resp_vc_sel_0_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_vcalloc_resp_vc_sel_0_1; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_vcalloc_resp_vc_sel_0_2; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_vcalloc_resp_vc_sel_0_3; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_out_credit_available_2_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_out_credit_available_1_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_out_credit_available_1_1; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_out_credit_available_1_2; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_out_credit_available_1_3; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_out_credit_available_0_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_out_credit_available_0_1; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_out_credit_available_0_2; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_out_credit_available_0_3; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_salloc_req_0_ready; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_salloc_req_0_valid; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_salloc_req_0_bits_vc_sel_2_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_salloc_req_0_bits_vc_sel_1_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_salloc_req_0_bits_vc_sel_1_1; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_salloc_req_0_bits_vc_sel_1_2; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_salloc_req_0_bits_vc_sel_1_3; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_salloc_req_0_bits_vc_sel_0_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_salloc_req_0_bits_vc_sel_0_1; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_salloc_req_0_bits_vc_sel_0_2; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_salloc_req_0_bits_vc_sel_0_3; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_salloc_req_0_bits_tail; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_out_0_valid; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_out_0_bits_flit_head; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_out_0_bits_flit_tail; // @[Router.scala 116:13]
  wire [63:0] ingress_unit_2_from_2_io_out_0_bits_flit_payload; // @[Router.scala 116:13]
  wire [1:0] ingress_unit_2_from_2_io_out_0_bits_flit_flow_ingress_node; // @[Router.scala 116:13]
  wire [1:0] ingress_unit_2_from_2_io_out_0_bits_flit_flow_egress_node; // @[Router.scala 116:13]
  wire [1:0] ingress_unit_2_from_2_io_out_0_bits_out_virt_channel; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_in_ready; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_in_valid; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_in_bits_head; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_2_io_in_bits_tail; // @[Router.scala 116:13]
  wire [63:0] ingress_unit_2_from_2_io_in_bits_payload; // @[Router.scala 116:13]
  wire [1:0] ingress_unit_2_from_2_io_in_bits_egress_id; // @[Router.scala 116:13]
  wire  output_unit_0_to_1_clock; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_reset; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_in_0_valid; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_in_0_bits_head; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_in_0_bits_tail; // @[Router.scala 122:13]
  wire [63:0] output_unit_0_to_1_io_in_0_bits_payload; // @[Router.scala 122:13]
  wire [1:0] output_unit_0_to_1_io_in_0_bits_flow_ingress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_0_to_1_io_in_0_bits_flow_egress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_0_to_1_io_in_0_bits_virt_channel_id; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_credit_available_0; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_credit_available_1; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_credit_available_2; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_credit_available_3; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_channel_status_0_occupied; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_channel_status_1_occupied; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_channel_status_2_occupied; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_channel_status_3_occupied; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_allocs_0_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_allocs_1_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_allocs_2_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_allocs_3_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_credit_alloc_0_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_credit_alloc_1_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_credit_alloc_2_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_credit_alloc_3_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_out_flit_0_valid; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_out_flit_0_bits_head; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_out_flit_0_bits_tail; // @[Router.scala 122:13]
  wire [63:0] output_unit_0_to_1_io_out_flit_0_bits_payload; // @[Router.scala 122:13]
  wire [1:0] output_unit_0_to_1_io_out_flit_0_bits_flow_ingress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_0_to_1_io_out_flit_0_bits_flow_egress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_0_to_1_io_out_flit_0_bits_virt_channel_id; // @[Router.scala 122:13]
  wire [3:0] output_unit_0_to_1_io_out_credit_return; // @[Router.scala 122:13]
  wire [3:0] output_unit_0_to_1_io_out_vc_free; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_clock; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_reset; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_in_0_valid; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_in_0_bits_head; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_in_0_bits_tail; // @[Router.scala 122:13]
  wire [63:0] output_unit_1_to_3_io_in_0_bits_payload; // @[Router.scala 122:13]
  wire [1:0] output_unit_1_to_3_io_in_0_bits_flow_ingress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_1_to_3_io_in_0_bits_flow_egress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_1_to_3_io_in_0_bits_virt_channel_id; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_credit_available_0; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_credit_available_1; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_credit_available_2; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_credit_available_3; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_channel_status_0_occupied; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_channel_status_1_occupied; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_channel_status_2_occupied; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_channel_status_3_occupied; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_allocs_0_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_allocs_1_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_allocs_2_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_allocs_3_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_credit_alloc_0_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_credit_alloc_1_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_credit_alloc_2_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_credit_alloc_3_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_out_flit_0_valid; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_out_flit_0_bits_head; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_out_flit_0_bits_tail; // @[Router.scala 122:13]
  wire [63:0] output_unit_1_to_3_io_out_flit_0_bits_payload; // @[Router.scala 122:13]
  wire [1:0] output_unit_1_to_3_io_out_flit_0_bits_flow_ingress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_1_to_3_io_out_flit_0_bits_flow_egress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_1_to_3_io_out_flit_0_bits_virt_channel_id; // @[Router.scala 122:13]
  wire [3:0] output_unit_1_to_3_io_out_credit_return; // @[Router.scala 122:13]
  wire [3:0] output_unit_1_to_3_io_out_vc_free; // @[Router.scala 122:13]
  wire  egress_unit_2_to_2_clock; // @[Router.scala 125:13]
  wire  egress_unit_2_to_2_reset; // @[Router.scala 125:13]
  wire  egress_unit_2_to_2_io_in_0_valid; // @[Router.scala 125:13]
  wire  egress_unit_2_to_2_io_in_0_bits_head; // @[Router.scala 125:13]
  wire  egress_unit_2_to_2_io_in_0_bits_tail; // @[Router.scala 125:13]
  wire [63:0] egress_unit_2_to_2_io_in_0_bits_payload; // @[Router.scala 125:13]
  wire [1:0] egress_unit_2_to_2_io_in_0_bits_flow_ingress_node; // @[Router.scala 125:13]
  wire  egress_unit_2_to_2_io_credit_available_0; // @[Router.scala 125:13]
  wire  egress_unit_2_to_2_io_channel_status_0_occupied; // @[Router.scala 125:13]
  wire  egress_unit_2_to_2_io_allocs_0_alloc; // @[Router.scala 125:13]
  wire  egress_unit_2_to_2_io_credit_alloc_0_alloc; // @[Router.scala 125:13]
  wire  egress_unit_2_to_2_io_credit_alloc_0_tail; // @[Router.scala 125:13]
  wire  egress_unit_2_to_2_io_out_valid; // @[Router.scala 125:13]
  wire  egress_unit_2_to_2_io_out_bits_head; // @[Router.scala 125:13]
  wire  egress_unit_2_to_2_io_out_bits_tail; // @[Router.scala 125:13]
  wire [63:0] egress_unit_2_to_2_io_out_bits_payload; // @[Router.scala 125:13]
  wire [1:0] egress_unit_2_to_2_io_out_bits_ingress_id; // @[Router.scala 125:13]
  wire  switch_clock; // @[Router.scala 129:24]
  wire  switch_reset; // @[Router.scala 129:24]
  wire  switch_io_in_2_0_valid; // @[Router.scala 129:24]
  wire  switch_io_in_2_0_bits_flit_head; // @[Router.scala 129:24]
  wire  switch_io_in_2_0_bits_flit_tail; // @[Router.scala 129:24]
  wire [63:0] switch_io_in_2_0_bits_flit_payload; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_2_0_bits_flit_flow_ingress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_2_0_bits_flit_flow_egress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_2_0_bits_out_virt_channel; // @[Router.scala 129:24]
  wire  switch_io_in_1_0_valid; // @[Router.scala 129:24]
  wire  switch_io_in_1_0_bits_flit_head; // @[Router.scala 129:24]
  wire  switch_io_in_1_0_bits_flit_tail; // @[Router.scala 129:24]
  wire [63:0] switch_io_in_1_0_bits_flit_payload; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_1_0_bits_flit_flow_ingress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_1_0_bits_flit_flow_egress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_1_0_bits_out_virt_channel; // @[Router.scala 129:24]
  wire  switch_io_in_0_0_valid; // @[Router.scala 129:24]
  wire  switch_io_in_0_0_bits_flit_head; // @[Router.scala 129:24]
  wire  switch_io_in_0_0_bits_flit_tail; // @[Router.scala 129:24]
  wire [63:0] switch_io_in_0_0_bits_flit_payload; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_0_0_bits_flit_flow_ingress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_0_0_bits_flit_flow_egress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_0_0_bits_out_virt_channel; // @[Router.scala 129:24]
  wire  switch_io_out_2_0_valid; // @[Router.scala 129:24]
  wire  switch_io_out_2_0_bits_head; // @[Router.scala 129:24]
  wire  switch_io_out_2_0_bits_tail; // @[Router.scala 129:24]
  wire [63:0] switch_io_out_2_0_bits_payload; // @[Router.scala 129:24]
  wire [1:0] switch_io_out_2_0_bits_flow_ingress_node; // @[Router.scala 129:24]
  wire  switch_io_out_1_0_valid; // @[Router.scala 129:24]
  wire  switch_io_out_1_0_bits_head; // @[Router.scala 129:24]
  wire  switch_io_out_1_0_bits_tail; // @[Router.scala 129:24]
  wire [63:0] switch_io_out_1_0_bits_payload; // @[Router.scala 129:24]
  wire [1:0] switch_io_out_1_0_bits_flow_ingress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_out_1_0_bits_flow_egress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_out_1_0_bits_virt_channel_id; // @[Router.scala 129:24]
  wire  switch_io_out_0_0_valid; // @[Router.scala 129:24]
  wire  switch_io_out_0_0_bits_head; // @[Router.scala 129:24]
  wire  switch_io_out_0_0_bits_tail; // @[Router.scala 129:24]
  wire [63:0] switch_io_out_0_0_bits_payload; // @[Router.scala 129:24]
  wire [1:0] switch_io_out_0_0_bits_flow_ingress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_out_0_0_bits_flow_egress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_out_0_0_bits_virt_channel_id; // @[Router.scala 129:24]
  wire  switch_io_sel_2_0_2_0; // @[Router.scala 129:24]
  wire  switch_io_sel_2_0_1_0; // @[Router.scala 129:24]
  wire  switch_io_sel_2_0_0_0; // @[Router.scala 129:24]
  wire  switch_io_sel_1_0_2_0; // @[Router.scala 129:24]
  wire  switch_io_sel_1_0_1_0; // @[Router.scala 129:24]
  wire  switch_io_sel_1_0_0_0; // @[Router.scala 129:24]
  wire  switch_io_sel_0_0_2_0; // @[Router.scala 129:24]
  wire  switch_io_sel_0_0_1_0; // @[Router.scala 129:24]
  wire  switch_io_sel_0_0_0_0; // @[Router.scala 129:24]
  wire  switch_allocator_clock; // @[Router.scala 130:34]
  wire  switch_allocator_reset; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_ready; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_valid; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_bits_vc_sel_2_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_bits_vc_sel_1_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_bits_vc_sel_1_1; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_bits_vc_sel_1_2; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_bits_vc_sel_1_3; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_bits_vc_sel_0_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_bits_vc_sel_0_1; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_bits_vc_sel_0_2; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_bits_vc_sel_0_3; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_bits_tail; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_ready; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_valid; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_vc_sel_2_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_vc_sel_1_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_vc_sel_1_1; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_vc_sel_1_2; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_vc_sel_1_3; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_vc_sel_0_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_vc_sel_0_1; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_vc_sel_0_2; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_vc_sel_0_3; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_tail; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_ready; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_valid; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_2_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_1_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_1_1; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_1_2; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_1_3; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_0_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_0_1; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_0_2; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_0_3; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_tail; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_2_0_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_2_0_tail; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_1_0_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_1_1_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_1_2_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_1_3_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_0_0_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_0_1_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_0_2_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_0_3_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_2_0_2_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_2_0_1_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_2_0_0_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_1_0_2_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_1_0_1_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_1_0_0_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_0_0_2_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_0_0_1_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_0_0_0_0; // @[Router.scala 130:34]
  wire  vc_allocator_clock; // @[Router.scala 131:30]
  wire  vc_allocator_reset; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_ready; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_valid; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_bits_vc_sel_2_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_bits_vc_sel_1_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_bits_vc_sel_1_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_bits_vc_sel_1_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_bits_vc_sel_1_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_bits_vc_sel_0_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_bits_vc_sel_0_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_bits_vc_sel_0_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_bits_vc_sel_0_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_ready; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_valid; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_bits_vc_sel_2_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_bits_vc_sel_1_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_bits_vc_sel_1_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_bits_vc_sel_1_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_bits_vc_sel_1_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_bits_vc_sel_0_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_bits_vc_sel_0_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_bits_vc_sel_0_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_bits_vc_sel_0_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_ready; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_valid; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_2_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_1_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_1_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_1_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_1_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_0_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_0_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_0_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_0_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_2_vc_sel_2_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_2_vc_sel_1_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_2_vc_sel_1_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_2_vc_sel_1_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_2_vc_sel_1_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_2_vc_sel_0_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_2_vc_sel_0_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_2_vc_sel_0_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_2_vc_sel_0_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_1_vc_sel_2_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_1_vc_sel_1_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_1_vc_sel_1_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_1_vc_sel_1_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_1_vc_sel_1_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_1_vc_sel_0_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_1_vc_sel_0_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_1_vc_sel_0_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_1_vc_sel_0_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_2_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_1_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_1_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_1_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_1_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_0_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_0_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_0_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_0_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_2_0_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_1_0_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_1_1_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_1_2_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_1_3_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_0_0_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_0_1_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_0_2_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_0_3_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_2_0_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_1_0_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_1_1_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_1_2_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_1_3_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_0_0_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_0_1_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_0_2_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_0_3_alloc; // @[Router.scala 131:30]
  wire [1:0] route_computer_io_req_2_bits_flow_ingress_node; // @[Router.scala 134:32]
  wire [1:0] route_computer_io_req_2_bits_flow_egress_node; // @[Router.scala 134:32]
  wire [1:0] route_computer_io_req_1_bits_src_virt_id; // @[Router.scala 134:32]
  wire [1:0] route_computer_io_req_1_bits_flow_ingress_node; // @[Router.scala 134:32]
  wire [1:0] route_computer_io_req_1_bits_flow_egress_node; // @[Router.scala 134:32]
  wire [1:0] route_computer_io_req_0_bits_src_virt_id; // @[Router.scala 134:32]
  wire [1:0] route_computer_io_req_0_bits_flow_ingress_node; // @[Router.scala 134:32]
  wire [1:0] route_computer_io_req_0_bits_flow_egress_node; // @[Router.scala 134:32]
  wire  route_computer_io_resp_2_vc_sel_1_0; // @[Router.scala 134:32]
  wire  route_computer_io_resp_2_vc_sel_1_1; // @[Router.scala 134:32]
  wire  route_computer_io_resp_2_vc_sel_1_2; // @[Router.scala 134:32]
  wire  route_computer_io_resp_2_vc_sel_1_3; // @[Router.scala 134:32]
  wire  route_computer_io_resp_2_vc_sel_0_0; // @[Router.scala 134:32]
  wire  route_computer_io_resp_2_vc_sel_0_1; // @[Router.scala 134:32]
  wire  route_computer_io_resp_2_vc_sel_0_2; // @[Router.scala 134:32]
  wire  route_computer_io_resp_2_vc_sel_0_3; // @[Router.scala 134:32]
  wire  route_computer_io_resp_1_vc_sel_1_0; // @[Router.scala 134:32]
  wire  route_computer_io_resp_1_vc_sel_1_1; // @[Router.scala 134:32]
  wire  route_computer_io_resp_1_vc_sel_1_2; // @[Router.scala 134:32]
  wire  route_computer_io_resp_1_vc_sel_1_3; // @[Router.scala 134:32]
  wire  route_computer_io_resp_1_vc_sel_0_0; // @[Router.scala 134:32]
  wire  route_computer_io_resp_1_vc_sel_0_1; // @[Router.scala 134:32]
  wire  route_computer_io_resp_1_vc_sel_0_2; // @[Router.scala 134:32]
  wire  route_computer_io_resp_1_vc_sel_0_3; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_1_0; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_1_1; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_1_2; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_1_3; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_0_0; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_0_1; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_0_2; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_0_3; // @[Router.scala 134:32]
  wire [19:0] plusarg_reader_out; // @[PlusArg.scala 80:11]
  wire  _fires_count_T = vc_allocator_io_req_0_ready & vc_allocator_io_req_0_valid; // @[Decoupled.scala 51:35]
  wire  _fires_count_T_1 = vc_allocator_io_req_1_ready & vc_allocator_io_req_1_valid; // @[Decoupled.scala 51:35]
  wire  _fires_count_T_2 = vc_allocator_io_req_2_ready & vc_allocator_io_req_2_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _fires_count_T_3 = _fires_count_T_1 + _fires_count_T_2; // @[Bitwise.scala 51:90]
  wire [1:0] _GEN_5 = {{1'd0}, _fires_count_T}; // @[Bitwise.scala 51:90]
  wire [2:0] _fires_count_T_5 = _GEN_5 + _fires_count_T_3; // @[Bitwise.scala 51:90]
  reg  switch_io_sel_REG_2_0_2_0; // @[Router.scala 176:14]
  reg  switch_io_sel_REG_2_0_1_0; // @[Router.scala 176:14]
  reg  switch_io_sel_REG_2_0_0_0; // @[Router.scala 176:14]
  reg  switch_io_sel_REG_1_0_2_0; // @[Router.scala 176:14]
  reg  switch_io_sel_REG_1_0_1_0; // @[Router.scala 176:14]
  reg  switch_io_sel_REG_1_0_0_0; // @[Router.scala 176:14]
  reg  switch_io_sel_REG_0_0_2_0; // @[Router.scala 176:14]
  reg  switch_io_sel_REG_0_0_1_0; // @[Router.scala 176:14]
  reg  switch_io_sel_REG_0_0_0_0; // @[Router.scala 176:14]
  reg [63:0] debug_tsc; // @[Router.scala 193:28]
  wire [63:0] _debug_tsc_T_1 = debug_tsc + 64'h1; // @[Router.scala 194:28]
  reg [63:0] debug_sample; // @[Router.scala 195:31]
  wire [63:0] _debug_sample_T_1 = debug_sample + 64'h1; // @[Router.scala 196:34]
  wire [19:0] _T_1 = plusarg_reader_out - 20'h1; // @[Router.scala 198:40]
  wire [63:0] _GEN_6 = {{44'd0}, _T_1}; // @[Router.scala 198:24]
  wire  _T_2 = debug_sample == _GEN_6; // @[Router.scala 198:24]
  reg [63:0] util_ctr; // @[Router.scala 201:29]
  reg  fired; // @[Router.scala 202:26]
  wire [63:0] _GEN_7 = {{63'd0}, auto_dest_nodes_in_0_flit_0_valid}; // @[Router.scala 203:28]
  wire [63:0] _util_ctr_T_1 = util_ctr + _GEN_7; // @[Router.scala 203:28]
  wire  _T_8 = plusarg_reader_out != 20'h0 & _T_2 & fired; // @[Router.scala 205:71]
  reg [63:0] util_ctr_1; // @[Router.scala 201:29]
  reg  fired_1; // @[Router.scala 202:26]
  wire [63:0] _GEN_9 = {{63'd0}, auto_dest_nodes_in_1_flit_0_valid}; // @[Router.scala 203:28]
  wire [63:0] _util_ctr_T_3 = util_ctr_1 + _GEN_9; // @[Router.scala 203:28]
  wire  _T_16 = plusarg_reader_out != 20'h0 & _T_2 & fired_1; // @[Router.scala 205:71]
  wire  bundleIn_0_2_flit_ready = ingress_unit_2_from_2_io_in_ready; // @[Nodes.scala 1215:84 Router.scala 142:68]
  wire  _T_19 = bundleIn_0_2_flit_ready & auto_ingress_nodes_in_flit_valid; // @[Decoupled.scala 51:35]
  reg [63:0] util_ctr_2; // @[Router.scala 201:29]
  reg  fired_2; // @[Router.scala 202:26]
  wire [63:0] _GEN_11 = {{63'd0}, _T_19}; // @[Router.scala 203:28]
  wire [63:0] _util_ctr_T_5 = util_ctr_2 + _GEN_11; // @[Router.scala 203:28]
  wire  _T_25 = plusarg_reader_out != 20'h0 & _T_2 & fired_2; // @[Router.scala 205:71]
  wire  x1_2_flit_valid = egress_unit_2_to_2_io_out_valid; // @[Nodes.scala 1212:84 Router.scala 144:65]
  reg [63:0] util_ctr_3; // @[Router.scala 201:29]
  reg  fired_3; // @[Router.scala 202:26]
  wire [63:0] _GEN_13 = {{63'd0}, x1_2_flit_valid}; // @[Router.scala 203:28]
  wire [63:0] _util_ctr_T_7 = util_ctr_3 + _GEN_13; // @[Router.scala 203:28]
  wire  _T_34 = plusarg_reader_out != 20'h0 & _T_2 & fired_3; // @[Router.scala 205:71]
  wire [1:0] fires_count = _fires_count_T_5[1:0]; // @[Bitwise.scala 51:90]
  NoCMonitor_4 monitor ( // @[Nodes.scala 24:25]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_flit_0_valid(monitor_io_in_flit_0_valid),
    .io_in_flit_0_bits_head(monitor_io_in_flit_0_bits_head),
    .io_in_flit_0_bits_tail(monitor_io_in_flit_0_bits_tail),
    .io_in_flit_0_bits_flow_ingress_node(monitor_io_in_flit_0_bits_flow_ingress_node),
    .io_in_flit_0_bits_flow_egress_node(monitor_io_in_flit_0_bits_flow_egress_node),
    .io_in_flit_0_bits_virt_channel_id(monitor_io_in_flit_0_bits_virt_channel_id)
  );
  NoCMonitor_5 monitor_1 ( // @[Nodes.scala 24:25]
    .clock(monitor_1_clock),
    .reset(monitor_1_reset),
    .io_in_flit_0_valid(monitor_1_io_in_flit_0_valid),
    .io_in_flit_0_bits_head(monitor_1_io_in_flit_0_bits_head),
    .io_in_flit_0_bits_tail(monitor_1_io_in_flit_0_bits_tail),
    .io_in_flit_0_bits_flow_ingress_node(monitor_1_io_in_flit_0_bits_flow_ingress_node),
    .io_in_flit_0_bits_flow_egress_node(monitor_1_io_in_flit_0_bits_flow_egress_node),
    .io_in_flit_0_bits_virt_channel_id(monitor_1_io_in_flit_0_bits_virt_channel_id)
  );
  InputUnit_4 input_unit_0_from_1 ( // @[Router.scala 112:13]
    .clock(input_unit_0_from_1_clock),
    .reset(input_unit_0_from_1_reset),
    .io_router_req_valid(input_unit_0_from_1_io_router_req_valid),
    .io_router_req_bits_src_virt_id(input_unit_0_from_1_io_router_req_bits_src_virt_id),
    .io_router_req_bits_flow_ingress_node(input_unit_0_from_1_io_router_req_bits_flow_ingress_node),
    .io_router_req_bits_flow_egress_node(input_unit_0_from_1_io_router_req_bits_flow_egress_node),
    .io_router_resp_vc_sel_1_0(input_unit_0_from_1_io_router_resp_vc_sel_1_0),
    .io_router_resp_vc_sel_1_1(input_unit_0_from_1_io_router_resp_vc_sel_1_1),
    .io_router_resp_vc_sel_1_2(input_unit_0_from_1_io_router_resp_vc_sel_1_2),
    .io_router_resp_vc_sel_1_3(input_unit_0_from_1_io_router_resp_vc_sel_1_3),
    .io_router_resp_vc_sel_0_0(input_unit_0_from_1_io_router_resp_vc_sel_0_0),
    .io_router_resp_vc_sel_0_1(input_unit_0_from_1_io_router_resp_vc_sel_0_1),
    .io_router_resp_vc_sel_0_2(input_unit_0_from_1_io_router_resp_vc_sel_0_2),
    .io_router_resp_vc_sel_0_3(input_unit_0_from_1_io_router_resp_vc_sel_0_3),
    .io_vcalloc_req_ready(input_unit_0_from_1_io_vcalloc_req_ready),
    .io_vcalloc_req_valid(input_unit_0_from_1_io_vcalloc_req_valid),
    .io_vcalloc_req_bits_vc_sel_2_0(input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_2_0),
    .io_vcalloc_req_bits_vc_sel_1_0(input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_1_0),
    .io_vcalloc_req_bits_vc_sel_1_1(input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_1_1),
    .io_vcalloc_req_bits_vc_sel_1_2(input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_1_2),
    .io_vcalloc_req_bits_vc_sel_1_3(input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_1_3),
    .io_vcalloc_req_bits_vc_sel_0_0(input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_0_0),
    .io_vcalloc_req_bits_vc_sel_0_1(input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_0_1),
    .io_vcalloc_req_bits_vc_sel_0_2(input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_0_2),
    .io_vcalloc_req_bits_vc_sel_0_3(input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_0_3),
    .io_vcalloc_resp_vc_sel_2_0(input_unit_0_from_1_io_vcalloc_resp_vc_sel_2_0),
    .io_vcalloc_resp_vc_sel_1_0(input_unit_0_from_1_io_vcalloc_resp_vc_sel_1_0),
    .io_vcalloc_resp_vc_sel_1_1(input_unit_0_from_1_io_vcalloc_resp_vc_sel_1_1),
    .io_vcalloc_resp_vc_sel_1_2(input_unit_0_from_1_io_vcalloc_resp_vc_sel_1_2),
    .io_vcalloc_resp_vc_sel_1_3(input_unit_0_from_1_io_vcalloc_resp_vc_sel_1_3),
    .io_vcalloc_resp_vc_sel_0_0(input_unit_0_from_1_io_vcalloc_resp_vc_sel_0_0),
    .io_vcalloc_resp_vc_sel_0_1(input_unit_0_from_1_io_vcalloc_resp_vc_sel_0_1),
    .io_vcalloc_resp_vc_sel_0_2(input_unit_0_from_1_io_vcalloc_resp_vc_sel_0_2),
    .io_vcalloc_resp_vc_sel_0_3(input_unit_0_from_1_io_vcalloc_resp_vc_sel_0_3),
    .io_out_credit_available_2_0(input_unit_0_from_1_io_out_credit_available_2_0),
    .io_out_credit_available_1_0(input_unit_0_from_1_io_out_credit_available_1_0),
    .io_out_credit_available_1_1(input_unit_0_from_1_io_out_credit_available_1_1),
    .io_out_credit_available_1_2(input_unit_0_from_1_io_out_credit_available_1_2),
    .io_out_credit_available_1_3(input_unit_0_from_1_io_out_credit_available_1_3),
    .io_out_credit_available_0_0(input_unit_0_from_1_io_out_credit_available_0_0),
    .io_out_credit_available_0_1(input_unit_0_from_1_io_out_credit_available_0_1),
    .io_out_credit_available_0_2(input_unit_0_from_1_io_out_credit_available_0_2),
    .io_out_credit_available_0_3(input_unit_0_from_1_io_out_credit_available_0_3),
    .io_salloc_req_0_ready(input_unit_0_from_1_io_salloc_req_0_ready),
    .io_salloc_req_0_valid(input_unit_0_from_1_io_salloc_req_0_valid),
    .io_salloc_req_0_bits_vc_sel_2_0(input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_2_0),
    .io_salloc_req_0_bits_vc_sel_1_0(input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_1_0),
    .io_salloc_req_0_bits_vc_sel_1_1(input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_1_1),
    .io_salloc_req_0_bits_vc_sel_1_2(input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_1_2),
    .io_salloc_req_0_bits_vc_sel_1_3(input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_1_3),
    .io_salloc_req_0_bits_vc_sel_0_0(input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_0_0),
    .io_salloc_req_0_bits_vc_sel_0_1(input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_0_1),
    .io_salloc_req_0_bits_vc_sel_0_2(input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_0_2),
    .io_salloc_req_0_bits_vc_sel_0_3(input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_0_3),
    .io_salloc_req_0_bits_tail(input_unit_0_from_1_io_salloc_req_0_bits_tail),
    .io_out_0_valid(input_unit_0_from_1_io_out_0_valid),
    .io_out_0_bits_flit_head(input_unit_0_from_1_io_out_0_bits_flit_head),
    .io_out_0_bits_flit_tail(input_unit_0_from_1_io_out_0_bits_flit_tail),
    .io_out_0_bits_flit_payload(input_unit_0_from_1_io_out_0_bits_flit_payload),
    .io_out_0_bits_flit_flow_ingress_node(input_unit_0_from_1_io_out_0_bits_flit_flow_ingress_node),
    .io_out_0_bits_flit_flow_egress_node(input_unit_0_from_1_io_out_0_bits_flit_flow_egress_node),
    .io_out_0_bits_out_virt_channel(input_unit_0_from_1_io_out_0_bits_out_virt_channel),
    .io_debug_va_stall(input_unit_0_from_1_io_debug_va_stall),
    .io_debug_sa_stall(input_unit_0_from_1_io_debug_sa_stall),
    .io_in_flit_0_valid(input_unit_0_from_1_io_in_flit_0_valid),
    .io_in_flit_0_bits_head(input_unit_0_from_1_io_in_flit_0_bits_head),
    .io_in_flit_0_bits_tail(input_unit_0_from_1_io_in_flit_0_bits_tail),
    .io_in_flit_0_bits_payload(input_unit_0_from_1_io_in_flit_0_bits_payload),
    .io_in_flit_0_bits_flow_ingress_node(input_unit_0_from_1_io_in_flit_0_bits_flow_ingress_node),
    .io_in_flit_0_bits_flow_egress_node(input_unit_0_from_1_io_in_flit_0_bits_flow_egress_node),
    .io_in_flit_0_bits_virt_channel_id(input_unit_0_from_1_io_in_flit_0_bits_virt_channel_id),
    .io_in_credit_return(input_unit_0_from_1_io_in_credit_return),
    .io_in_vc_free(input_unit_0_from_1_io_in_vc_free)
  );
  InputUnit_5 input_unit_1_from_3 ( // @[Router.scala 112:13]
    .clock(input_unit_1_from_3_clock),
    .reset(input_unit_1_from_3_reset),
    .io_router_req_valid(input_unit_1_from_3_io_router_req_valid),
    .io_router_req_bits_src_virt_id(input_unit_1_from_3_io_router_req_bits_src_virt_id),
    .io_router_req_bits_flow_ingress_node(input_unit_1_from_3_io_router_req_bits_flow_ingress_node),
    .io_router_req_bits_flow_egress_node(input_unit_1_from_3_io_router_req_bits_flow_egress_node),
    .io_router_resp_vc_sel_1_0(input_unit_1_from_3_io_router_resp_vc_sel_1_0),
    .io_router_resp_vc_sel_1_1(input_unit_1_from_3_io_router_resp_vc_sel_1_1),
    .io_router_resp_vc_sel_1_2(input_unit_1_from_3_io_router_resp_vc_sel_1_2),
    .io_router_resp_vc_sel_1_3(input_unit_1_from_3_io_router_resp_vc_sel_1_3),
    .io_router_resp_vc_sel_0_0(input_unit_1_from_3_io_router_resp_vc_sel_0_0),
    .io_router_resp_vc_sel_0_1(input_unit_1_from_3_io_router_resp_vc_sel_0_1),
    .io_router_resp_vc_sel_0_2(input_unit_1_from_3_io_router_resp_vc_sel_0_2),
    .io_router_resp_vc_sel_0_3(input_unit_1_from_3_io_router_resp_vc_sel_0_3),
    .io_vcalloc_req_ready(input_unit_1_from_3_io_vcalloc_req_ready),
    .io_vcalloc_req_valid(input_unit_1_from_3_io_vcalloc_req_valid),
    .io_vcalloc_req_bits_vc_sel_2_0(input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_2_0),
    .io_vcalloc_req_bits_vc_sel_1_0(input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_1_0),
    .io_vcalloc_req_bits_vc_sel_1_1(input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_1_1),
    .io_vcalloc_req_bits_vc_sel_1_2(input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_1_2),
    .io_vcalloc_req_bits_vc_sel_1_3(input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_1_3),
    .io_vcalloc_req_bits_vc_sel_0_0(input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_0_0),
    .io_vcalloc_req_bits_vc_sel_0_1(input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_0_1),
    .io_vcalloc_req_bits_vc_sel_0_2(input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_0_2),
    .io_vcalloc_req_bits_vc_sel_0_3(input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_0_3),
    .io_vcalloc_resp_vc_sel_2_0(input_unit_1_from_3_io_vcalloc_resp_vc_sel_2_0),
    .io_vcalloc_resp_vc_sel_1_0(input_unit_1_from_3_io_vcalloc_resp_vc_sel_1_0),
    .io_vcalloc_resp_vc_sel_1_1(input_unit_1_from_3_io_vcalloc_resp_vc_sel_1_1),
    .io_vcalloc_resp_vc_sel_1_2(input_unit_1_from_3_io_vcalloc_resp_vc_sel_1_2),
    .io_vcalloc_resp_vc_sel_1_3(input_unit_1_from_3_io_vcalloc_resp_vc_sel_1_3),
    .io_vcalloc_resp_vc_sel_0_0(input_unit_1_from_3_io_vcalloc_resp_vc_sel_0_0),
    .io_vcalloc_resp_vc_sel_0_1(input_unit_1_from_3_io_vcalloc_resp_vc_sel_0_1),
    .io_vcalloc_resp_vc_sel_0_2(input_unit_1_from_3_io_vcalloc_resp_vc_sel_0_2),
    .io_vcalloc_resp_vc_sel_0_3(input_unit_1_from_3_io_vcalloc_resp_vc_sel_0_3),
    .io_out_credit_available_2_0(input_unit_1_from_3_io_out_credit_available_2_0),
    .io_out_credit_available_1_0(input_unit_1_from_3_io_out_credit_available_1_0),
    .io_out_credit_available_1_1(input_unit_1_from_3_io_out_credit_available_1_1),
    .io_out_credit_available_1_2(input_unit_1_from_3_io_out_credit_available_1_2),
    .io_out_credit_available_1_3(input_unit_1_from_3_io_out_credit_available_1_3),
    .io_out_credit_available_0_0(input_unit_1_from_3_io_out_credit_available_0_0),
    .io_out_credit_available_0_1(input_unit_1_from_3_io_out_credit_available_0_1),
    .io_out_credit_available_0_2(input_unit_1_from_3_io_out_credit_available_0_2),
    .io_out_credit_available_0_3(input_unit_1_from_3_io_out_credit_available_0_3),
    .io_salloc_req_0_ready(input_unit_1_from_3_io_salloc_req_0_ready),
    .io_salloc_req_0_valid(input_unit_1_from_3_io_salloc_req_0_valid),
    .io_salloc_req_0_bits_vc_sel_2_0(input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_2_0),
    .io_salloc_req_0_bits_vc_sel_1_0(input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_1_0),
    .io_salloc_req_0_bits_vc_sel_1_1(input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_1_1),
    .io_salloc_req_0_bits_vc_sel_1_2(input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_1_2),
    .io_salloc_req_0_bits_vc_sel_1_3(input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_1_3),
    .io_salloc_req_0_bits_vc_sel_0_0(input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_0_0),
    .io_salloc_req_0_bits_vc_sel_0_1(input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_0_1),
    .io_salloc_req_0_bits_vc_sel_0_2(input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_0_2),
    .io_salloc_req_0_bits_vc_sel_0_3(input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_0_3),
    .io_salloc_req_0_bits_tail(input_unit_1_from_3_io_salloc_req_0_bits_tail),
    .io_out_0_valid(input_unit_1_from_3_io_out_0_valid),
    .io_out_0_bits_flit_head(input_unit_1_from_3_io_out_0_bits_flit_head),
    .io_out_0_bits_flit_tail(input_unit_1_from_3_io_out_0_bits_flit_tail),
    .io_out_0_bits_flit_payload(input_unit_1_from_3_io_out_0_bits_flit_payload),
    .io_out_0_bits_flit_flow_ingress_node(input_unit_1_from_3_io_out_0_bits_flit_flow_ingress_node),
    .io_out_0_bits_flit_flow_egress_node(input_unit_1_from_3_io_out_0_bits_flit_flow_egress_node),
    .io_out_0_bits_out_virt_channel(input_unit_1_from_3_io_out_0_bits_out_virt_channel),
    .io_debug_va_stall(input_unit_1_from_3_io_debug_va_stall),
    .io_debug_sa_stall(input_unit_1_from_3_io_debug_sa_stall),
    .io_in_flit_0_valid(input_unit_1_from_3_io_in_flit_0_valid),
    .io_in_flit_0_bits_head(input_unit_1_from_3_io_in_flit_0_bits_head),
    .io_in_flit_0_bits_tail(input_unit_1_from_3_io_in_flit_0_bits_tail),
    .io_in_flit_0_bits_payload(input_unit_1_from_3_io_in_flit_0_bits_payload),
    .io_in_flit_0_bits_flow_ingress_node(input_unit_1_from_3_io_in_flit_0_bits_flow_ingress_node),
    .io_in_flit_0_bits_flow_egress_node(input_unit_1_from_3_io_in_flit_0_bits_flow_egress_node),
    .io_in_flit_0_bits_virt_channel_id(input_unit_1_from_3_io_in_flit_0_bits_virt_channel_id),
    .io_in_credit_return(input_unit_1_from_3_io_in_credit_return),
    .io_in_vc_free(input_unit_1_from_3_io_in_vc_free)
  );
  IngressUnit_2 ingress_unit_2_from_2 ( // @[Router.scala 116:13]
    .clock(ingress_unit_2_from_2_clock),
    .reset(ingress_unit_2_from_2_reset),
    .io_router_req_valid(ingress_unit_2_from_2_io_router_req_valid),
    .io_router_req_bits_flow_ingress_node(ingress_unit_2_from_2_io_router_req_bits_flow_ingress_node),
    .io_router_req_bits_flow_egress_node(ingress_unit_2_from_2_io_router_req_bits_flow_egress_node),
    .io_router_resp_vc_sel_1_0(ingress_unit_2_from_2_io_router_resp_vc_sel_1_0),
    .io_router_resp_vc_sel_1_1(ingress_unit_2_from_2_io_router_resp_vc_sel_1_1),
    .io_router_resp_vc_sel_1_2(ingress_unit_2_from_2_io_router_resp_vc_sel_1_2),
    .io_router_resp_vc_sel_1_3(ingress_unit_2_from_2_io_router_resp_vc_sel_1_3),
    .io_router_resp_vc_sel_0_0(ingress_unit_2_from_2_io_router_resp_vc_sel_0_0),
    .io_router_resp_vc_sel_0_1(ingress_unit_2_from_2_io_router_resp_vc_sel_0_1),
    .io_router_resp_vc_sel_0_2(ingress_unit_2_from_2_io_router_resp_vc_sel_0_2),
    .io_router_resp_vc_sel_0_3(ingress_unit_2_from_2_io_router_resp_vc_sel_0_3),
    .io_vcalloc_req_ready(ingress_unit_2_from_2_io_vcalloc_req_ready),
    .io_vcalloc_req_valid(ingress_unit_2_from_2_io_vcalloc_req_valid),
    .io_vcalloc_req_bits_vc_sel_2_0(ingress_unit_2_from_2_io_vcalloc_req_bits_vc_sel_2_0),
    .io_vcalloc_req_bits_vc_sel_1_0(ingress_unit_2_from_2_io_vcalloc_req_bits_vc_sel_1_0),
    .io_vcalloc_req_bits_vc_sel_1_1(ingress_unit_2_from_2_io_vcalloc_req_bits_vc_sel_1_1),
    .io_vcalloc_req_bits_vc_sel_1_2(ingress_unit_2_from_2_io_vcalloc_req_bits_vc_sel_1_2),
    .io_vcalloc_req_bits_vc_sel_1_3(ingress_unit_2_from_2_io_vcalloc_req_bits_vc_sel_1_3),
    .io_vcalloc_req_bits_vc_sel_0_0(ingress_unit_2_from_2_io_vcalloc_req_bits_vc_sel_0_0),
    .io_vcalloc_req_bits_vc_sel_0_1(ingress_unit_2_from_2_io_vcalloc_req_bits_vc_sel_0_1),
    .io_vcalloc_req_bits_vc_sel_0_2(ingress_unit_2_from_2_io_vcalloc_req_bits_vc_sel_0_2),
    .io_vcalloc_req_bits_vc_sel_0_3(ingress_unit_2_from_2_io_vcalloc_req_bits_vc_sel_0_3),
    .io_vcalloc_resp_vc_sel_2_0(ingress_unit_2_from_2_io_vcalloc_resp_vc_sel_2_0),
    .io_vcalloc_resp_vc_sel_1_0(ingress_unit_2_from_2_io_vcalloc_resp_vc_sel_1_0),
    .io_vcalloc_resp_vc_sel_1_1(ingress_unit_2_from_2_io_vcalloc_resp_vc_sel_1_1),
    .io_vcalloc_resp_vc_sel_1_2(ingress_unit_2_from_2_io_vcalloc_resp_vc_sel_1_2),
    .io_vcalloc_resp_vc_sel_1_3(ingress_unit_2_from_2_io_vcalloc_resp_vc_sel_1_3),
    .io_vcalloc_resp_vc_sel_0_0(ingress_unit_2_from_2_io_vcalloc_resp_vc_sel_0_0),
    .io_vcalloc_resp_vc_sel_0_1(ingress_unit_2_from_2_io_vcalloc_resp_vc_sel_0_1),
    .io_vcalloc_resp_vc_sel_0_2(ingress_unit_2_from_2_io_vcalloc_resp_vc_sel_0_2),
    .io_vcalloc_resp_vc_sel_0_3(ingress_unit_2_from_2_io_vcalloc_resp_vc_sel_0_3),
    .io_out_credit_available_2_0(ingress_unit_2_from_2_io_out_credit_available_2_0),
    .io_out_credit_available_1_0(ingress_unit_2_from_2_io_out_credit_available_1_0),
    .io_out_credit_available_1_1(ingress_unit_2_from_2_io_out_credit_available_1_1),
    .io_out_credit_available_1_2(ingress_unit_2_from_2_io_out_credit_available_1_2),
    .io_out_credit_available_1_3(ingress_unit_2_from_2_io_out_credit_available_1_3),
    .io_out_credit_available_0_0(ingress_unit_2_from_2_io_out_credit_available_0_0),
    .io_out_credit_available_0_1(ingress_unit_2_from_2_io_out_credit_available_0_1),
    .io_out_credit_available_0_2(ingress_unit_2_from_2_io_out_credit_available_0_2),
    .io_out_credit_available_0_3(ingress_unit_2_from_2_io_out_credit_available_0_3),
    .io_salloc_req_0_ready(ingress_unit_2_from_2_io_salloc_req_0_ready),
    .io_salloc_req_0_valid(ingress_unit_2_from_2_io_salloc_req_0_valid),
    .io_salloc_req_0_bits_vc_sel_2_0(ingress_unit_2_from_2_io_salloc_req_0_bits_vc_sel_2_0),
    .io_salloc_req_0_bits_vc_sel_1_0(ingress_unit_2_from_2_io_salloc_req_0_bits_vc_sel_1_0),
    .io_salloc_req_0_bits_vc_sel_1_1(ingress_unit_2_from_2_io_salloc_req_0_bits_vc_sel_1_1),
    .io_salloc_req_0_bits_vc_sel_1_2(ingress_unit_2_from_2_io_salloc_req_0_bits_vc_sel_1_2),
    .io_salloc_req_0_bits_vc_sel_1_3(ingress_unit_2_from_2_io_salloc_req_0_bits_vc_sel_1_3),
    .io_salloc_req_0_bits_vc_sel_0_0(ingress_unit_2_from_2_io_salloc_req_0_bits_vc_sel_0_0),
    .io_salloc_req_0_bits_vc_sel_0_1(ingress_unit_2_from_2_io_salloc_req_0_bits_vc_sel_0_1),
    .io_salloc_req_0_bits_vc_sel_0_2(ingress_unit_2_from_2_io_salloc_req_0_bits_vc_sel_0_2),
    .io_salloc_req_0_bits_vc_sel_0_3(ingress_unit_2_from_2_io_salloc_req_0_bits_vc_sel_0_3),
    .io_salloc_req_0_bits_tail(ingress_unit_2_from_2_io_salloc_req_0_bits_tail),
    .io_out_0_valid(ingress_unit_2_from_2_io_out_0_valid),
    .io_out_0_bits_flit_head(ingress_unit_2_from_2_io_out_0_bits_flit_head),
    .io_out_0_bits_flit_tail(ingress_unit_2_from_2_io_out_0_bits_flit_tail),
    .io_out_0_bits_flit_payload(ingress_unit_2_from_2_io_out_0_bits_flit_payload),
    .io_out_0_bits_flit_flow_ingress_node(ingress_unit_2_from_2_io_out_0_bits_flit_flow_ingress_node),
    .io_out_0_bits_flit_flow_egress_node(ingress_unit_2_from_2_io_out_0_bits_flit_flow_egress_node),
    .io_out_0_bits_out_virt_channel(ingress_unit_2_from_2_io_out_0_bits_out_virt_channel),
    .io_in_ready(ingress_unit_2_from_2_io_in_ready),
    .io_in_valid(ingress_unit_2_from_2_io_in_valid),
    .io_in_bits_head(ingress_unit_2_from_2_io_in_bits_head),
    .io_in_bits_tail(ingress_unit_2_from_2_io_in_bits_tail),
    .io_in_bits_payload(ingress_unit_2_from_2_io_in_bits_payload),
    .io_in_bits_egress_id(ingress_unit_2_from_2_io_in_bits_egress_id)
  );
  OutputUnit output_unit_0_to_1 ( // @[Router.scala 122:13]
    .clock(output_unit_0_to_1_clock),
    .reset(output_unit_0_to_1_reset),
    .io_in_0_valid(output_unit_0_to_1_io_in_0_valid),
    .io_in_0_bits_head(output_unit_0_to_1_io_in_0_bits_head),
    .io_in_0_bits_tail(output_unit_0_to_1_io_in_0_bits_tail),
    .io_in_0_bits_payload(output_unit_0_to_1_io_in_0_bits_payload),
    .io_in_0_bits_flow_ingress_node(output_unit_0_to_1_io_in_0_bits_flow_ingress_node),
    .io_in_0_bits_flow_egress_node(output_unit_0_to_1_io_in_0_bits_flow_egress_node),
    .io_in_0_bits_virt_channel_id(output_unit_0_to_1_io_in_0_bits_virt_channel_id),
    .io_credit_available_0(output_unit_0_to_1_io_credit_available_0),
    .io_credit_available_1(output_unit_0_to_1_io_credit_available_1),
    .io_credit_available_2(output_unit_0_to_1_io_credit_available_2),
    .io_credit_available_3(output_unit_0_to_1_io_credit_available_3),
    .io_channel_status_0_occupied(output_unit_0_to_1_io_channel_status_0_occupied),
    .io_channel_status_1_occupied(output_unit_0_to_1_io_channel_status_1_occupied),
    .io_channel_status_2_occupied(output_unit_0_to_1_io_channel_status_2_occupied),
    .io_channel_status_3_occupied(output_unit_0_to_1_io_channel_status_3_occupied),
    .io_allocs_0_alloc(output_unit_0_to_1_io_allocs_0_alloc),
    .io_allocs_1_alloc(output_unit_0_to_1_io_allocs_1_alloc),
    .io_allocs_2_alloc(output_unit_0_to_1_io_allocs_2_alloc),
    .io_allocs_3_alloc(output_unit_0_to_1_io_allocs_3_alloc),
    .io_credit_alloc_0_alloc(output_unit_0_to_1_io_credit_alloc_0_alloc),
    .io_credit_alloc_1_alloc(output_unit_0_to_1_io_credit_alloc_1_alloc),
    .io_credit_alloc_2_alloc(output_unit_0_to_1_io_credit_alloc_2_alloc),
    .io_credit_alloc_3_alloc(output_unit_0_to_1_io_credit_alloc_3_alloc),
    .io_out_flit_0_valid(output_unit_0_to_1_io_out_flit_0_valid),
    .io_out_flit_0_bits_head(output_unit_0_to_1_io_out_flit_0_bits_head),
    .io_out_flit_0_bits_tail(output_unit_0_to_1_io_out_flit_0_bits_tail),
    .io_out_flit_0_bits_payload(output_unit_0_to_1_io_out_flit_0_bits_payload),
    .io_out_flit_0_bits_flow_ingress_node(output_unit_0_to_1_io_out_flit_0_bits_flow_ingress_node),
    .io_out_flit_0_bits_flow_egress_node(output_unit_0_to_1_io_out_flit_0_bits_flow_egress_node),
    .io_out_flit_0_bits_virt_channel_id(output_unit_0_to_1_io_out_flit_0_bits_virt_channel_id),
    .io_out_credit_return(output_unit_0_to_1_io_out_credit_return),
    .io_out_vc_free(output_unit_0_to_1_io_out_vc_free)
  );
  OutputUnit output_unit_1_to_3 ( // @[Router.scala 122:13]
    .clock(output_unit_1_to_3_clock),
    .reset(output_unit_1_to_3_reset),
    .io_in_0_valid(output_unit_1_to_3_io_in_0_valid),
    .io_in_0_bits_head(output_unit_1_to_3_io_in_0_bits_head),
    .io_in_0_bits_tail(output_unit_1_to_3_io_in_0_bits_tail),
    .io_in_0_bits_payload(output_unit_1_to_3_io_in_0_bits_payload),
    .io_in_0_bits_flow_ingress_node(output_unit_1_to_3_io_in_0_bits_flow_ingress_node),
    .io_in_0_bits_flow_egress_node(output_unit_1_to_3_io_in_0_bits_flow_egress_node),
    .io_in_0_bits_virt_channel_id(output_unit_1_to_3_io_in_0_bits_virt_channel_id),
    .io_credit_available_0(output_unit_1_to_3_io_credit_available_0),
    .io_credit_available_1(output_unit_1_to_3_io_credit_available_1),
    .io_credit_available_2(output_unit_1_to_3_io_credit_available_2),
    .io_credit_available_3(output_unit_1_to_3_io_credit_available_3),
    .io_channel_status_0_occupied(output_unit_1_to_3_io_channel_status_0_occupied),
    .io_channel_status_1_occupied(output_unit_1_to_3_io_channel_status_1_occupied),
    .io_channel_status_2_occupied(output_unit_1_to_3_io_channel_status_2_occupied),
    .io_channel_status_3_occupied(output_unit_1_to_3_io_channel_status_3_occupied),
    .io_allocs_0_alloc(output_unit_1_to_3_io_allocs_0_alloc),
    .io_allocs_1_alloc(output_unit_1_to_3_io_allocs_1_alloc),
    .io_allocs_2_alloc(output_unit_1_to_3_io_allocs_2_alloc),
    .io_allocs_3_alloc(output_unit_1_to_3_io_allocs_3_alloc),
    .io_credit_alloc_0_alloc(output_unit_1_to_3_io_credit_alloc_0_alloc),
    .io_credit_alloc_1_alloc(output_unit_1_to_3_io_credit_alloc_1_alloc),
    .io_credit_alloc_2_alloc(output_unit_1_to_3_io_credit_alloc_2_alloc),
    .io_credit_alloc_3_alloc(output_unit_1_to_3_io_credit_alloc_3_alloc),
    .io_out_flit_0_valid(output_unit_1_to_3_io_out_flit_0_valid),
    .io_out_flit_0_bits_head(output_unit_1_to_3_io_out_flit_0_bits_head),
    .io_out_flit_0_bits_tail(output_unit_1_to_3_io_out_flit_0_bits_tail),
    .io_out_flit_0_bits_payload(output_unit_1_to_3_io_out_flit_0_bits_payload),
    .io_out_flit_0_bits_flow_ingress_node(output_unit_1_to_3_io_out_flit_0_bits_flow_ingress_node),
    .io_out_flit_0_bits_flow_egress_node(output_unit_1_to_3_io_out_flit_0_bits_flow_egress_node),
    .io_out_flit_0_bits_virt_channel_id(output_unit_1_to_3_io_out_flit_0_bits_virt_channel_id),
    .io_out_credit_return(output_unit_1_to_3_io_out_credit_return),
    .io_out_vc_free(output_unit_1_to_3_io_out_vc_free)
  );
  EgressUnit egress_unit_2_to_2 ( // @[Router.scala 125:13]
    .clock(egress_unit_2_to_2_clock),
    .reset(egress_unit_2_to_2_reset),
    .io_in_0_valid(egress_unit_2_to_2_io_in_0_valid),
    .io_in_0_bits_head(egress_unit_2_to_2_io_in_0_bits_head),
    .io_in_0_bits_tail(egress_unit_2_to_2_io_in_0_bits_tail),
    .io_in_0_bits_payload(egress_unit_2_to_2_io_in_0_bits_payload),
    .io_in_0_bits_flow_ingress_node(egress_unit_2_to_2_io_in_0_bits_flow_ingress_node),
    .io_credit_available_0(egress_unit_2_to_2_io_credit_available_0),
    .io_channel_status_0_occupied(egress_unit_2_to_2_io_channel_status_0_occupied),
    .io_allocs_0_alloc(egress_unit_2_to_2_io_allocs_0_alloc),
    .io_credit_alloc_0_alloc(egress_unit_2_to_2_io_credit_alloc_0_alloc),
    .io_credit_alloc_0_tail(egress_unit_2_to_2_io_credit_alloc_0_tail),
    .io_out_valid(egress_unit_2_to_2_io_out_valid),
    .io_out_bits_head(egress_unit_2_to_2_io_out_bits_head),
    .io_out_bits_tail(egress_unit_2_to_2_io_out_bits_tail),
    .io_out_bits_payload(egress_unit_2_to_2_io_out_bits_payload),
    .io_out_bits_ingress_id(egress_unit_2_to_2_io_out_bits_ingress_id)
  );
  Switch switch ( // @[Router.scala 129:24]
    .clock(switch_clock),
    .reset(switch_reset),
    .io_in_2_0_valid(switch_io_in_2_0_valid),
    .io_in_2_0_bits_flit_head(switch_io_in_2_0_bits_flit_head),
    .io_in_2_0_bits_flit_tail(switch_io_in_2_0_bits_flit_tail),
    .io_in_2_0_bits_flit_payload(switch_io_in_2_0_bits_flit_payload),
    .io_in_2_0_bits_flit_flow_ingress_node(switch_io_in_2_0_bits_flit_flow_ingress_node),
    .io_in_2_0_bits_flit_flow_egress_node(switch_io_in_2_0_bits_flit_flow_egress_node),
    .io_in_2_0_bits_out_virt_channel(switch_io_in_2_0_bits_out_virt_channel),
    .io_in_1_0_valid(switch_io_in_1_0_valid),
    .io_in_1_0_bits_flit_head(switch_io_in_1_0_bits_flit_head),
    .io_in_1_0_bits_flit_tail(switch_io_in_1_0_bits_flit_tail),
    .io_in_1_0_bits_flit_payload(switch_io_in_1_0_bits_flit_payload),
    .io_in_1_0_bits_flit_flow_ingress_node(switch_io_in_1_0_bits_flit_flow_ingress_node),
    .io_in_1_0_bits_flit_flow_egress_node(switch_io_in_1_0_bits_flit_flow_egress_node),
    .io_in_1_0_bits_out_virt_channel(switch_io_in_1_0_bits_out_virt_channel),
    .io_in_0_0_valid(switch_io_in_0_0_valid),
    .io_in_0_0_bits_flit_head(switch_io_in_0_0_bits_flit_head),
    .io_in_0_0_bits_flit_tail(switch_io_in_0_0_bits_flit_tail),
    .io_in_0_0_bits_flit_payload(switch_io_in_0_0_bits_flit_payload),
    .io_in_0_0_bits_flit_flow_ingress_node(switch_io_in_0_0_bits_flit_flow_ingress_node),
    .io_in_0_0_bits_flit_flow_egress_node(switch_io_in_0_0_bits_flit_flow_egress_node),
    .io_in_0_0_bits_out_virt_channel(switch_io_in_0_0_bits_out_virt_channel),
    .io_out_2_0_valid(switch_io_out_2_0_valid),
    .io_out_2_0_bits_head(switch_io_out_2_0_bits_head),
    .io_out_2_0_bits_tail(switch_io_out_2_0_bits_tail),
    .io_out_2_0_bits_payload(switch_io_out_2_0_bits_payload),
    .io_out_2_0_bits_flow_ingress_node(switch_io_out_2_0_bits_flow_ingress_node),
    .io_out_1_0_valid(switch_io_out_1_0_valid),
    .io_out_1_0_bits_head(switch_io_out_1_0_bits_head),
    .io_out_1_0_bits_tail(switch_io_out_1_0_bits_tail),
    .io_out_1_0_bits_payload(switch_io_out_1_0_bits_payload),
    .io_out_1_0_bits_flow_ingress_node(switch_io_out_1_0_bits_flow_ingress_node),
    .io_out_1_0_bits_flow_egress_node(switch_io_out_1_0_bits_flow_egress_node),
    .io_out_1_0_bits_virt_channel_id(switch_io_out_1_0_bits_virt_channel_id),
    .io_out_0_0_valid(switch_io_out_0_0_valid),
    .io_out_0_0_bits_head(switch_io_out_0_0_bits_head),
    .io_out_0_0_bits_tail(switch_io_out_0_0_bits_tail),
    .io_out_0_0_bits_payload(switch_io_out_0_0_bits_payload),
    .io_out_0_0_bits_flow_ingress_node(switch_io_out_0_0_bits_flow_ingress_node),
    .io_out_0_0_bits_flow_egress_node(switch_io_out_0_0_bits_flow_egress_node),
    .io_out_0_0_bits_virt_channel_id(switch_io_out_0_0_bits_virt_channel_id),
    .io_sel_2_0_2_0(switch_io_sel_2_0_2_0),
    .io_sel_2_0_1_0(switch_io_sel_2_0_1_0),
    .io_sel_2_0_0_0(switch_io_sel_2_0_0_0),
    .io_sel_1_0_2_0(switch_io_sel_1_0_2_0),
    .io_sel_1_0_1_0(switch_io_sel_1_0_1_0),
    .io_sel_1_0_0_0(switch_io_sel_1_0_0_0),
    .io_sel_0_0_2_0(switch_io_sel_0_0_2_0),
    .io_sel_0_0_1_0(switch_io_sel_0_0_1_0),
    .io_sel_0_0_0_0(switch_io_sel_0_0_0_0)
  );
  SwitchAllocator switch_allocator ( // @[Router.scala 130:34]
    .clock(switch_allocator_clock),
    .reset(switch_allocator_reset),
    .io_req_2_0_ready(switch_allocator_io_req_2_0_ready),
    .io_req_2_0_valid(switch_allocator_io_req_2_0_valid),
    .io_req_2_0_bits_vc_sel_2_0(switch_allocator_io_req_2_0_bits_vc_sel_2_0),
    .io_req_2_0_bits_vc_sel_1_0(switch_allocator_io_req_2_0_bits_vc_sel_1_0),
    .io_req_2_0_bits_vc_sel_1_1(switch_allocator_io_req_2_0_bits_vc_sel_1_1),
    .io_req_2_0_bits_vc_sel_1_2(switch_allocator_io_req_2_0_bits_vc_sel_1_2),
    .io_req_2_0_bits_vc_sel_1_3(switch_allocator_io_req_2_0_bits_vc_sel_1_3),
    .io_req_2_0_bits_vc_sel_0_0(switch_allocator_io_req_2_0_bits_vc_sel_0_0),
    .io_req_2_0_bits_vc_sel_0_1(switch_allocator_io_req_2_0_bits_vc_sel_0_1),
    .io_req_2_0_bits_vc_sel_0_2(switch_allocator_io_req_2_0_bits_vc_sel_0_2),
    .io_req_2_0_bits_vc_sel_0_3(switch_allocator_io_req_2_0_bits_vc_sel_0_3),
    .io_req_2_0_bits_tail(switch_allocator_io_req_2_0_bits_tail),
    .io_req_1_0_ready(switch_allocator_io_req_1_0_ready),
    .io_req_1_0_valid(switch_allocator_io_req_1_0_valid),
    .io_req_1_0_bits_vc_sel_2_0(switch_allocator_io_req_1_0_bits_vc_sel_2_0),
    .io_req_1_0_bits_vc_sel_1_0(switch_allocator_io_req_1_0_bits_vc_sel_1_0),
    .io_req_1_0_bits_vc_sel_1_1(switch_allocator_io_req_1_0_bits_vc_sel_1_1),
    .io_req_1_0_bits_vc_sel_1_2(switch_allocator_io_req_1_0_bits_vc_sel_1_2),
    .io_req_1_0_bits_vc_sel_1_3(switch_allocator_io_req_1_0_bits_vc_sel_1_3),
    .io_req_1_0_bits_vc_sel_0_0(switch_allocator_io_req_1_0_bits_vc_sel_0_0),
    .io_req_1_0_bits_vc_sel_0_1(switch_allocator_io_req_1_0_bits_vc_sel_0_1),
    .io_req_1_0_bits_vc_sel_0_2(switch_allocator_io_req_1_0_bits_vc_sel_0_2),
    .io_req_1_0_bits_vc_sel_0_3(switch_allocator_io_req_1_0_bits_vc_sel_0_3),
    .io_req_1_0_bits_tail(switch_allocator_io_req_1_0_bits_tail),
    .io_req_0_0_ready(switch_allocator_io_req_0_0_ready),
    .io_req_0_0_valid(switch_allocator_io_req_0_0_valid),
    .io_req_0_0_bits_vc_sel_2_0(switch_allocator_io_req_0_0_bits_vc_sel_2_0),
    .io_req_0_0_bits_vc_sel_1_0(switch_allocator_io_req_0_0_bits_vc_sel_1_0),
    .io_req_0_0_bits_vc_sel_1_1(switch_allocator_io_req_0_0_bits_vc_sel_1_1),
    .io_req_0_0_bits_vc_sel_1_2(switch_allocator_io_req_0_0_bits_vc_sel_1_2),
    .io_req_0_0_bits_vc_sel_1_3(switch_allocator_io_req_0_0_bits_vc_sel_1_3),
    .io_req_0_0_bits_vc_sel_0_0(switch_allocator_io_req_0_0_bits_vc_sel_0_0),
    .io_req_0_0_bits_vc_sel_0_1(switch_allocator_io_req_0_0_bits_vc_sel_0_1),
    .io_req_0_0_bits_vc_sel_0_2(switch_allocator_io_req_0_0_bits_vc_sel_0_2),
    .io_req_0_0_bits_vc_sel_0_3(switch_allocator_io_req_0_0_bits_vc_sel_0_3),
    .io_req_0_0_bits_tail(switch_allocator_io_req_0_0_bits_tail),
    .io_credit_alloc_2_0_alloc(switch_allocator_io_credit_alloc_2_0_alloc),
    .io_credit_alloc_2_0_tail(switch_allocator_io_credit_alloc_2_0_tail),
    .io_credit_alloc_1_0_alloc(switch_allocator_io_credit_alloc_1_0_alloc),
    .io_credit_alloc_1_1_alloc(switch_allocator_io_credit_alloc_1_1_alloc),
    .io_credit_alloc_1_2_alloc(switch_allocator_io_credit_alloc_1_2_alloc),
    .io_credit_alloc_1_3_alloc(switch_allocator_io_credit_alloc_1_3_alloc),
    .io_credit_alloc_0_0_alloc(switch_allocator_io_credit_alloc_0_0_alloc),
    .io_credit_alloc_0_1_alloc(switch_allocator_io_credit_alloc_0_1_alloc),
    .io_credit_alloc_0_2_alloc(switch_allocator_io_credit_alloc_0_2_alloc),
    .io_credit_alloc_0_3_alloc(switch_allocator_io_credit_alloc_0_3_alloc),
    .io_switch_sel_2_0_2_0(switch_allocator_io_switch_sel_2_0_2_0),
    .io_switch_sel_2_0_1_0(switch_allocator_io_switch_sel_2_0_1_0),
    .io_switch_sel_2_0_0_0(switch_allocator_io_switch_sel_2_0_0_0),
    .io_switch_sel_1_0_2_0(switch_allocator_io_switch_sel_1_0_2_0),
    .io_switch_sel_1_0_1_0(switch_allocator_io_switch_sel_1_0_1_0),
    .io_switch_sel_1_0_0_0(switch_allocator_io_switch_sel_1_0_0_0),
    .io_switch_sel_0_0_2_0(switch_allocator_io_switch_sel_0_0_2_0),
    .io_switch_sel_0_0_1_0(switch_allocator_io_switch_sel_0_0_1_0),
    .io_switch_sel_0_0_0_0(switch_allocator_io_switch_sel_0_0_0_0)
  );
  RotatingSingleVCAllocator vc_allocator ( // @[Router.scala 131:30]
    .clock(vc_allocator_clock),
    .reset(vc_allocator_reset),
    .io_req_2_ready(vc_allocator_io_req_2_ready),
    .io_req_2_valid(vc_allocator_io_req_2_valid),
    .io_req_2_bits_vc_sel_2_0(vc_allocator_io_req_2_bits_vc_sel_2_0),
    .io_req_2_bits_vc_sel_1_0(vc_allocator_io_req_2_bits_vc_sel_1_0),
    .io_req_2_bits_vc_sel_1_1(vc_allocator_io_req_2_bits_vc_sel_1_1),
    .io_req_2_bits_vc_sel_1_2(vc_allocator_io_req_2_bits_vc_sel_1_2),
    .io_req_2_bits_vc_sel_1_3(vc_allocator_io_req_2_bits_vc_sel_1_3),
    .io_req_2_bits_vc_sel_0_0(vc_allocator_io_req_2_bits_vc_sel_0_0),
    .io_req_2_bits_vc_sel_0_1(vc_allocator_io_req_2_bits_vc_sel_0_1),
    .io_req_2_bits_vc_sel_0_2(vc_allocator_io_req_2_bits_vc_sel_0_2),
    .io_req_2_bits_vc_sel_0_3(vc_allocator_io_req_2_bits_vc_sel_0_3),
    .io_req_1_ready(vc_allocator_io_req_1_ready),
    .io_req_1_valid(vc_allocator_io_req_1_valid),
    .io_req_1_bits_vc_sel_2_0(vc_allocator_io_req_1_bits_vc_sel_2_0),
    .io_req_1_bits_vc_sel_1_0(vc_allocator_io_req_1_bits_vc_sel_1_0),
    .io_req_1_bits_vc_sel_1_1(vc_allocator_io_req_1_bits_vc_sel_1_1),
    .io_req_1_bits_vc_sel_1_2(vc_allocator_io_req_1_bits_vc_sel_1_2),
    .io_req_1_bits_vc_sel_1_3(vc_allocator_io_req_1_bits_vc_sel_1_3),
    .io_req_1_bits_vc_sel_0_0(vc_allocator_io_req_1_bits_vc_sel_0_0),
    .io_req_1_bits_vc_sel_0_1(vc_allocator_io_req_1_bits_vc_sel_0_1),
    .io_req_1_bits_vc_sel_0_2(vc_allocator_io_req_1_bits_vc_sel_0_2),
    .io_req_1_bits_vc_sel_0_3(vc_allocator_io_req_1_bits_vc_sel_0_3),
    .io_req_0_ready(vc_allocator_io_req_0_ready),
    .io_req_0_valid(vc_allocator_io_req_0_valid),
    .io_req_0_bits_vc_sel_2_0(vc_allocator_io_req_0_bits_vc_sel_2_0),
    .io_req_0_bits_vc_sel_1_0(vc_allocator_io_req_0_bits_vc_sel_1_0),
    .io_req_0_bits_vc_sel_1_1(vc_allocator_io_req_0_bits_vc_sel_1_1),
    .io_req_0_bits_vc_sel_1_2(vc_allocator_io_req_0_bits_vc_sel_1_2),
    .io_req_0_bits_vc_sel_1_3(vc_allocator_io_req_0_bits_vc_sel_1_3),
    .io_req_0_bits_vc_sel_0_0(vc_allocator_io_req_0_bits_vc_sel_0_0),
    .io_req_0_bits_vc_sel_0_1(vc_allocator_io_req_0_bits_vc_sel_0_1),
    .io_req_0_bits_vc_sel_0_2(vc_allocator_io_req_0_bits_vc_sel_0_2),
    .io_req_0_bits_vc_sel_0_3(vc_allocator_io_req_0_bits_vc_sel_0_3),
    .io_resp_2_vc_sel_2_0(vc_allocator_io_resp_2_vc_sel_2_0),
    .io_resp_2_vc_sel_1_0(vc_allocator_io_resp_2_vc_sel_1_0),
    .io_resp_2_vc_sel_1_1(vc_allocator_io_resp_2_vc_sel_1_1),
    .io_resp_2_vc_sel_1_2(vc_allocator_io_resp_2_vc_sel_1_2),
    .io_resp_2_vc_sel_1_3(vc_allocator_io_resp_2_vc_sel_1_3),
    .io_resp_2_vc_sel_0_0(vc_allocator_io_resp_2_vc_sel_0_0),
    .io_resp_2_vc_sel_0_1(vc_allocator_io_resp_2_vc_sel_0_1),
    .io_resp_2_vc_sel_0_2(vc_allocator_io_resp_2_vc_sel_0_2),
    .io_resp_2_vc_sel_0_3(vc_allocator_io_resp_2_vc_sel_0_3),
    .io_resp_1_vc_sel_2_0(vc_allocator_io_resp_1_vc_sel_2_0),
    .io_resp_1_vc_sel_1_0(vc_allocator_io_resp_1_vc_sel_1_0),
    .io_resp_1_vc_sel_1_1(vc_allocator_io_resp_1_vc_sel_1_1),
    .io_resp_1_vc_sel_1_2(vc_allocator_io_resp_1_vc_sel_1_2),
    .io_resp_1_vc_sel_1_3(vc_allocator_io_resp_1_vc_sel_1_3),
    .io_resp_1_vc_sel_0_0(vc_allocator_io_resp_1_vc_sel_0_0),
    .io_resp_1_vc_sel_0_1(vc_allocator_io_resp_1_vc_sel_0_1),
    .io_resp_1_vc_sel_0_2(vc_allocator_io_resp_1_vc_sel_0_2),
    .io_resp_1_vc_sel_0_3(vc_allocator_io_resp_1_vc_sel_0_3),
    .io_resp_0_vc_sel_2_0(vc_allocator_io_resp_0_vc_sel_2_0),
    .io_resp_0_vc_sel_1_0(vc_allocator_io_resp_0_vc_sel_1_0),
    .io_resp_0_vc_sel_1_1(vc_allocator_io_resp_0_vc_sel_1_1),
    .io_resp_0_vc_sel_1_2(vc_allocator_io_resp_0_vc_sel_1_2),
    .io_resp_0_vc_sel_1_3(vc_allocator_io_resp_0_vc_sel_1_3),
    .io_resp_0_vc_sel_0_0(vc_allocator_io_resp_0_vc_sel_0_0),
    .io_resp_0_vc_sel_0_1(vc_allocator_io_resp_0_vc_sel_0_1),
    .io_resp_0_vc_sel_0_2(vc_allocator_io_resp_0_vc_sel_0_2),
    .io_resp_0_vc_sel_0_3(vc_allocator_io_resp_0_vc_sel_0_3),
    .io_channel_status_2_0_occupied(vc_allocator_io_channel_status_2_0_occupied),
    .io_channel_status_1_0_occupied(vc_allocator_io_channel_status_1_0_occupied),
    .io_channel_status_1_1_occupied(vc_allocator_io_channel_status_1_1_occupied),
    .io_channel_status_1_2_occupied(vc_allocator_io_channel_status_1_2_occupied),
    .io_channel_status_1_3_occupied(vc_allocator_io_channel_status_1_3_occupied),
    .io_channel_status_0_0_occupied(vc_allocator_io_channel_status_0_0_occupied),
    .io_channel_status_0_1_occupied(vc_allocator_io_channel_status_0_1_occupied),
    .io_channel_status_0_2_occupied(vc_allocator_io_channel_status_0_2_occupied),
    .io_channel_status_0_3_occupied(vc_allocator_io_channel_status_0_3_occupied),
    .io_out_allocs_2_0_alloc(vc_allocator_io_out_allocs_2_0_alloc),
    .io_out_allocs_1_0_alloc(vc_allocator_io_out_allocs_1_0_alloc),
    .io_out_allocs_1_1_alloc(vc_allocator_io_out_allocs_1_1_alloc),
    .io_out_allocs_1_2_alloc(vc_allocator_io_out_allocs_1_2_alloc),
    .io_out_allocs_1_3_alloc(vc_allocator_io_out_allocs_1_3_alloc),
    .io_out_allocs_0_0_alloc(vc_allocator_io_out_allocs_0_0_alloc),
    .io_out_allocs_0_1_alloc(vc_allocator_io_out_allocs_0_1_alloc),
    .io_out_allocs_0_2_alloc(vc_allocator_io_out_allocs_0_2_alloc),
    .io_out_allocs_0_3_alloc(vc_allocator_io_out_allocs_0_3_alloc)
  );
  RouteComputer_2 route_computer ( // @[Router.scala 134:32]
    .io_req_2_bits_flow_ingress_node(route_computer_io_req_2_bits_flow_ingress_node),
    .io_req_2_bits_flow_egress_node(route_computer_io_req_2_bits_flow_egress_node),
    .io_req_1_bits_src_virt_id(route_computer_io_req_1_bits_src_virt_id),
    .io_req_1_bits_flow_ingress_node(route_computer_io_req_1_bits_flow_ingress_node),
    .io_req_1_bits_flow_egress_node(route_computer_io_req_1_bits_flow_egress_node),
    .io_req_0_bits_src_virt_id(route_computer_io_req_0_bits_src_virt_id),
    .io_req_0_bits_flow_ingress_node(route_computer_io_req_0_bits_flow_ingress_node),
    .io_req_0_bits_flow_egress_node(route_computer_io_req_0_bits_flow_egress_node),
    .io_resp_2_vc_sel_1_0(route_computer_io_resp_2_vc_sel_1_0),
    .io_resp_2_vc_sel_1_1(route_computer_io_resp_2_vc_sel_1_1),
    .io_resp_2_vc_sel_1_2(route_computer_io_resp_2_vc_sel_1_2),
    .io_resp_2_vc_sel_1_3(route_computer_io_resp_2_vc_sel_1_3),
    .io_resp_2_vc_sel_0_0(route_computer_io_resp_2_vc_sel_0_0),
    .io_resp_2_vc_sel_0_1(route_computer_io_resp_2_vc_sel_0_1),
    .io_resp_2_vc_sel_0_2(route_computer_io_resp_2_vc_sel_0_2),
    .io_resp_2_vc_sel_0_3(route_computer_io_resp_2_vc_sel_0_3),
    .io_resp_1_vc_sel_1_0(route_computer_io_resp_1_vc_sel_1_0),
    .io_resp_1_vc_sel_1_1(route_computer_io_resp_1_vc_sel_1_1),
    .io_resp_1_vc_sel_1_2(route_computer_io_resp_1_vc_sel_1_2),
    .io_resp_1_vc_sel_1_3(route_computer_io_resp_1_vc_sel_1_3),
    .io_resp_1_vc_sel_0_0(route_computer_io_resp_1_vc_sel_0_0),
    .io_resp_1_vc_sel_0_1(route_computer_io_resp_1_vc_sel_0_1),
    .io_resp_1_vc_sel_0_2(route_computer_io_resp_1_vc_sel_0_2),
    .io_resp_1_vc_sel_0_3(route_computer_io_resp_1_vc_sel_0_3),
    .io_resp_0_vc_sel_1_0(route_computer_io_resp_0_vc_sel_1_0),
    .io_resp_0_vc_sel_1_1(route_computer_io_resp_0_vc_sel_1_1),
    .io_resp_0_vc_sel_1_2(route_computer_io_resp_0_vc_sel_1_2),
    .io_resp_0_vc_sel_1_3(route_computer_io_resp_0_vc_sel_1_3),
    .io_resp_0_vc_sel_0_0(route_computer_io_resp_0_vc_sel_0_0),
    .io_resp_0_vc_sel_0_1(route_computer_io_resp_0_vc_sel_0_1),
    .io_resp_0_vc_sel_0_2(route_computer_io_resp_0_vc_sel_0_2),
    .io_resp_0_vc_sel_0_3(route_computer_io_resp_0_vc_sel_0_3)
  );
  plusarg_reader #(.FORMAT("noc_util_sample_rate=%d"), .DEFAULT(0), .WIDTH(20)) plusarg_reader ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_out)
  );
  assign auto_debug_out_va_stall_0 = input_unit_0_from_1_io_debug_va_stall; // @[Nodes.scala 1212:84 Router.scala 190:92]
  assign auto_debug_out_va_stall_1 = input_unit_1_from_3_io_debug_va_stall; // @[Nodes.scala 1212:84 Router.scala 190:92]
  assign auto_debug_out_sa_stall_0 = input_unit_0_from_1_io_debug_sa_stall; // @[Nodes.scala 1212:84 Router.scala 191:92]
  assign auto_debug_out_sa_stall_1 = input_unit_1_from_3_io_debug_sa_stall; // @[Nodes.scala 1212:84 Router.scala 191:92]
  assign auto_egress_nodes_out_flit_valid = egress_unit_2_to_2_io_out_valid; // @[Nodes.scala 1212:84 Router.scala 144:65]
  assign auto_egress_nodes_out_flit_bits_head = egress_unit_2_to_2_io_out_bits_head; // @[Nodes.scala 1212:84 Router.scala 144:65]
  assign auto_egress_nodes_out_flit_bits_tail = egress_unit_2_to_2_io_out_bits_tail; // @[Nodes.scala 1212:84 Router.scala 144:65]
  assign auto_egress_nodes_out_flit_bits_payload = egress_unit_2_to_2_io_out_bits_payload; // @[Nodes.scala 1212:84 Router.scala 144:65]
  assign auto_egress_nodes_out_flit_bits_ingress_id = egress_unit_2_to_2_io_out_bits_ingress_id; // @[Nodes.scala 1212:84 Router.scala 144:65]
  assign auto_ingress_nodes_in_flit_ready = ingress_unit_2_from_2_io_in_ready; // @[Nodes.scala 1215:84 Router.scala 142:68]
  assign auto_source_nodes_out_1_flit_0_valid = output_unit_1_to_3_io_out_flit_0_valid; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_1_flit_0_bits_head = output_unit_1_to_3_io_out_flit_0_bits_head; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_1_flit_0_bits_tail = output_unit_1_to_3_io_out_flit_0_bits_tail; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_1_flit_0_bits_payload = output_unit_1_to_3_io_out_flit_0_bits_payload; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_1_flit_0_bits_flow_ingress_node = output_unit_1_to_3_io_out_flit_0_bits_flow_ingress_node
    ; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_1_flit_0_bits_flow_egress_node = output_unit_1_to_3_io_out_flit_0_bits_flow_egress_node; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_1_flit_0_bits_virt_channel_id = output_unit_1_to_3_io_out_flit_0_bits_virt_channel_id; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_0_flit_0_valid = output_unit_0_to_1_io_out_flit_0_valid; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_0_flit_0_bits_head = output_unit_0_to_1_io_out_flit_0_bits_head; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_0_flit_0_bits_tail = output_unit_0_to_1_io_out_flit_0_bits_tail; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_0_flit_0_bits_payload = output_unit_0_to_1_io_out_flit_0_bits_payload; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_0_flit_0_bits_flow_ingress_node = output_unit_0_to_1_io_out_flit_0_bits_flow_ingress_node
    ; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_0_flit_0_bits_flow_egress_node = output_unit_0_to_1_io_out_flit_0_bits_flow_egress_node; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_0_flit_0_bits_virt_channel_id = output_unit_0_to_1_io_out_flit_0_bits_virt_channel_id; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_dest_nodes_in_1_credit_return = input_unit_1_from_3_io_in_credit_return; // @[Nodes.scala 1215:84 Router.scala 141:68]
  assign auto_dest_nodes_in_1_vc_free = input_unit_1_from_3_io_in_vc_free; // @[Nodes.scala 1215:84 Router.scala 141:68]
  assign auto_dest_nodes_in_0_credit_return = input_unit_0_from_1_io_in_credit_return; // @[Nodes.scala 1215:84 Router.scala 141:68]
  assign auto_dest_nodes_in_0_vc_free = input_unit_0_from_1_io_in_vc_free; // @[Nodes.scala 1215:84 Router.scala 141:68]
  assign monitor_clock = clock;
  assign monitor_reset = reset;
  assign monitor_io_in_flit_0_valid = auto_dest_nodes_in_0_flit_0_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_io_in_flit_0_bits_head = auto_dest_nodes_in_0_flit_0_bits_head; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_io_in_flit_0_bits_tail = auto_dest_nodes_in_0_flit_0_bits_tail; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_io_in_flit_0_bits_flow_ingress_node = auto_dest_nodes_in_0_flit_0_bits_flow_ingress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_io_in_flit_0_bits_flow_egress_node = auto_dest_nodes_in_0_flit_0_bits_flow_egress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_io_in_flit_0_bits_virt_channel_id = auto_dest_nodes_in_0_flit_0_bits_virt_channel_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_1_clock = clock;
  assign monitor_1_reset = reset;
  assign monitor_1_io_in_flit_0_valid = auto_dest_nodes_in_1_flit_0_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_1_io_in_flit_0_bits_head = auto_dest_nodes_in_1_flit_0_bits_head; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_1_io_in_flit_0_bits_tail = auto_dest_nodes_in_1_flit_0_bits_tail; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_1_io_in_flit_0_bits_flow_ingress_node = auto_dest_nodes_in_1_flit_0_bits_flow_ingress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_1_io_in_flit_0_bits_flow_egress_node = auto_dest_nodes_in_1_flit_0_bits_flow_egress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_1_io_in_flit_0_bits_virt_channel_id = auto_dest_nodes_in_1_flit_0_bits_virt_channel_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_1_clock = clock;
  assign input_unit_0_from_1_reset = reset;
  assign input_unit_0_from_1_io_router_resp_vc_sel_1_0 = route_computer_io_resp_0_vc_sel_1_0; // @[Router.scala 148:38]
  assign input_unit_0_from_1_io_router_resp_vc_sel_1_1 = route_computer_io_resp_0_vc_sel_1_1; // @[Router.scala 148:38]
  assign input_unit_0_from_1_io_router_resp_vc_sel_1_2 = route_computer_io_resp_0_vc_sel_1_2; // @[Router.scala 148:38]
  assign input_unit_0_from_1_io_router_resp_vc_sel_1_3 = route_computer_io_resp_0_vc_sel_1_3; // @[Router.scala 148:38]
  assign input_unit_0_from_1_io_router_resp_vc_sel_0_0 = route_computer_io_resp_0_vc_sel_0_0; // @[Router.scala 148:38]
  assign input_unit_0_from_1_io_router_resp_vc_sel_0_1 = route_computer_io_resp_0_vc_sel_0_1; // @[Router.scala 148:38]
  assign input_unit_0_from_1_io_router_resp_vc_sel_0_2 = route_computer_io_resp_0_vc_sel_0_2; // @[Router.scala 148:38]
  assign input_unit_0_from_1_io_router_resp_vc_sel_0_3 = route_computer_io_resp_0_vc_sel_0_3; // @[Router.scala 148:38]
  assign input_unit_0_from_1_io_vcalloc_req_ready = vc_allocator_io_req_0_ready; // @[Router.scala 151:23]
  assign input_unit_0_from_1_io_vcalloc_resp_vc_sel_2_0 = vc_allocator_io_resp_0_vc_sel_2_0; // @[Router.scala 153:39]
  assign input_unit_0_from_1_io_vcalloc_resp_vc_sel_1_0 = vc_allocator_io_resp_0_vc_sel_1_0; // @[Router.scala 153:39]
  assign input_unit_0_from_1_io_vcalloc_resp_vc_sel_1_1 = vc_allocator_io_resp_0_vc_sel_1_1; // @[Router.scala 153:39]
  assign input_unit_0_from_1_io_vcalloc_resp_vc_sel_1_2 = vc_allocator_io_resp_0_vc_sel_1_2; // @[Router.scala 153:39]
  assign input_unit_0_from_1_io_vcalloc_resp_vc_sel_1_3 = vc_allocator_io_resp_0_vc_sel_1_3; // @[Router.scala 153:39]
  assign input_unit_0_from_1_io_vcalloc_resp_vc_sel_0_0 = vc_allocator_io_resp_0_vc_sel_0_0; // @[Router.scala 153:39]
  assign input_unit_0_from_1_io_vcalloc_resp_vc_sel_0_1 = vc_allocator_io_resp_0_vc_sel_0_1; // @[Router.scala 153:39]
  assign input_unit_0_from_1_io_vcalloc_resp_vc_sel_0_2 = vc_allocator_io_resp_0_vc_sel_0_2; // @[Router.scala 153:39]
  assign input_unit_0_from_1_io_vcalloc_resp_vc_sel_0_3 = vc_allocator_io_resp_0_vc_sel_0_3; // @[Router.scala 153:39]
  assign input_unit_0_from_1_io_out_credit_available_2_0 = egress_unit_2_to_2_io_credit_available_0; // @[Router.scala 162:42]
  assign input_unit_0_from_1_io_out_credit_available_1_0 = output_unit_1_to_3_io_credit_available_0; // @[Router.scala 162:42]
  assign input_unit_0_from_1_io_out_credit_available_1_1 = output_unit_1_to_3_io_credit_available_1; // @[Router.scala 162:42]
  assign input_unit_0_from_1_io_out_credit_available_1_2 = output_unit_1_to_3_io_credit_available_2; // @[Router.scala 162:42]
  assign input_unit_0_from_1_io_out_credit_available_1_3 = output_unit_1_to_3_io_credit_available_3; // @[Router.scala 162:42]
  assign input_unit_0_from_1_io_out_credit_available_0_0 = output_unit_0_to_1_io_credit_available_0; // @[Router.scala 162:42]
  assign input_unit_0_from_1_io_out_credit_available_0_1 = output_unit_0_to_1_io_credit_available_1; // @[Router.scala 162:42]
  assign input_unit_0_from_1_io_out_credit_available_0_2 = output_unit_0_to_1_io_credit_available_2; // @[Router.scala 162:42]
  assign input_unit_0_from_1_io_out_credit_available_0_3 = output_unit_0_to_1_io_credit_available_3; // @[Router.scala 162:42]
  assign input_unit_0_from_1_io_salloc_req_0_ready = switch_allocator_io_req_0_0_ready; // @[Router.scala 165:23]
  assign input_unit_0_from_1_io_in_flit_0_valid = auto_dest_nodes_in_0_flit_0_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_1_io_in_flit_0_bits_head = auto_dest_nodes_in_0_flit_0_bits_head; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_1_io_in_flit_0_bits_tail = auto_dest_nodes_in_0_flit_0_bits_tail; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_1_io_in_flit_0_bits_payload = auto_dest_nodes_in_0_flit_0_bits_payload; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_1_io_in_flit_0_bits_flow_ingress_node = auto_dest_nodes_in_0_flit_0_bits_flow_ingress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_1_io_in_flit_0_bits_flow_egress_node = auto_dest_nodes_in_0_flit_0_bits_flow_egress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_1_io_in_flit_0_bits_virt_channel_id = auto_dest_nodes_in_0_flit_0_bits_virt_channel_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_1_from_3_clock = clock;
  assign input_unit_1_from_3_reset = reset;
  assign input_unit_1_from_3_io_router_resp_vc_sel_1_0 = route_computer_io_resp_1_vc_sel_1_0; // @[Router.scala 148:38]
  assign input_unit_1_from_3_io_router_resp_vc_sel_1_1 = route_computer_io_resp_1_vc_sel_1_1; // @[Router.scala 148:38]
  assign input_unit_1_from_3_io_router_resp_vc_sel_1_2 = route_computer_io_resp_1_vc_sel_1_2; // @[Router.scala 148:38]
  assign input_unit_1_from_3_io_router_resp_vc_sel_1_3 = route_computer_io_resp_1_vc_sel_1_3; // @[Router.scala 148:38]
  assign input_unit_1_from_3_io_router_resp_vc_sel_0_0 = route_computer_io_resp_1_vc_sel_0_0; // @[Router.scala 148:38]
  assign input_unit_1_from_3_io_router_resp_vc_sel_0_1 = route_computer_io_resp_1_vc_sel_0_1; // @[Router.scala 148:38]
  assign input_unit_1_from_3_io_router_resp_vc_sel_0_2 = route_computer_io_resp_1_vc_sel_0_2; // @[Router.scala 148:38]
  assign input_unit_1_from_3_io_router_resp_vc_sel_0_3 = route_computer_io_resp_1_vc_sel_0_3; // @[Router.scala 148:38]
  assign input_unit_1_from_3_io_vcalloc_req_ready = vc_allocator_io_req_1_ready; // @[Router.scala 151:23]
  assign input_unit_1_from_3_io_vcalloc_resp_vc_sel_2_0 = vc_allocator_io_resp_1_vc_sel_2_0; // @[Router.scala 153:39]
  assign input_unit_1_from_3_io_vcalloc_resp_vc_sel_1_0 = vc_allocator_io_resp_1_vc_sel_1_0; // @[Router.scala 153:39]
  assign input_unit_1_from_3_io_vcalloc_resp_vc_sel_1_1 = vc_allocator_io_resp_1_vc_sel_1_1; // @[Router.scala 153:39]
  assign input_unit_1_from_3_io_vcalloc_resp_vc_sel_1_2 = vc_allocator_io_resp_1_vc_sel_1_2; // @[Router.scala 153:39]
  assign input_unit_1_from_3_io_vcalloc_resp_vc_sel_1_3 = vc_allocator_io_resp_1_vc_sel_1_3; // @[Router.scala 153:39]
  assign input_unit_1_from_3_io_vcalloc_resp_vc_sel_0_0 = vc_allocator_io_resp_1_vc_sel_0_0; // @[Router.scala 153:39]
  assign input_unit_1_from_3_io_vcalloc_resp_vc_sel_0_1 = vc_allocator_io_resp_1_vc_sel_0_1; // @[Router.scala 153:39]
  assign input_unit_1_from_3_io_vcalloc_resp_vc_sel_0_2 = vc_allocator_io_resp_1_vc_sel_0_2; // @[Router.scala 153:39]
  assign input_unit_1_from_3_io_vcalloc_resp_vc_sel_0_3 = vc_allocator_io_resp_1_vc_sel_0_3; // @[Router.scala 153:39]
  assign input_unit_1_from_3_io_out_credit_available_2_0 = egress_unit_2_to_2_io_credit_available_0; // @[Router.scala 162:42]
  assign input_unit_1_from_3_io_out_credit_available_1_0 = output_unit_1_to_3_io_credit_available_0; // @[Router.scala 162:42]
  assign input_unit_1_from_3_io_out_credit_available_1_1 = output_unit_1_to_3_io_credit_available_1; // @[Router.scala 162:42]
  assign input_unit_1_from_3_io_out_credit_available_1_2 = output_unit_1_to_3_io_credit_available_2; // @[Router.scala 162:42]
  assign input_unit_1_from_3_io_out_credit_available_1_3 = output_unit_1_to_3_io_credit_available_3; // @[Router.scala 162:42]
  assign input_unit_1_from_3_io_out_credit_available_0_0 = output_unit_0_to_1_io_credit_available_0; // @[Router.scala 162:42]
  assign input_unit_1_from_3_io_out_credit_available_0_1 = output_unit_0_to_1_io_credit_available_1; // @[Router.scala 162:42]
  assign input_unit_1_from_3_io_out_credit_available_0_2 = output_unit_0_to_1_io_credit_available_2; // @[Router.scala 162:42]
  assign input_unit_1_from_3_io_out_credit_available_0_3 = output_unit_0_to_1_io_credit_available_3; // @[Router.scala 162:42]
  assign input_unit_1_from_3_io_salloc_req_0_ready = switch_allocator_io_req_1_0_ready; // @[Router.scala 165:23]
  assign input_unit_1_from_3_io_in_flit_0_valid = auto_dest_nodes_in_1_flit_0_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_1_from_3_io_in_flit_0_bits_head = auto_dest_nodes_in_1_flit_0_bits_head; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_1_from_3_io_in_flit_0_bits_tail = auto_dest_nodes_in_1_flit_0_bits_tail; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_1_from_3_io_in_flit_0_bits_payload = auto_dest_nodes_in_1_flit_0_bits_payload; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_1_from_3_io_in_flit_0_bits_flow_ingress_node = auto_dest_nodes_in_1_flit_0_bits_flow_ingress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_1_from_3_io_in_flit_0_bits_flow_egress_node = auto_dest_nodes_in_1_flit_0_bits_flow_egress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_1_from_3_io_in_flit_0_bits_virt_channel_id = auto_dest_nodes_in_1_flit_0_bits_virt_channel_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign ingress_unit_2_from_2_clock = clock;
  assign ingress_unit_2_from_2_reset = reset;
  assign ingress_unit_2_from_2_io_router_resp_vc_sel_1_0 = route_computer_io_resp_2_vc_sel_1_0; // @[Router.scala 148:38]
  assign ingress_unit_2_from_2_io_router_resp_vc_sel_1_1 = route_computer_io_resp_2_vc_sel_1_1; // @[Router.scala 148:38]
  assign ingress_unit_2_from_2_io_router_resp_vc_sel_1_2 = route_computer_io_resp_2_vc_sel_1_2; // @[Router.scala 148:38]
  assign ingress_unit_2_from_2_io_router_resp_vc_sel_1_3 = route_computer_io_resp_2_vc_sel_1_3; // @[Router.scala 148:38]
  assign ingress_unit_2_from_2_io_router_resp_vc_sel_0_0 = route_computer_io_resp_2_vc_sel_0_0; // @[Router.scala 148:38]
  assign ingress_unit_2_from_2_io_router_resp_vc_sel_0_1 = route_computer_io_resp_2_vc_sel_0_1; // @[Router.scala 148:38]
  assign ingress_unit_2_from_2_io_router_resp_vc_sel_0_2 = route_computer_io_resp_2_vc_sel_0_2; // @[Router.scala 148:38]
  assign ingress_unit_2_from_2_io_router_resp_vc_sel_0_3 = route_computer_io_resp_2_vc_sel_0_3; // @[Router.scala 148:38]
  assign ingress_unit_2_from_2_io_vcalloc_req_ready = vc_allocator_io_req_2_ready; // @[Router.scala 151:23]
  assign ingress_unit_2_from_2_io_vcalloc_resp_vc_sel_2_0 = vc_allocator_io_resp_2_vc_sel_2_0; // @[Router.scala 153:39]
  assign ingress_unit_2_from_2_io_vcalloc_resp_vc_sel_1_0 = vc_allocator_io_resp_2_vc_sel_1_0; // @[Router.scala 153:39]
  assign ingress_unit_2_from_2_io_vcalloc_resp_vc_sel_1_1 = vc_allocator_io_resp_2_vc_sel_1_1; // @[Router.scala 153:39]
  assign ingress_unit_2_from_2_io_vcalloc_resp_vc_sel_1_2 = vc_allocator_io_resp_2_vc_sel_1_2; // @[Router.scala 153:39]
  assign ingress_unit_2_from_2_io_vcalloc_resp_vc_sel_1_3 = vc_allocator_io_resp_2_vc_sel_1_3; // @[Router.scala 153:39]
  assign ingress_unit_2_from_2_io_vcalloc_resp_vc_sel_0_0 = vc_allocator_io_resp_2_vc_sel_0_0; // @[Router.scala 153:39]
  assign ingress_unit_2_from_2_io_vcalloc_resp_vc_sel_0_1 = vc_allocator_io_resp_2_vc_sel_0_1; // @[Router.scala 153:39]
  assign ingress_unit_2_from_2_io_vcalloc_resp_vc_sel_0_2 = vc_allocator_io_resp_2_vc_sel_0_2; // @[Router.scala 153:39]
  assign ingress_unit_2_from_2_io_vcalloc_resp_vc_sel_0_3 = vc_allocator_io_resp_2_vc_sel_0_3; // @[Router.scala 153:39]
  assign ingress_unit_2_from_2_io_out_credit_available_2_0 = egress_unit_2_to_2_io_credit_available_0; // @[Router.scala 162:42]
  assign ingress_unit_2_from_2_io_out_credit_available_1_0 = output_unit_1_to_3_io_credit_available_0; // @[Router.scala 162:42]
  assign ingress_unit_2_from_2_io_out_credit_available_1_1 = output_unit_1_to_3_io_credit_available_1; // @[Router.scala 162:42]
  assign ingress_unit_2_from_2_io_out_credit_available_1_2 = output_unit_1_to_3_io_credit_available_2; // @[Router.scala 162:42]
  assign ingress_unit_2_from_2_io_out_credit_available_1_3 = output_unit_1_to_3_io_credit_available_3; // @[Router.scala 162:42]
  assign ingress_unit_2_from_2_io_out_credit_available_0_0 = output_unit_0_to_1_io_credit_available_0; // @[Router.scala 162:42]
  assign ingress_unit_2_from_2_io_out_credit_available_0_1 = output_unit_0_to_1_io_credit_available_1; // @[Router.scala 162:42]
  assign ingress_unit_2_from_2_io_out_credit_available_0_2 = output_unit_0_to_1_io_credit_available_2; // @[Router.scala 162:42]
  assign ingress_unit_2_from_2_io_out_credit_available_0_3 = output_unit_0_to_1_io_credit_available_3; // @[Router.scala 162:42]
  assign ingress_unit_2_from_2_io_salloc_req_0_ready = switch_allocator_io_req_2_0_ready; // @[Router.scala 165:23]
  assign ingress_unit_2_from_2_io_in_valid = auto_ingress_nodes_in_flit_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign ingress_unit_2_from_2_io_in_bits_head = auto_ingress_nodes_in_flit_bits_head; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign ingress_unit_2_from_2_io_in_bits_tail = auto_ingress_nodes_in_flit_bits_tail; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign ingress_unit_2_from_2_io_in_bits_payload = auto_ingress_nodes_in_flit_bits_payload; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign ingress_unit_2_from_2_io_in_bits_egress_id = auto_ingress_nodes_in_flit_bits_egress_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign output_unit_0_to_1_clock = clock;
  assign output_unit_0_to_1_reset = reset;
  assign output_unit_0_to_1_io_in_0_valid = switch_io_out_0_0_valid; // @[Router.scala 172:29]
  assign output_unit_0_to_1_io_in_0_bits_head = switch_io_out_0_0_bits_head; // @[Router.scala 172:29]
  assign output_unit_0_to_1_io_in_0_bits_tail = switch_io_out_0_0_bits_tail; // @[Router.scala 172:29]
  assign output_unit_0_to_1_io_in_0_bits_payload = switch_io_out_0_0_bits_payload; // @[Router.scala 172:29]
  assign output_unit_0_to_1_io_in_0_bits_flow_ingress_node = switch_io_out_0_0_bits_flow_ingress_node; // @[Router.scala 172:29]
  assign output_unit_0_to_1_io_in_0_bits_flow_egress_node = switch_io_out_0_0_bits_flow_egress_node; // @[Router.scala 172:29]
  assign output_unit_0_to_1_io_in_0_bits_virt_channel_id = switch_io_out_0_0_bits_virt_channel_id; // @[Router.scala 172:29]
  assign output_unit_0_to_1_io_allocs_0_alloc = vc_allocator_io_out_allocs_0_0_alloc; // @[Router.scala 157:33]
  assign output_unit_0_to_1_io_allocs_1_alloc = vc_allocator_io_out_allocs_0_1_alloc; // @[Router.scala 157:33]
  assign output_unit_0_to_1_io_allocs_2_alloc = vc_allocator_io_out_allocs_0_2_alloc; // @[Router.scala 157:33]
  assign output_unit_0_to_1_io_allocs_3_alloc = vc_allocator_io_out_allocs_0_3_alloc; // @[Router.scala 157:33]
  assign output_unit_0_to_1_io_credit_alloc_0_alloc = switch_allocator_io_credit_alloc_0_0_alloc; // @[Router.scala 167:39]
  assign output_unit_0_to_1_io_credit_alloc_1_alloc = switch_allocator_io_credit_alloc_0_1_alloc; // @[Router.scala 167:39]
  assign output_unit_0_to_1_io_credit_alloc_2_alloc = switch_allocator_io_credit_alloc_0_2_alloc; // @[Router.scala 167:39]
  assign output_unit_0_to_1_io_credit_alloc_3_alloc = switch_allocator_io_credit_alloc_0_3_alloc; // @[Router.scala 167:39]
  assign output_unit_0_to_1_io_out_credit_return = auto_source_nodes_out_0_credit_return; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign output_unit_0_to_1_io_out_vc_free = auto_source_nodes_out_0_vc_free; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign output_unit_1_to_3_clock = clock;
  assign output_unit_1_to_3_reset = reset;
  assign output_unit_1_to_3_io_in_0_valid = switch_io_out_1_0_valid; // @[Router.scala 172:29]
  assign output_unit_1_to_3_io_in_0_bits_head = switch_io_out_1_0_bits_head; // @[Router.scala 172:29]
  assign output_unit_1_to_3_io_in_0_bits_tail = switch_io_out_1_0_bits_tail; // @[Router.scala 172:29]
  assign output_unit_1_to_3_io_in_0_bits_payload = switch_io_out_1_0_bits_payload; // @[Router.scala 172:29]
  assign output_unit_1_to_3_io_in_0_bits_flow_ingress_node = switch_io_out_1_0_bits_flow_ingress_node; // @[Router.scala 172:29]
  assign output_unit_1_to_3_io_in_0_bits_flow_egress_node = switch_io_out_1_0_bits_flow_egress_node; // @[Router.scala 172:29]
  assign output_unit_1_to_3_io_in_0_bits_virt_channel_id = switch_io_out_1_0_bits_virt_channel_id; // @[Router.scala 172:29]
  assign output_unit_1_to_3_io_allocs_0_alloc = vc_allocator_io_out_allocs_1_0_alloc; // @[Router.scala 157:33]
  assign output_unit_1_to_3_io_allocs_1_alloc = vc_allocator_io_out_allocs_1_1_alloc; // @[Router.scala 157:33]
  assign output_unit_1_to_3_io_allocs_2_alloc = vc_allocator_io_out_allocs_1_2_alloc; // @[Router.scala 157:33]
  assign output_unit_1_to_3_io_allocs_3_alloc = vc_allocator_io_out_allocs_1_3_alloc; // @[Router.scala 157:33]
  assign output_unit_1_to_3_io_credit_alloc_0_alloc = switch_allocator_io_credit_alloc_1_0_alloc; // @[Router.scala 167:39]
  assign output_unit_1_to_3_io_credit_alloc_1_alloc = switch_allocator_io_credit_alloc_1_1_alloc; // @[Router.scala 167:39]
  assign output_unit_1_to_3_io_credit_alloc_2_alloc = switch_allocator_io_credit_alloc_1_2_alloc; // @[Router.scala 167:39]
  assign output_unit_1_to_3_io_credit_alloc_3_alloc = switch_allocator_io_credit_alloc_1_3_alloc; // @[Router.scala 167:39]
  assign output_unit_1_to_3_io_out_credit_return = auto_source_nodes_out_1_credit_return; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign output_unit_1_to_3_io_out_vc_free = auto_source_nodes_out_1_vc_free; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign egress_unit_2_to_2_clock = clock;
  assign egress_unit_2_to_2_reset = reset;
  assign egress_unit_2_to_2_io_in_0_valid = switch_io_out_2_0_valid; // @[Router.scala 172:29]
  assign egress_unit_2_to_2_io_in_0_bits_head = switch_io_out_2_0_bits_head; // @[Router.scala 172:29]
  assign egress_unit_2_to_2_io_in_0_bits_tail = switch_io_out_2_0_bits_tail; // @[Router.scala 172:29]
  assign egress_unit_2_to_2_io_in_0_bits_payload = switch_io_out_2_0_bits_payload; // @[Router.scala 172:29]
  assign egress_unit_2_to_2_io_in_0_bits_flow_ingress_node = switch_io_out_2_0_bits_flow_ingress_node; // @[Router.scala 172:29]
  assign egress_unit_2_to_2_io_allocs_0_alloc = vc_allocator_io_out_allocs_2_0_alloc; // @[Router.scala 157:33]
  assign egress_unit_2_to_2_io_credit_alloc_0_alloc = switch_allocator_io_credit_alloc_2_0_alloc; // @[Router.scala 167:39]
  assign egress_unit_2_to_2_io_credit_alloc_0_tail = switch_allocator_io_credit_alloc_2_0_tail; // @[Router.scala 167:39]
  assign switch_clock = clock;
  assign switch_reset = reset;
  assign switch_io_in_2_0_valid = ingress_unit_2_from_2_io_out_0_valid; // @[Router.scala 170:23]
  assign switch_io_in_2_0_bits_flit_head = ingress_unit_2_from_2_io_out_0_bits_flit_head; // @[Router.scala 170:23]
  assign switch_io_in_2_0_bits_flit_tail = ingress_unit_2_from_2_io_out_0_bits_flit_tail; // @[Router.scala 170:23]
  assign switch_io_in_2_0_bits_flit_payload = ingress_unit_2_from_2_io_out_0_bits_flit_payload; // @[Router.scala 170:23]
  assign switch_io_in_2_0_bits_flit_flow_ingress_node = ingress_unit_2_from_2_io_out_0_bits_flit_flow_ingress_node; // @[Router.scala 170:23]
  assign switch_io_in_2_0_bits_flit_flow_egress_node = ingress_unit_2_from_2_io_out_0_bits_flit_flow_egress_node; // @[Router.scala 170:23]
  assign switch_io_in_2_0_bits_out_virt_channel = ingress_unit_2_from_2_io_out_0_bits_out_virt_channel; // @[Router.scala 170:23]
  assign switch_io_in_1_0_valid = input_unit_1_from_3_io_out_0_valid; // @[Router.scala 170:23]
  assign switch_io_in_1_0_bits_flit_head = input_unit_1_from_3_io_out_0_bits_flit_head; // @[Router.scala 170:23]
  assign switch_io_in_1_0_bits_flit_tail = input_unit_1_from_3_io_out_0_bits_flit_tail; // @[Router.scala 170:23]
  assign switch_io_in_1_0_bits_flit_payload = input_unit_1_from_3_io_out_0_bits_flit_payload; // @[Router.scala 170:23]
  assign switch_io_in_1_0_bits_flit_flow_ingress_node = input_unit_1_from_3_io_out_0_bits_flit_flow_ingress_node; // @[Router.scala 170:23]
  assign switch_io_in_1_0_bits_flit_flow_egress_node = input_unit_1_from_3_io_out_0_bits_flit_flow_egress_node; // @[Router.scala 170:23]
  assign switch_io_in_1_0_bits_out_virt_channel = input_unit_1_from_3_io_out_0_bits_out_virt_channel; // @[Router.scala 170:23]
  assign switch_io_in_0_0_valid = input_unit_0_from_1_io_out_0_valid; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_head = input_unit_0_from_1_io_out_0_bits_flit_head; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_tail = input_unit_0_from_1_io_out_0_bits_flit_tail; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_payload = input_unit_0_from_1_io_out_0_bits_flit_payload; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_flow_ingress_node = input_unit_0_from_1_io_out_0_bits_flit_flow_ingress_node; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_flow_egress_node = input_unit_0_from_1_io_out_0_bits_flit_flow_egress_node; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_out_virt_channel = input_unit_0_from_1_io_out_0_bits_out_virt_channel; // @[Router.scala 170:23]
  assign switch_io_sel_2_0_2_0 = switch_io_sel_REG_2_0_2_0; // @[Router.scala 173:19]
  assign switch_io_sel_2_0_1_0 = switch_io_sel_REG_2_0_1_0; // @[Router.scala 173:19]
  assign switch_io_sel_2_0_0_0 = switch_io_sel_REG_2_0_0_0; // @[Router.scala 173:19]
  assign switch_io_sel_1_0_2_0 = switch_io_sel_REG_1_0_2_0; // @[Router.scala 173:19]
  assign switch_io_sel_1_0_1_0 = switch_io_sel_REG_1_0_1_0; // @[Router.scala 173:19]
  assign switch_io_sel_1_0_0_0 = switch_io_sel_REG_1_0_0_0; // @[Router.scala 173:19]
  assign switch_io_sel_0_0_2_0 = switch_io_sel_REG_0_0_2_0; // @[Router.scala 173:19]
  assign switch_io_sel_0_0_1_0 = switch_io_sel_REG_0_0_1_0; // @[Router.scala 173:19]
  assign switch_io_sel_0_0_0_0 = switch_io_sel_REG_0_0_0_0; // @[Router.scala 173:19]
  assign switch_allocator_clock = clock;
  assign switch_allocator_reset = reset;
  assign switch_allocator_io_req_2_0_valid = ingress_unit_2_from_2_io_salloc_req_0_valid; // @[Router.scala 165:23]
  assign switch_allocator_io_req_2_0_bits_vc_sel_2_0 = ingress_unit_2_from_2_io_salloc_req_0_bits_vc_sel_2_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_2_0_bits_vc_sel_1_0 = ingress_unit_2_from_2_io_salloc_req_0_bits_vc_sel_1_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_2_0_bits_vc_sel_1_1 = ingress_unit_2_from_2_io_salloc_req_0_bits_vc_sel_1_1; // @[Router.scala 165:23]
  assign switch_allocator_io_req_2_0_bits_vc_sel_1_2 = ingress_unit_2_from_2_io_salloc_req_0_bits_vc_sel_1_2; // @[Router.scala 165:23]
  assign switch_allocator_io_req_2_0_bits_vc_sel_1_3 = ingress_unit_2_from_2_io_salloc_req_0_bits_vc_sel_1_3; // @[Router.scala 165:23]
  assign switch_allocator_io_req_2_0_bits_vc_sel_0_0 = ingress_unit_2_from_2_io_salloc_req_0_bits_vc_sel_0_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_2_0_bits_vc_sel_0_1 = ingress_unit_2_from_2_io_salloc_req_0_bits_vc_sel_0_1; // @[Router.scala 165:23]
  assign switch_allocator_io_req_2_0_bits_vc_sel_0_2 = ingress_unit_2_from_2_io_salloc_req_0_bits_vc_sel_0_2; // @[Router.scala 165:23]
  assign switch_allocator_io_req_2_0_bits_vc_sel_0_3 = ingress_unit_2_from_2_io_salloc_req_0_bits_vc_sel_0_3; // @[Router.scala 165:23]
  assign switch_allocator_io_req_2_0_bits_tail = ingress_unit_2_from_2_io_salloc_req_0_bits_tail; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_valid = input_unit_1_from_3_io_salloc_req_0_valid; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_vc_sel_2_0 = input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_2_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_vc_sel_1_0 = input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_1_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_vc_sel_1_1 = input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_1_1; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_vc_sel_1_2 = input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_1_2; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_vc_sel_1_3 = input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_1_3; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_vc_sel_0_0 = input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_0_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_vc_sel_0_1 = input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_0_1; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_vc_sel_0_2 = input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_0_2; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_vc_sel_0_3 = input_unit_1_from_3_io_salloc_req_0_bits_vc_sel_0_3; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_tail = input_unit_1_from_3_io_salloc_req_0_bits_tail; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_valid = input_unit_0_from_1_io_salloc_req_0_valid; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_2_0 = input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_2_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_1_0 = input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_1_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_1_1 = input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_1_1; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_1_2 = input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_1_2; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_1_3 = input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_1_3; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_0_0 = input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_0_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_0_1 = input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_0_1; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_0_2 = input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_0_2; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_0_3 = input_unit_0_from_1_io_salloc_req_0_bits_vc_sel_0_3; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_tail = input_unit_0_from_1_io_salloc_req_0_bits_tail; // @[Router.scala 165:23]
  assign vc_allocator_clock = clock;
  assign vc_allocator_reset = reset;
  assign vc_allocator_io_req_2_valid = ingress_unit_2_from_2_io_vcalloc_req_valid; // @[Router.scala 151:23]
  assign vc_allocator_io_req_2_bits_vc_sel_2_0 = ingress_unit_2_from_2_io_vcalloc_req_bits_vc_sel_2_0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_2_bits_vc_sel_1_0 = ingress_unit_2_from_2_io_vcalloc_req_bits_vc_sel_1_0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_2_bits_vc_sel_1_1 = ingress_unit_2_from_2_io_vcalloc_req_bits_vc_sel_1_1; // @[Router.scala 151:23]
  assign vc_allocator_io_req_2_bits_vc_sel_1_2 = ingress_unit_2_from_2_io_vcalloc_req_bits_vc_sel_1_2; // @[Router.scala 151:23]
  assign vc_allocator_io_req_2_bits_vc_sel_1_3 = ingress_unit_2_from_2_io_vcalloc_req_bits_vc_sel_1_3; // @[Router.scala 151:23]
  assign vc_allocator_io_req_2_bits_vc_sel_0_0 = ingress_unit_2_from_2_io_vcalloc_req_bits_vc_sel_0_0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_2_bits_vc_sel_0_1 = ingress_unit_2_from_2_io_vcalloc_req_bits_vc_sel_0_1; // @[Router.scala 151:23]
  assign vc_allocator_io_req_2_bits_vc_sel_0_2 = ingress_unit_2_from_2_io_vcalloc_req_bits_vc_sel_0_2; // @[Router.scala 151:23]
  assign vc_allocator_io_req_2_bits_vc_sel_0_3 = ingress_unit_2_from_2_io_vcalloc_req_bits_vc_sel_0_3; // @[Router.scala 151:23]
  assign vc_allocator_io_req_1_valid = input_unit_1_from_3_io_vcalloc_req_valid; // @[Router.scala 151:23]
  assign vc_allocator_io_req_1_bits_vc_sel_2_0 = input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_2_0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_1_bits_vc_sel_1_0 = input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_1_0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_1_bits_vc_sel_1_1 = input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_1_1; // @[Router.scala 151:23]
  assign vc_allocator_io_req_1_bits_vc_sel_1_2 = input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_1_2; // @[Router.scala 151:23]
  assign vc_allocator_io_req_1_bits_vc_sel_1_3 = input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_1_3; // @[Router.scala 151:23]
  assign vc_allocator_io_req_1_bits_vc_sel_0_0 = input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_0_0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_1_bits_vc_sel_0_1 = input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_0_1; // @[Router.scala 151:23]
  assign vc_allocator_io_req_1_bits_vc_sel_0_2 = input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_0_2; // @[Router.scala 151:23]
  assign vc_allocator_io_req_1_bits_vc_sel_0_3 = input_unit_1_from_3_io_vcalloc_req_bits_vc_sel_0_3; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_valid = input_unit_0_from_1_io_vcalloc_req_valid; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_2_0 = input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_2_0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_1_0 = input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_1_0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_1_1 = input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_1_1; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_1_2 = input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_1_2; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_1_3 = input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_1_3; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_0_0 = input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_0_0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_0_1 = input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_0_1; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_0_2 = input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_0_2; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_0_3 = input_unit_0_from_1_io_vcalloc_req_bits_vc_sel_0_3; // @[Router.scala 151:23]
  assign vc_allocator_io_channel_status_2_0_occupied = egress_unit_2_to_2_io_channel_status_0_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_1_0_occupied = output_unit_1_to_3_io_channel_status_0_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_1_1_occupied = output_unit_1_to_3_io_channel_status_1_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_1_2_occupied = output_unit_1_to_3_io_channel_status_2_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_1_3_occupied = output_unit_1_to_3_io_channel_status_3_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_0_0_occupied = output_unit_0_to_1_io_channel_status_0_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_0_1_occupied = output_unit_0_to_1_io_channel_status_1_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_0_2_occupied = output_unit_0_to_1_io_channel_status_2_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_0_3_occupied = output_unit_0_to_1_io_channel_status_3_occupied; // @[Router.scala 159:23]
  assign route_computer_io_req_2_bits_flow_ingress_node = ingress_unit_2_from_2_io_router_req_bits_flow_ingress_node; // @[Router.scala 146:23]
  assign route_computer_io_req_2_bits_flow_egress_node = ingress_unit_2_from_2_io_router_req_bits_flow_egress_node; // @[Router.scala 146:23]
  assign route_computer_io_req_1_bits_src_virt_id = input_unit_1_from_3_io_router_req_bits_src_virt_id; // @[Router.scala 146:23]
  assign route_computer_io_req_1_bits_flow_ingress_node = input_unit_1_from_3_io_router_req_bits_flow_ingress_node; // @[Router.scala 146:23]
  assign route_computer_io_req_1_bits_flow_egress_node = input_unit_1_from_3_io_router_req_bits_flow_egress_node; // @[Router.scala 146:23]
  assign route_computer_io_req_0_bits_src_virt_id = input_unit_0_from_1_io_router_req_bits_src_virt_id; // @[Router.scala 146:23]
  assign route_computer_io_req_0_bits_flow_ingress_node = input_unit_0_from_1_io_router_req_bits_flow_ingress_node; // @[Router.scala 146:23]
  assign route_computer_io_req_0_bits_flow_egress_node = input_unit_0_from_1_io_router_req_bits_flow_egress_node; // @[Router.scala 146:23]
  always @(posedge clock) begin
    switch_io_sel_REG_2_0_2_0 <= switch_allocator_io_switch_sel_2_0_2_0; // @[Router.scala 176:14]
    switch_io_sel_REG_2_0_1_0 <= switch_allocator_io_switch_sel_2_0_1_0; // @[Router.scala 176:14]
    switch_io_sel_REG_2_0_0_0 <= switch_allocator_io_switch_sel_2_0_0_0; // @[Router.scala 176:14]
    switch_io_sel_REG_1_0_2_0 <= switch_allocator_io_switch_sel_1_0_2_0; // @[Router.scala 176:14]
    switch_io_sel_REG_1_0_1_0 <= switch_allocator_io_switch_sel_1_0_1_0; // @[Router.scala 176:14]
    switch_io_sel_REG_1_0_0_0 <= switch_allocator_io_switch_sel_1_0_0_0; // @[Router.scala 176:14]
    switch_io_sel_REG_0_0_2_0 <= switch_allocator_io_switch_sel_0_0_2_0; // @[Router.scala 176:14]
    switch_io_sel_REG_0_0_1_0 <= switch_allocator_io_switch_sel_0_0_1_0; // @[Router.scala 176:14]
    switch_io_sel_REG_0_0_0_0 <= switch_allocator_io_switch_sel_0_0_0_0; // @[Router.scala 176:14]
    if (reset) begin // @[Router.scala 193:28]
      debug_tsc <= 64'h0; // @[Router.scala 193:28]
    end else begin
      debug_tsc <= _debug_tsc_T_1; // @[Router.scala 194:15]
    end
    if (reset) begin // @[Router.scala 195:31]
      debug_sample <= 64'h0; // @[Router.scala 195:31]
    end else if (debug_sample == _GEN_6) begin // @[Router.scala 198:47]
      debug_sample <= 64'h0; // @[Router.scala 198:62]
    end else begin
      debug_sample <= _debug_sample_T_1; // @[Router.scala 196:18]
    end
    if (reset) begin // @[Router.scala 201:29]
      util_ctr <= 64'h0; // @[Router.scala 201:29]
    end else begin
      util_ctr <= _util_ctr_T_1; // @[Router.scala 203:16]
    end
    if (reset) begin // @[Router.scala 202:26]
      fired <= 1'h0; // @[Router.scala 202:26]
    end else if (plusarg_reader_out != 20'h0 & _T_2 & fired) begin // @[Router.scala 205:81]
      fired <= auto_dest_nodes_in_0_flit_0_valid; // @[Router.scala 208:15]
    end else begin
      fired <= fired | auto_dest_nodes_in_0_flit_0_valid; // @[Router.scala 204:13]
    end
    if (reset) begin // @[Router.scala 201:29]
      util_ctr_1 <= 64'h0; // @[Router.scala 201:29]
    end else begin
      util_ctr_1 <= _util_ctr_T_3; // @[Router.scala 203:16]
    end
    if (reset) begin // @[Router.scala 202:26]
      fired_1 <= 1'h0; // @[Router.scala 202:26]
    end else if (plusarg_reader_out != 20'h0 & _T_2 & fired_1) begin // @[Router.scala 205:81]
      fired_1 <= auto_dest_nodes_in_1_flit_0_valid; // @[Router.scala 208:15]
    end else begin
      fired_1 <= fired_1 | auto_dest_nodes_in_1_flit_0_valid; // @[Router.scala 204:13]
    end
    if (reset) begin // @[Router.scala 201:29]
      util_ctr_2 <= 64'h0; // @[Router.scala 201:29]
    end else begin
      util_ctr_2 <= _util_ctr_T_5; // @[Router.scala 203:16]
    end
    if (reset) begin // @[Router.scala 202:26]
      fired_2 <= 1'h0; // @[Router.scala 202:26]
    end else if (plusarg_reader_out != 20'h0 & _T_2 & fired_2) begin // @[Router.scala 205:81]
      fired_2 <= _T_19; // @[Router.scala 208:15]
    end else begin
      fired_2 <= fired_2 | _T_19; // @[Router.scala 204:13]
    end
    if (reset) begin // @[Router.scala 201:29]
      util_ctr_3 <= 64'h0; // @[Router.scala 201:29]
    end else begin
      util_ctr_3 <= _util_ctr_T_7; // @[Router.scala 203:16]
    end
    if (reset) begin // @[Router.scala 202:26]
      fired_3 <= 1'h0; // @[Router.scala 202:26]
    end else if (plusarg_reader_out != 20'h0 & _T_2 & fired_3) begin // @[Router.scala 205:81]
      fired_3 <= x1_2_flit_valid; // @[Router.scala 208:15]
    end else begin
      fired_3 <= fired_3 | x1_2_flit_valid; // @[Router.scala 204:13]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8 & ~reset) begin
          $fwrite(32'h80000002,"nocsample %d 1 2 %d\n",debug_tsc,util_ctr); // @[Router.scala 207:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_16 & ~reset) begin
          $fwrite(32'h80000002,"nocsample %d 3 2 %d\n",debug_tsc,util_ctr_1); // @[Router.scala 207:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_25 & ~reset) begin
          $fwrite(32'h80000002,"nocsample %d i2 2 %d\n",debug_tsc,util_ctr_2); // @[Router.scala 207:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_34 & ~reset) begin
          $fwrite(32'h80000002,"nocsample %d 2 e2 %d\n",debug_tsc,util_ctr_3); // @[Router.scala 207:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  switch_io_sel_REG_2_0_2_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  switch_io_sel_REG_2_0_1_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  switch_io_sel_REG_2_0_0_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  switch_io_sel_REG_1_0_2_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  switch_io_sel_REG_1_0_1_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  switch_io_sel_REG_1_0_0_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  switch_io_sel_REG_0_0_2_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  switch_io_sel_REG_0_0_1_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  switch_io_sel_REG_0_0_0_0 = _RAND_8[0:0];
  _RAND_9 = {2{`RANDOM}};
  debug_tsc = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  debug_sample = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  util_ctr = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  fired = _RAND_12[0:0];
  _RAND_13 = {2{`RANDOM}};
  util_ctr_1 = _RAND_13[63:0];
  _RAND_14 = {1{`RANDOM}};
  fired_1 = _RAND_14[0:0];
  _RAND_15 = {2{`RANDOM}};
  util_ctr_2 = _RAND_15[63:0];
  _RAND_16 = {1{`RANDOM}};
  fired_2 = _RAND_16[0:0];
  _RAND_17 = {2{`RANDOM}};
  util_ctr_3 = _RAND_17[63:0];
  _RAND_18 = {1{`RANDOM}};
  fired_3 = _RAND_18[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ClockSinkDomain_2(
  output [1:0]  auto_routers_debug_out_va_stall_0,
  output [1:0]  auto_routers_debug_out_va_stall_1,
  output [1:0]  auto_routers_debug_out_sa_stall_0,
  output [1:0]  auto_routers_debug_out_sa_stall_1,
  output        auto_routers_egress_nodes_out_flit_valid,
  output        auto_routers_egress_nodes_out_flit_bits_head,
  output        auto_routers_egress_nodes_out_flit_bits_tail,
  output [63:0] auto_routers_egress_nodes_out_flit_bits_payload,
  output [1:0]  auto_routers_egress_nodes_out_flit_bits_ingress_id,
  output        auto_routers_ingress_nodes_in_flit_ready,
  input         auto_routers_ingress_nodes_in_flit_valid,
  input         auto_routers_ingress_nodes_in_flit_bits_head,
  input         auto_routers_ingress_nodes_in_flit_bits_tail,
  input  [63:0] auto_routers_ingress_nodes_in_flit_bits_payload,
  input  [1:0]  auto_routers_ingress_nodes_in_flit_bits_egress_id,
  output        auto_routers_source_nodes_out_1_flit_0_valid,
  output        auto_routers_source_nodes_out_1_flit_0_bits_head,
  output        auto_routers_source_nodes_out_1_flit_0_bits_tail,
  output [63:0] auto_routers_source_nodes_out_1_flit_0_bits_payload,
  output [1:0]  auto_routers_source_nodes_out_1_flit_0_bits_flow_ingress_node,
  output [1:0]  auto_routers_source_nodes_out_1_flit_0_bits_flow_egress_node,
  output [1:0]  auto_routers_source_nodes_out_1_flit_0_bits_virt_channel_id,
  input  [3:0]  auto_routers_source_nodes_out_1_credit_return,
  input  [3:0]  auto_routers_source_nodes_out_1_vc_free,
  output        auto_routers_source_nodes_out_0_flit_0_valid,
  output        auto_routers_source_nodes_out_0_flit_0_bits_head,
  output        auto_routers_source_nodes_out_0_flit_0_bits_tail,
  output [63:0] auto_routers_source_nodes_out_0_flit_0_bits_payload,
  output [1:0]  auto_routers_source_nodes_out_0_flit_0_bits_flow_ingress_node,
  output [1:0]  auto_routers_source_nodes_out_0_flit_0_bits_flow_egress_node,
  output [1:0]  auto_routers_source_nodes_out_0_flit_0_bits_virt_channel_id,
  input  [3:0]  auto_routers_source_nodes_out_0_credit_return,
  input  [3:0]  auto_routers_source_nodes_out_0_vc_free,
  input         auto_routers_dest_nodes_in_1_flit_0_valid,
  input         auto_routers_dest_nodes_in_1_flit_0_bits_head,
  input         auto_routers_dest_nodes_in_1_flit_0_bits_tail,
  input  [63:0] auto_routers_dest_nodes_in_1_flit_0_bits_payload,
  input  [1:0]  auto_routers_dest_nodes_in_1_flit_0_bits_flow_ingress_node,
  input  [1:0]  auto_routers_dest_nodes_in_1_flit_0_bits_flow_egress_node,
  input  [1:0]  auto_routers_dest_nodes_in_1_flit_0_bits_virt_channel_id,
  output [3:0]  auto_routers_dest_nodes_in_1_credit_return,
  output [3:0]  auto_routers_dest_nodes_in_1_vc_free,
  input         auto_routers_dest_nodes_in_0_flit_0_valid,
  input         auto_routers_dest_nodes_in_0_flit_0_bits_head,
  input         auto_routers_dest_nodes_in_0_flit_0_bits_tail,
  input  [63:0] auto_routers_dest_nodes_in_0_flit_0_bits_payload,
  input  [1:0]  auto_routers_dest_nodes_in_0_flit_0_bits_flow_ingress_node,
  input  [1:0]  auto_routers_dest_nodes_in_0_flit_0_bits_flow_egress_node,
  input  [1:0]  auto_routers_dest_nodes_in_0_flit_0_bits_virt_channel_id,
  output [3:0]  auto_routers_dest_nodes_in_0_credit_return,
  output [3:0]  auto_routers_dest_nodes_in_0_vc_free,
  input         auto_clock_in_clock,
  input         auto_clock_in_reset
);
  wire  routers_clock; // @[NoC.scala 64:22]
  wire  routers_reset; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_debug_out_va_stall_0; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_debug_out_va_stall_1; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_debug_out_sa_stall_0; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_debug_out_sa_stall_1; // @[NoC.scala 64:22]
  wire  routers_auto_egress_nodes_out_flit_valid; // @[NoC.scala 64:22]
  wire  routers_auto_egress_nodes_out_flit_bits_head; // @[NoC.scala 64:22]
  wire  routers_auto_egress_nodes_out_flit_bits_tail; // @[NoC.scala 64:22]
  wire [63:0] routers_auto_egress_nodes_out_flit_bits_payload; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_egress_nodes_out_flit_bits_ingress_id; // @[NoC.scala 64:22]
  wire  routers_auto_ingress_nodes_in_flit_ready; // @[NoC.scala 64:22]
  wire  routers_auto_ingress_nodes_in_flit_valid; // @[NoC.scala 64:22]
  wire  routers_auto_ingress_nodes_in_flit_bits_head; // @[NoC.scala 64:22]
  wire  routers_auto_ingress_nodes_in_flit_bits_tail; // @[NoC.scala 64:22]
  wire [63:0] routers_auto_ingress_nodes_in_flit_bits_payload; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_ingress_nodes_in_flit_bits_egress_id; // @[NoC.scala 64:22]
  wire  routers_auto_source_nodes_out_1_flit_0_valid; // @[NoC.scala 64:22]
  wire  routers_auto_source_nodes_out_1_flit_0_bits_head; // @[NoC.scala 64:22]
  wire  routers_auto_source_nodes_out_1_flit_0_bits_tail; // @[NoC.scala 64:22]
  wire [63:0] routers_auto_source_nodes_out_1_flit_0_bits_payload; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_source_nodes_out_1_flit_0_bits_flow_ingress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_source_nodes_out_1_flit_0_bits_flow_egress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_source_nodes_out_1_flit_0_bits_virt_channel_id; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_source_nodes_out_1_credit_return; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_source_nodes_out_1_vc_free; // @[NoC.scala 64:22]
  wire  routers_auto_source_nodes_out_0_flit_0_valid; // @[NoC.scala 64:22]
  wire  routers_auto_source_nodes_out_0_flit_0_bits_head; // @[NoC.scala 64:22]
  wire  routers_auto_source_nodes_out_0_flit_0_bits_tail; // @[NoC.scala 64:22]
  wire [63:0] routers_auto_source_nodes_out_0_flit_0_bits_payload; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_source_nodes_out_0_flit_0_bits_flow_ingress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_source_nodes_out_0_flit_0_bits_flow_egress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_source_nodes_out_0_flit_0_bits_virt_channel_id; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_source_nodes_out_0_credit_return; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_source_nodes_out_0_vc_free; // @[NoC.scala 64:22]
  wire  routers_auto_dest_nodes_in_1_flit_0_valid; // @[NoC.scala 64:22]
  wire  routers_auto_dest_nodes_in_1_flit_0_bits_head; // @[NoC.scala 64:22]
  wire  routers_auto_dest_nodes_in_1_flit_0_bits_tail; // @[NoC.scala 64:22]
  wire [63:0] routers_auto_dest_nodes_in_1_flit_0_bits_payload; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_dest_nodes_in_1_flit_0_bits_flow_ingress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_dest_nodes_in_1_flit_0_bits_flow_egress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_dest_nodes_in_1_flit_0_bits_virt_channel_id; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_dest_nodes_in_1_credit_return; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_dest_nodes_in_1_vc_free; // @[NoC.scala 64:22]
  wire  routers_auto_dest_nodes_in_0_flit_0_valid; // @[NoC.scala 64:22]
  wire  routers_auto_dest_nodes_in_0_flit_0_bits_head; // @[NoC.scala 64:22]
  wire  routers_auto_dest_nodes_in_0_flit_0_bits_tail; // @[NoC.scala 64:22]
  wire [63:0] routers_auto_dest_nodes_in_0_flit_0_bits_payload; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_dest_nodes_in_0_flit_0_bits_flow_ingress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_dest_nodes_in_0_flit_0_bits_flow_egress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_dest_nodes_in_0_flit_0_bits_virt_channel_id; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_dest_nodes_in_0_credit_return; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_dest_nodes_in_0_vc_free; // @[NoC.scala 64:22]
  Router_2 routers ( // @[NoC.scala 64:22]
    .clock(routers_clock),
    .reset(routers_reset),
    .auto_debug_out_va_stall_0(routers_auto_debug_out_va_stall_0),
    .auto_debug_out_va_stall_1(routers_auto_debug_out_va_stall_1),
    .auto_debug_out_sa_stall_0(routers_auto_debug_out_sa_stall_0),
    .auto_debug_out_sa_stall_1(routers_auto_debug_out_sa_stall_1),
    .auto_egress_nodes_out_flit_valid(routers_auto_egress_nodes_out_flit_valid),
    .auto_egress_nodes_out_flit_bits_head(routers_auto_egress_nodes_out_flit_bits_head),
    .auto_egress_nodes_out_flit_bits_tail(routers_auto_egress_nodes_out_flit_bits_tail),
    .auto_egress_nodes_out_flit_bits_payload(routers_auto_egress_nodes_out_flit_bits_payload),
    .auto_egress_nodes_out_flit_bits_ingress_id(routers_auto_egress_nodes_out_flit_bits_ingress_id),
    .auto_ingress_nodes_in_flit_ready(routers_auto_ingress_nodes_in_flit_ready),
    .auto_ingress_nodes_in_flit_valid(routers_auto_ingress_nodes_in_flit_valid),
    .auto_ingress_nodes_in_flit_bits_head(routers_auto_ingress_nodes_in_flit_bits_head),
    .auto_ingress_nodes_in_flit_bits_tail(routers_auto_ingress_nodes_in_flit_bits_tail),
    .auto_ingress_nodes_in_flit_bits_payload(routers_auto_ingress_nodes_in_flit_bits_payload),
    .auto_ingress_nodes_in_flit_bits_egress_id(routers_auto_ingress_nodes_in_flit_bits_egress_id),
    .auto_source_nodes_out_1_flit_0_valid(routers_auto_source_nodes_out_1_flit_0_valid),
    .auto_source_nodes_out_1_flit_0_bits_head(routers_auto_source_nodes_out_1_flit_0_bits_head),
    .auto_source_nodes_out_1_flit_0_bits_tail(routers_auto_source_nodes_out_1_flit_0_bits_tail),
    .auto_source_nodes_out_1_flit_0_bits_payload(routers_auto_source_nodes_out_1_flit_0_bits_payload),
    .auto_source_nodes_out_1_flit_0_bits_flow_ingress_node(routers_auto_source_nodes_out_1_flit_0_bits_flow_ingress_node
      ),
    .auto_source_nodes_out_1_flit_0_bits_flow_egress_node(routers_auto_source_nodes_out_1_flit_0_bits_flow_egress_node),
    .auto_source_nodes_out_1_flit_0_bits_virt_channel_id(routers_auto_source_nodes_out_1_flit_0_bits_virt_channel_id),
    .auto_source_nodes_out_1_credit_return(routers_auto_source_nodes_out_1_credit_return),
    .auto_source_nodes_out_1_vc_free(routers_auto_source_nodes_out_1_vc_free),
    .auto_source_nodes_out_0_flit_0_valid(routers_auto_source_nodes_out_0_flit_0_valid),
    .auto_source_nodes_out_0_flit_0_bits_head(routers_auto_source_nodes_out_0_flit_0_bits_head),
    .auto_source_nodes_out_0_flit_0_bits_tail(routers_auto_source_nodes_out_0_flit_0_bits_tail),
    .auto_source_nodes_out_0_flit_0_bits_payload(routers_auto_source_nodes_out_0_flit_0_bits_payload),
    .auto_source_nodes_out_0_flit_0_bits_flow_ingress_node(routers_auto_source_nodes_out_0_flit_0_bits_flow_ingress_node
      ),
    .auto_source_nodes_out_0_flit_0_bits_flow_egress_node(routers_auto_source_nodes_out_0_flit_0_bits_flow_egress_node),
    .auto_source_nodes_out_0_flit_0_bits_virt_channel_id(routers_auto_source_nodes_out_0_flit_0_bits_virt_channel_id),
    .auto_source_nodes_out_0_credit_return(routers_auto_source_nodes_out_0_credit_return),
    .auto_source_nodes_out_0_vc_free(routers_auto_source_nodes_out_0_vc_free),
    .auto_dest_nodes_in_1_flit_0_valid(routers_auto_dest_nodes_in_1_flit_0_valid),
    .auto_dest_nodes_in_1_flit_0_bits_head(routers_auto_dest_nodes_in_1_flit_0_bits_head),
    .auto_dest_nodes_in_1_flit_0_bits_tail(routers_auto_dest_nodes_in_1_flit_0_bits_tail),
    .auto_dest_nodes_in_1_flit_0_bits_payload(routers_auto_dest_nodes_in_1_flit_0_bits_payload),
    .auto_dest_nodes_in_1_flit_0_bits_flow_ingress_node(routers_auto_dest_nodes_in_1_flit_0_bits_flow_ingress_node),
    .auto_dest_nodes_in_1_flit_0_bits_flow_egress_node(routers_auto_dest_nodes_in_1_flit_0_bits_flow_egress_node),
    .auto_dest_nodes_in_1_flit_0_bits_virt_channel_id(routers_auto_dest_nodes_in_1_flit_0_bits_virt_channel_id),
    .auto_dest_nodes_in_1_credit_return(routers_auto_dest_nodes_in_1_credit_return),
    .auto_dest_nodes_in_1_vc_free(routers_auto_dest_nodes_in_1_vc_free),
    .auto_dest_nodes_in_0_flit_0_valid(routers_auto_dest_nodes_in_0_flit_0_valid),
    .auto_dest_nodes_in_0_flit_0_bits_head(routers_auto_dest_nodes_in_0_flit_0_bits_head),
    .auto_dest_nodes_in_0_flit_0_bits_tail(routers_auto_dest_nodes_in_0_flit_0_bits_tail),
    .auto_dest_nodes_in_0_flit_0_bits_payload(routers_auto_dest_nodes_in_0_flit_0_bits_payload),
    .auto_dest_nodes_in_0_flit_0_bits_flow_ingress_node(routers_auto_dest_nodes_in_0_flit_0_bits_flow_ingress_node),
    .auto_dest_nodes_in_0_flit_0_bits_flow_egress_node(routers_auto_dest_nodes_in_0_flit_0_bits_flow_egress_node),
    .auto_dest_nodes_in_0_flit_0_bits_virt_channel_id(routers_auto_dest_nodes_in_0_flit_0_bits_virt_channel_id),
    .auto_dest_nodes_in_0_credit_return(routers_auto_dest_nodes_in_0_credit_return),
    .auto_dest_nodes_in_0_vc_free(routers_auto_dest_nodes_in_0_vc_free)
  );
  assign auto_routers_debug_out_va_stall_0 = routers_auto_debug_out_va_stall_0; // @[LazyModule.scala 368:12]
  assign auto_routers_debug_out_va_stall_1 = routers_auto_debug_out_va_stall_1; // @[LazyModule.scala 368:12]
  assign auto_routers_debug_out_sa_stall_0 = routers_auto_debug_out_sa_stall_0; // @[LazyModule.scala 368:12]
  assign auto_routers_debug_out_sa_stall_1 = routers_auto_debug_out_sa_stall_1; // @[LazyModule.scala 368:12]
  assign auto_routers_egress_nodes_out_flit_valid = routers_auto_egress_nodes_out_flit_valid; // @[LazyModule.scala 368:12]
  assign auto_routers_egress_nodes_out_flit_bits_head = routers_auto_egress_nodes_out_flit_bits_head; // @[LazyModule.scala 368:12]
  assign auto_routers_egress_nodes_out_flit_bits_tail = routers_auto_egress_nodes_out_flit_bits_tail; // @[LazyModule.scala 368:12]
  assign auto_routers_egress_nodes_out_flit_bits_payload = routers_auto_egress_nodes_out_flit_bits_payload; // @[LazyModule.scala 368:12]
  assign auto_routers_egress_nodes_out_flit_bits_ingress_id = routers_auto_egress_nodes_out_flit_bits_ingress_id; // @[LazyModule.scala 368:12]
  assign auto_routers_ingress_nodes_in_flit_ready = routers_auto_ingress_nodes_in_flit_ready; // @[LazyModule.scala 366:16]
  assign auto_routers_source_nodes_out_1_flit_0_valid = routers_auto_source_nodes_out_1_flit_0_valid; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_1_flit_0_bits_head = routers_auto_source_nodes_out_1_flit_0_bits_head; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_1_flit_0_bits_tail = routers_auto_source_nodes_out_1_flit_0_bits_tail; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_1_flit_0_bits_payload = routers_auto_source_nodes_out_1_flit_0_bits_payload; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_1_flit_0_bits_flow_ingress_node =
    routers_auto_source_nodes_out_1_flit_0_bits_flow_ingress_node; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_1_flit_0_bits_flow_egress_node =
    routers_auto_source_nodes_out_1_flit_0_bits_flow_egress_node; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_1_flit_0_bits_virt_channel_id =
    routers_auto_source_nodes_out_1_flit_0_bits_virt_channel_id; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_0_flit_0_valid = routers_auto_source_nodes_out_0_flit_0_valid; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_0_flit_0_bits_head = routers_auto_source_nodes_out_0_flit_0_bits_head; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_0_flit_0_bits_tail = routers_auto_source_nodes_out_0_flit_0_bits_tail; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_0_flit_0_bits_payload = routers_auto_source_nodes_out_0_flit_0_bits_payload; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_0_flit_0_bits_flow_ingress_node =
    routers_auto_source_nodes_out_0_flit_0_bits_flow_ingress_node; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_0_flit_0_bits_flow_egress_node =
    routers_auto_source_nodes_out_0_flit_0_bits_flow_egress_node; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_0_flit_0_bits_virt_channel_id =
    routers_auto_source_nodes_out_0_flit_0_bits_virt_channel_id; // @[LazyModule.scala 368:12]
  assign auto_routers_dest_nodes_in_1_credit_return = routers_auto_dest_nodes_in_1_credit_return; // @[LazyModule.scala 366:16]
  assign auto_routers_dest_nodes_in_1_vc_free = routers_auto_dest_nodes_in_1_vc_free; // @[LazyModule.scala 366:16]
  assign auto_routers_dest_nodes_in_0_credit_return = routers_auto_dest_nodes_in_0_credit_return; // @[LazyModule.scala 366:16]
  assign auto_routers_dest_nodes_in_0_vc_free = routers_auto_dest_nodes_in_0_vc_free; // @[LazyModule.scala 366:16]
  assign routers_clock = auto_clock_in_clock; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign routers_reset = auto_clock_in_reset; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign routers_auto_ingress_nodes_in_flit_valid = auto_routers_ingress_nodes_in_flit_valid; // @[LazyModule.scala 366:16]
  assign routers_auto_ingress_nodes_in_flit_bits_head = auto_routers_ingress_nodes_in_flit_bits_head; // @[LazyModule.scala 366:16]
  assign routers_auto_ingress_nodes_in_flit_bits_tail = auto_routers_ingress_nodes_in_flit_bits_tail; // @[LazyModule.scala 366:16]
  assign routers_auto_ingress_nodes_in_flit_bits_payload = auto_routers_ingress_nodes_in_flit_bits_payload; // @[LazyModule.scala 366:16]
  assign routers_auto_ingress_nodes_in_flit_bits_egress_id = auto_routers_ingress_nodes_in_flit_bits_egress_id; // @[LazyModule.scala 366:16]
  assign routers_auto_source_nodes_out_1_credit_return = auto_routers_source_nodes_out_1_credit_return; // @[LazyModule.scala 368:12]
  assign routers_auto_source_nodes_out_1_vc_free = auto_routers_source_nodes_out_1_vc_free; // @[LazyModule.scala 368:12]
  assign routers_auto_source_nodes_out_0_credit_return = auto_routers_source_nodes_out_0_credit_return; // @[LazyModule.scala 368:12]
  assign routers_auto_source_nodes_out_0_vc_free = auto_routers_source_nodes_out_0_vc_free; // @[LazyModule.scala 368:12]
  assign routers_auto_dest_nodes_in_1_flit_0_valid = auto_routers_dest_nodes_in_1_flit_0_valid; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_1_flit_0_bits_head = auto_routers_dest_nodes_in_1_flit_0_bits_head; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_1_flit_0_bits_tail = auto_routers_dest_nodes_in_1_flit_0_bits_tail; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_1_flit_0_bits_payload = auto_routers_dest_nodes_in_1_flit_0_bits_payload; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_1_flit_0_bits_flow_ingress_node =
    auto_routers_dest_nodes_in_1_flit_0_bits_flow_ingress_node; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_1_flit_0_bits_flow_egress_node =
    auto_routers_dest_nodes_in_1_flit_0_bits_flow_egress_node; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_1_flit_0_bits_virt_channel_id =
    auto_routers_dest_nodes_in_1_flit_0_bits_virt_channel_id; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_0_flit_0_valid = auto_routers_dest_nodes_in_0_flit_0_valid; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_0_flit_0_bits_head = auto_routers_dest_nodes_in_0_flit_0_bits_head; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_0_flit_0_bits_tail = auto_routers_dest_nodes_in_0_flit_0_bits_tail; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_0_flit_0_bits_payload = auto_routers_dest_nodes_in_0_flit_0_bits_payload; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_0_flit_0_bits_flow_ingress_node =
    auto_routers_dest_nodes_in_0_flit_0_bits_flow_ingress_node; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_0_flit_0_bits_flow_egress_node =
    auto_routers_dest_nodes_in_0_flit_0_bits_flow_egress_node; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_0_flit_0_bits_virt_channel_id =
    auto_routers_dest_nodes_in_0_flit_0_bits_virt_channel_id; // @[LazyModule.scala 366:16]
endmodule
module NoCMonitor_6(
  input        clock,
  input        reset,
  input        io_in_flit_0_valid,
  input        io_in_flit_0_bits_head,
  input        io_in_flit_0_bits_tail,
  input  [1:0] io_in_flit_0_bits_flow_ingress_node,
  input  [1:0] io_in_flit_0_bits_flow_egress_node,
  input  [1:0] io_in_flit_0_bits_virt_channel_id
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg  in_flight_0; // @[Monitor.scala 16:26]
  reg  in_flight_1; // @[Monitor.scala 16:26]
  reg  in_flight_2; // @[Monitor.scala 16:26]
  reg  in_flight_3; // @[Monitor.scala 16:26]
  wire  _GEN_0 = 2'h0 == io_in_flit_0_bits_virt_channel_id | in_flight_0; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_1 = 2'h1 == io_in_flit_0_bits_virt_channel_id | in_flight_1; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_2 = 2'h2 == io_in_flit_0_bits_virt_channel_id | in_flight_2; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_3 = 2'h3 == io_in_flit_0_bits_virt_channel_id | in_flight_3; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_5 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? in_flight_1 : in_flight_0; // @[Monitor.scala 22:{17,17}]
  wire  _GEN_6 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? in_flight_2 : _GEN_5; // @[Monitor.scala 22:{17,17}]
  wire  _GEN_7 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? in_flight_3 : _GEN_6; // @[Monitor.scala 22:{17,17}]
  wire  _T_2 = ~reset; // @[Monitor.scala 22:16]
  wire  _GEN_8 = io_in_flit_0_bits_head ? _GEN_0 : in_flight_0; // @[Monitor.scala 16:26 20:29]
  wire  _GEN_9 = io_in_flit_0_bits_head ? _GEN_1 : in_flight_1; // @[Monitor.scala 16:26 20:29]
  wire  _GEN_10 = io_in_flit_0_bits_head ? _GEN_2 : in_flight_2; // @[Monitor.scala 16:26 20:29]
  wire  _GEN_11 = io_in_flit_0_bits_head ? _GEN_3 : in_flight_3; // @[Monitor.scala 16:26 20:29]
  wire  _T_4 = io_in_flit_0_valid & io_in_flit_0_bits_head; // @[Monitor.scala 29:22]
  wire  _T_7 = io_in_flit_0_bits_flow_egress_node == 2'h3; // @[Types.scala 54:21]
  wire  _T_8 = io_in_flit_0_bits_flow_ingress_node == 2'h1 & _T_7; // @[Types.scala 53:39]
  wire  _T_19 = io_in_flit_0_bits_flow_egress_node == 2'h2; // @[Types.scala 54:21]
  wire  _T_20 = io_in_flit_0_bits_flow_ingress_node == 2'h0 & _T_19; // @[Types.scala 53:39]
  wire  _T_27 = io_in_flit_0_bits_flow_ingress_node == 2'h0 & _T_7; // @[Types.scala 53:39]
  wire  _T_39 = _T_20 | _T_27; // @[package.scala 73:59]
  wire  _T_40 = _T_20 | _T_27 | _T_8; // @[package.scala 73:59]
  wire  _GEN_29 = _T_4 & ~reset; // @[Monitor.scala 22:16]
  always @(posedge clock) begin
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_0 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h0 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_0 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_0 <= _GEN_8;
        end
      end else begin
        in_flight_0 <= _GEN_8;
      end
    end
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_1 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h1 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_1 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_1 <= _GEN_9;
        end
      end else begin
        in_flight_1 <= _GEN_9;
      end
    end
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_2 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h2 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_2 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_2 <= _GEN_10;
        end
      end else begin
        in_flight_2 <= _GEN_10;
      end
    end
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_3 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h3 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_3 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_3 <= _GEN_11;
        end
      end else begin
        in_flight_3 <= _GEN_11;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4 & ~reset & ~(~_GEN_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed: Flit head/tail sequencing is broken\n    at Monitor.scala:22 assert (!in_flight(flit.bits.virt_channel_id), \"Flit head/tail sequencing is broken\")\n"
            ); // @[Monitor.scala 22:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h0 | _T_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h1 | _T_40)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h2 | _T_40)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h3 | _T_39)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  in_flight_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  in_flight_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  in_flight_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  in_flight_3 = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (_T_4 & ~reset) begin
      assert(~_GEN_7); // @[Monitor.scala 22:16]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h0 | _T_8); // @[Monitor.scala 32:17]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h1 | _T_40); // @[Monitor.scala 32:17]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h2 | _T_40); // @[Monitor.scala 32:17]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h3 | _T_39); // @[Monitor.scala 32:17]
    end
  end
endmodule
module NoCMonitor_7(
  input        clock,
  input        reset,
  input        io_in_flit_0_valid,
  input        io_in_flit_0_bits_head,
  input        io_in_flit_0_bits_tail,
  input  [1:0] io_in_flit_0_bits_flow_ingress_node,
  input  [1:0] io_in_flit_0_bits_flow_egress_node,
  input  [1:0] io_in_flit_0_bits_virt_channel_id
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg  in_flight_0; // @[Monitor.scala 16:26]
  reg  in_flight_1; // @[Monitor.scala 16:26]
  reg  in_flight_2; // @[Monitor.scala 16:26]
  reg  in_flight_3; // @[Monitor.scala 16:26]
  wire  _GEN_0 = 2'h0 == io_in_flit_0_bits_virt_channel_id | in_flight_0; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_1 = 2'h1 == io_in_flit_0_bits_virt_channel_id | in_flight_1; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_2 = 2'h2 == io_in_flit_0_bits_virt_channel_id | in_flight_2; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_3 = 2'h3 == io_in_flit_0_bits_virt_channel_id | in_flight_3; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_5 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? in_flight_1 : in_flight_0; // @[Monitor.scala 22:{17,17}]
  wire  _GEN_6 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? in_flight_2 : _GEN_5; // @[Monitor.scala 22:{17,17}]
  wire  _GEN_7 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? in_flight_3 : _GEN_6; // @[Monitor.scala 22:{17,17}]
  wire  _T_2 = ~reset; // @[Monitor.scala 22:16]
  wire  _GEN_8 = io_in_flit_0_bits_head ? _GEN_0 : in_flight_0; // @[Monitor.scala 16:26 20:29]
  wire  _GEN_9 = io_in_flit_0_bits_head ? _GEN_1 : in_flight_1; // @[Monitor.scala 16:26 20:29]
  wire  _GEN_10 = io_in_flit_0_bits_head ? _GEN_2 : in_flight_2; // @[Monitor.scala 16:26 20:29]
  wire  _GEN_11 = io_in_flit_0_bits_head ? _GEN_3 : in_flight_3; // @[Monitor.scala 16:26 20:29]
  wire  _T_4 = io_in_flit_0_valid & io_in_flit_0_bits_head; // @[Monitor.scala 29:22]
  wire  _T_7 = io_in_flit_0_bits_flow_egress_node == 2'h3; // @[Types.scala 54:21]
  wire  _T_8 = io_in_flit_0_bits_flow_ingress_node == 2'h1 & _T_7; // @[Types.scala 53:39]
  wire  _T_26 = io_in_flit_0_bits_flow_egress_node == 2'h0; // @[Types.scala 54:21]
  wire  _T_27 = io_in_flit_0_bits_flow_ingress_node == 2'h2 & _T_26; // @[Types.scala 53:39]
  wire  _T_34 = io_in_flit_0_bits_flow_ingress_node == 2'h2 & _T_7; // @[Types.scala 53:39]
  wire  _T_40 = _T_8 | _T_27 | _T_34; // @[package.scala 73:59]
  wire  _GEN_29 = _T_4 & ~reset; // @[Monitor.scala 22:16]
  always @(posedge clock) begin
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_0 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h0 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_0 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_0 <= _GEN_8;
        end
      end else begin
        in_flight_0 <= _GEN_8;
      end
    end
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_1 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h1 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_1 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_1 <= _GEN_9;
        end
      end else begin
        in_flight_1 <= _GEN_9;
      end
    end
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_2 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h2 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_2 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_2 <= _GEN_10;
        end
      end else begin
        in_flight_2 <= _GEN_10;
      end
    end
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_3 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h3 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_3 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_3 <= _GEN_11;
        end
      end else begin
        in_flight_3 <= _GEN_11;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4 & ~reset & ~(~_GEN_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed: Flit head/tail sequencing is broken\n    at Monitor.scala:22 assert (!in_flight(flit.bits.virt_channel_id), \"Flit head/tail sequencing is broken\")\n"
            ); // @[Monitor.scala 22:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h0 | _T_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h1 | _T_40)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h2 | _T_40)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h3 | _T_40)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  in_flight_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  in_flight_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  in_flight_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  in_flight_3 = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (_T_4 & ~reset) begin
      assert(~_GEN_7); // @[Monitor.scala 22:16]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h0 | _T_8); // @[Monitor.scala 32:17]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h1 | _T_40); // @[Monitor.scala 32:17]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h2 | _T_40); // @[Monitor.scala 32:17]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h3 | _T_40); // @[Monitor.scala 32:17]
    end
  end
endmodule
module InputUnit_6(
  input         clock,
  input         reset,
  output        io_router_req_valid,
  output [1:0]  io_router_req_bits_src_virt_id,
  output [1:0]  io_router_req_bits_flow_ingress_node,
  output [1:0]  io_router_req_bits_flow_egress_node,
  input         io_router_resp_vc_sel_1_0,
  input         io_router_resp_vc_sel_1_1,
  input         io_router_resp_vc_sel_1_2,
  input         io_router_resp_vc_sel_1_3,
  input         io_router_resp_vc_sel_0_0,
  input         io_router_resp_vc_sel_0_1,
  input         io_router_resp_vc_sel_0_2,
  input         io_vcalloc_req_ready,
  output        io_vcalloc_req_valid,
  output        io_vcalloc_req_bits_vc_sel_2_0,
  output        io_vcalloc_req_bits_vc_sel_1_0,
  output        io_vcalloc_req_bits_vc_sel_1_1,
  output        io_vcalloc_req_bits_vc_sel_1_2,
  output        io_vcalloc_req_bits_vc_sel_1_3,
  output        io_vcalloc_req_bits_vc_sel_0_0,
  output        io_vcalloc_req_bits_vc_sel_0_1,
  output        io_vcalloc_req_bits_vc_sel_0_2,
  input         io_vcalloc_resp_vc_sel_2_0,
  input         io_vcalloc_resp_vc_sel_1_0,
  input         io_vcalloc_resp_vc_sel_1_1,
  input         io_vcalloc_resp_vc_sel_1_2,
  input         io_vcalloc_resp_vc_sel_1_3,
  input         io_vcalloc_resp_vc_sel_0_0,
  input         io_vcalloc_resp_vc_sel_0_1,
  input         io_vcalloc_resp_vc_sel_0_2,
  input         io_out_credit_available_2_0,
  input         io_out_credit_available_1_0,
  input         io_out_credit_available_1_1,
  input         io_out_credit_available_1_2,
  input         io_out_credit_available_1_3,
  input         io_out_credit_available_0_0,
  input         io_out_credit_available_0_1,
  input         io_out_credit_available_0_2,
  input         io_out_credit_available_0_3,
  input         io_salloc_req_0_ready,
  output        io_salloc_req_0_valid,
  output        io_salloc_req_0_bits_vc_sel_2_0,
  output        io_salloc_req_0_bits_vc_sel_1_0,
  output        io_salloc_req_0_bits_vc_sel_1_1,
  output        io_salloc_req_0_bits_vc_sel_1_2,
  output        io_salloc_req_0_bits_vc_sel_1_3,
  output        io_salloc_req_0_bits_vc_sel_0_0,
  output        io_salloc_req_0_bits_vc_sel_0_1,
  output        io_salloc_req_0_bits_vc_sel_0_2,
  output        io_salloc_req_0_bits_vc_sel_0_3,
  output        io_salloc_req_0_bits_tail,
  output        io_out_0_valid,
  output        io_out_0_bits_flit_head,
  output        io_out_0_bits_flit_tail,
  output [63:0] io_out_0_bits_flit_payload,
  output [1:0]  io_out_0_bits_flit_flow_ingress_node,
  output [1:0]  io_out_0_bits_flit_flow_egress_node,
  output [1:0]  io_out_0_bits_out_virt_channel,
  output [1:0]  io_debug_va_stall,
  output [1:0]  io_debug_sa_stall,
  input         io_in_flit_0_valid,
  input         io_in_flit_0_bits_head,
  input         io_in_flit_0_bits_tail,
  input  [63:0] io_in_flit_0_bits_payload,
  input  [1:0]  io_in_flit_0_bits_flow_ingress_node,
  input  [1:0]  io_in_flit_0_bits_flow_egress_node,
  input  [1:0]  io_in_flit_0_bits_virt_channel_id,
  output [3:0]  io_in_credit_return,
  output [3:0]  io_in_vc_free
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
`endif // RANDOMIZE_REG_INIT
  wire  input_buffer_clock; // @[InputUnit.scala 180:28]
  wire  input_buffer_reset; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_enq_0_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_enq_0_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_enq_0_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_enq_0_bits_payload; // @[InputUnit.scala 180:28]
  wire [1:0] input_buffer_io_enq_0_bits_virt_channel_id; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_0_ready; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_0_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_0_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_0_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_deq_0_bits_payload; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_ready; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_deq_1_bits_payload; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_ready; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_deq_2_bits_payload; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_3_ready; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_3_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_3_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_3_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_deq_3_bits_payload; // @[InputUnit.scala 180:28]
  wire  route_arbiter_io_in_0_valid; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_0_bits_flow_ingress_node; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_0_bits_flow_egress_node; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_1_ready; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_1_valid; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_1_bits_flow_ingress_node; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_1_bits_flow_egress_node; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_2_ready; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_2_valid; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_2_bits_flow_ingress_node; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_2_bits_flow_egress_node; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_3_ready; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_3_valid; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_3_bits_flow_ingress_node; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_3_bits_flow_egress_node; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_out_valid; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_out_bits_src_virt_id; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_out_bits_flow_ingress_node; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_out_bits_flow_egress_node; // @[InputUnit.scala 186:29]
  wire  salloc_arb_clock; // @[InputUnit.scala 279:26]
  wire  salloc_arb_reset; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_bits_vc_sel_2_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_bits_vc_sel_1_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_bits_tail; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_vc_sel_2_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_vc_sel_1_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_vc_sel_1_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_vc_sel_0_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_tail; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_2_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_1_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_1_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_1_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_0_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_0_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_tail; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_2_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_1_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_1_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_1_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_1_3; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_0_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_0_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_0_3; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_tail; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_2_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_1_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_1_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_1_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_1_3; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_0_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_0_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_0_3; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_tail; // @[InputUnit.scala 279:26]
  wire [3:0] salloc_arb_io_chosen_oh_0; // @[InputUnit.scala 279:26]
  reg [2:0] states_0_g; // @[InputUnit.scala 191:19]
  reg  states_0_vc_sel_2_0; // @[InputUnit.scala 191:19]
  reg  states_0_vc_sel_1_0; // @[InputUnit.scala 191:19]
  reg  states_0_vc_sel_0_0; // @[InputUnit.scala 191:19]
  reg [1:0] states_0_flow_ingress_node; // @[InputUnit.scala 191:19]
  reg [1:0] states_0_flow_egress_node; // @[InputUnit.scala 191:19]
  reg [2:0] states_1_g; // @[InputUnit.scala 191:19]
  reg  states_1_vc_sel_2_0; // @[InputUnit.scala 191:19]
  reg  states_1_vc_sel_1_0; // @[InputUnit.scala 191:19]
  reg  states_1_vc_sel_1_1; // @[InputUnit.scala 191:19]
  reg  states_1_vc_sel_0_0; // @[InputUnit.scala 191:19]
  reg [1:0] states_1_flow_ingress_node; // @[InputUnit.scala 191:19]
  reg [1:0] states_1_flow_egress_node; // @[InputUnit.scala 191:19]
  reg [2:0] states_2_g; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_2_0; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_1_0; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_1_1; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_1_2; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_0_0; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_0_1; // @[InputUnit.scala 191:19]
  reg [1:0] states_2_flow_ingress_node; // @[InputUnit.scala 191:19]
  reg [1:0] states_2_flow_egress_node; // @[InputUnit.scala 191:19]
  reg [2:0] states_3_g; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_2_0; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_1_0; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_1_1; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_1_2; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_1_3; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_0_0; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_0_1; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_0_2; // @[InputUnit.scala 191:19]
  reg [1:0] states_3_flow_ingress_node; // @[InputUnit.scala 191:19]
  reg [1:0] states_3_flow_egress_node; // @[InputUnit.scala 191:19]
  wire  _T = io_in_flit_0_valid & io_in_flit_0_bits_head; // @[InputUnit.scala 194:32]
  wire  _T_3 = ~reset; // @[InputUnit.scala 196:13]
  wire [2:0] _GEN_1 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? states_1_g : states_0_g; // @[InputUnit.scala 197:{27,27}]
  wire [2:0] _GEN_2 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? states_2_g : _GEN_1; // @[InputUnit.scala 197:{27,27}]
  wire [2:0] _GEN_3 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? states_3_g : _GEN_2; // @[InputUnit.scala 197:{27,27}]
  wire  at_dest = io_in_flit_0_bits_flow_egress_node == 2'h3; // @[InputUnit.scala 198:57]
  wire [2:0] _states_g_T = at_dest ? 3'h2 : 3'h1; // @[InputUnit.scala 199:26]
  wire [2:0] _GEN_4 = 2'h0 == io_in_flit_0_bits_virt_channel_id ? _states_g_T : states_0_g; // @[InputUnit.scala 191:19 199:{20,20}]
  wire [2:0] _GEN_5 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? _states_g_T : states_1_g; // @[InputUnit.scala 191:19 199:{20,20}]
  wire [2:0] _GEN_6 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? _states_g_T : states_2_g; // @[InputUnit.scala 191:19 199:{20,20}]
  wire [2:0] _GEN_7 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? _states_g_T : states_3_g; // @[InputUnit.scala 191:19 199:{20,20}]
  wire  _GEN_8 = 2'h0 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_0_vc_sel_0_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_9 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_1_vc_sel_0_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_10 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_0_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_11 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_0_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_14 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_0_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_15 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_0_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_19 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_0_2; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_24 = 2'h0 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_0_vc_sel_1_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_25 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_1_vc_sel_1_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_26 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_1_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_27 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_1_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_29 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_1_vc_sel_1_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_30 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_1_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_31 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_1_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_34 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_1_2; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_35 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_1_2; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_39 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_1_3; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_40 = 2'h0 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_0_vc_sel_2_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_41 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_1_vc_sel_2_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_42 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_2_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_43 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_2_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_44 = 2'h0 == io_in_flit_0_bits_virt_channel_id | _GEN_40; // @[InputUnit.scala 203:{44,44}]
  wire  _GEN_45 = 2'h1 == io_in_flit_0_bits_virt_channel_id | _GEN_41; // @[InputUnit.scala 203:{44,44}]
  wire  _GEN_46 = 2'h2 == io_in_flit_0_bits_virt_channel_id | _GEN_42; // @[InputUnit.scala 203:{44,44}]
  wire  _GEN_47 = 2'h3 == io_in_flit_0_bits_virt_channel_id | _GEN_43; // @[InputUnit.scala 203:{44,44}]
  wire [2:0] _GEN_72 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_4 : states_0_g; // @[InputUnit.scala 191:19 194:60]
  wire [2:0] _GEN_73 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_5 : states_1_g; // @[InputUnit.scala 191:19 194:60]
  wire [2:0] _GEN_74 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_6 : states_2_g; // @[InputUnit.scala 191:19 194:60]
  wire [2:0] _GEN_75 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_7 : states_3_g; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_76 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_8 : states_0_vc_sel_0_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_77 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_9 : states_1_vc_sel_0_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_78 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_10 : states_2_vc_sel_0_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_79 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_11 : states_3_vc_sel_0_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_82 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_14 : states_2_vc_sel_0_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_83 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_15 : states_3_vc_sel_0_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_87 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_19 : states_3_vc_sel_0_2; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_92 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_24 : states_0_vc_sel_1_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_93 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_25 : states_1_vc_sel_1_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_94 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_26 : states_2_vc_sel_1_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_95 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_27 : states_3_vc_sel_1_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_97 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_29 : states_1_vc_sel_1_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_98 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_30 : states_2_vc_sel_1_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_99 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_31 : states_3_vc_sel_1_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_102 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_34 : states_2_vc_sel_1_2; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_103 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_35 : states_3_vc_sel_1_2; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_107 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_39 : states_3_vc_sel_1_3; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_108 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_44 : states_0_vc_sel_2_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_109 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_45 : states_1_vc_sel_2_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_110 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_46 : states_2_vc_sel_2_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_111 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_47 : states_3_vc_sel_2_0; // @[InputUnit.scala 191:19 194:60]
  wire  _T_10 = route_arbiter_io_in_0_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_132 = _T_10 ? 3'h2 : _GEN_72; // @[InputUnit.scala 215:{23,29}]
  wire  _T_11 = route_arbiter_io_in_1_ready & route_arbiter_io_in_1_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_133 = _T_11 ? 3'h2 : _GEN_73; // @[InputUnit.scala 215:{23,29}]
  wire  _T_12 = route_arbiter_io_in_2_ready & route_arbiter_io_in_2_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_134 = _T_12 ? 3'h2 : _GEN_74; // @[InputUnit.scala 215:{23,29}]
  wire  _T_13 = route_arbiter_io_in_3_ready & route_arbiter_io_in_3_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_135 = _T_13 ? 3'h2 : _GEN_75; // @[InputUnit.scala 215:{23,29}]
  wire [2:0] _GEN_137 = 2'h1 == io_router_req_bits_src_virt_id ? states_1_g : states_0_g; // @[InputUnit.scala 224:{25,25}]
  wire [2:0] _GEN_138 = 2'h2 == io_router_req_bits_src_virt_id ? states_2_g : _GEN_137; // @[InputUnit.scala 224:{25,25}]
  wire [2:0] _GEN_139 = 2'h3 == io_router_req_bits_src_virt_id ? states_3_g : _GEN_138; // @[InputUnit.scala 224:{25,25}]
  wire [2:0] _GEN_140 = 2'h0 == io_router_req_bits_src_virt_id ? 3'h2 : _GEN_132; // @[InputUnit.scala 225:{18,18}]
  wire [2:0] _GEN_141 = 2'h1 == io_router_req_bits_src_virt_id ? 3'h2 : _GEN_133; // @[InputUnit.scala 225:{18,18}]
  wire [2:0] _GEN_142 = 2'h2 == io_router_req_bits_src_virt_id ? 3'h2 : _GEN_134; // @[InputUnit.scala 225:{18,18}]
  wire [2:0] _GEN_143 = 2'h3 == io_router_req_bits_src_virt_id ? 3'h2 : _GEN_135; // @[InputUnit.scala 225:{18,18}]
  wire  _GEN_144 = 2'h0 == io_router_req_bits_src_virt_id ? 1'h0 : _GEN_108; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_145 = 2'h0 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_0 : _GEN_92; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_149 = 2'h0 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_0 : _GEN_76; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_153 = 2'h1 == io_router_req_bits_src_virt_id ? 1'h0 : _GEN_109; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_154 = 2'h1 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_0 : _GEN_93; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_155 = 2'h1 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_1 : _GEN_97; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_158 = 2'h1 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_0 : _GEN_77; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_162 = 2'h2 == io_router_req_bits_src_virt_id ? 1'h0 : _GEN_110; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_163 = 2'h2 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_0 : _GEN_94; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_164 = 2'h2 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_1 : _GEN_98; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_165 = 2'h2 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_2 : _GEN_102; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_167 = 2'h2 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_0 : _GEN_78; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_168 = 2'h2 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_1 : _GEN_82; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_171 = 2'h3 == io_router_req_bits_src_virt_id ? 1'h0 : _GEN_111; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_172 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_0 : _GEN_95; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_173 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_1 : _GEN_99; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_174 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_2 : _GEN_103; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_175 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_3 : _GEN_107; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_176 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_0 : _GEN_79; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_177 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_1 : _GEN_83; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_178 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_2 : _GEN_87; // @[InputUnit.scala 227:25 228:26]
  wire [2:0] _GEN_180 = io_router_req_valid ? _GEN_140 : _GEN_132; // @[InputUnit.scala 222:31]
  wire [2:0] _GEN_181 = io_router_req_valid ? _GEN_141 : _GEN_133; // @[InputUnit.scala 222:31]
  wire [2:0] _GEN_182 = io_router_req_valid ? _GEN_142 : _GEN_134; // @[InputUnit.scala 222:31]
  wire [2:0] _GEN_183 = io_router_req_valid ? _GEN_143 : _GEN_135; // @[InputUnit.scala 222:31]
  wire  _GEN_184 = io_router_req_valid ? _GEN_144 : _GEN_108; // @[InputUnit.scala 222:31]
  wire  _GEN_185 = io_router_req_valid ? _GEN_145 : _GEN_92; // @[InputUnit.scala 222:31]
  wire  _GEN_189 = io_router_req_valid ? _GEN_149 : _GEN_76; // @[InputUnit.scala 222:31]
  wire  _GEN_193 = io_router_req_valid ? _GEN_153 : _GEN_109; // @[InputUnit.scala 222:31]
  wire  _GEN_194 = io_router_req_valid ? _GEN_154 : _GEN_93; // @[InputUnit.scala 222:31]
  wire  _GEN_195 = io_router_req_valid ? _GEN_155 : _GEN_97; // @[InputUnit.scala 222:31]
  wire  _GEN_198 = io_router_req_valid ? _GEN_158 : _GEN_77; // @[InputUnit.scala 222:31]
  wire  _GEN_202 = io_router_req_valid ? _GEN_162 : _GEN_110; // @[InputUnit.scala 222:31]
  wire  _GEN_203 = io_router_req_valid ? _GEN_163 : _GEN_94; // @[InputUnit.scala 222:31]
  wire  _GEN_204 = io_router_req_valid ? _GEN_164 : _GEN_98; // @[InputUnit.scala 222:31]
  wire  _GEN_205 = io_router_req_valid ? _GEN_165 : _GEN_102; // @[InputUnit.scala 222:31]
  wire  _GEN_207 = io_router_req_valid ? _GEN_167 : _GEN_78; // @[InputUnit.scala 222:31]
  wire  _GEN_208 = io_router_req_valid ? _GEN_168 : _GEN_82; // @[InputUnit.scala 222:31]
  wire  _GEN_211 = io_router_req_valid ? _GEN_171 : _GEN_111; // @[InputUnit.scala 222:31]
  wire  _GEN_212 = io_router_req_valid ? _GEN_172 : _GEN_95; // @[InputUnit.scala 222:31]
  wire  _GEN_213 = io_router_req_valid ? _GEN_173 : _GEN_99; // @[InputUnit.scala 222:31]
  wire  _GEN_214 = io_router_req_valid ? _GEN_174 : _GEN_103; // @[InputUnit.scala 222:31]
  wire  _GEN_215 = io_router_req_valid ? _GEN_175 : _GEN_107; // @[InputUnit.scala 222:31]
  wire  _GEN_216 = io_router_req_valid ? _GEN_176 : _GEN_79; // @[InputUnit.scala 222:31]
  wire  _GEN_217 = io_router_req_valid ? _GEN_177 : _GEN_83; // @[InputUnit.scala 222:31]
  wire  _GEN_218 = io_router_req_valid ? _GEN_178 : _GEN_87; // @[InputUnit.scala 222:31]
  reg [3:0] mask; // @[InputUnit.scala 233:21]
  wire  vcalloc_vals_1 = states_1_g == 3'h2; // @[InputUnit.scala 249:32]
  wire  vcalloc_vals_0 = states_0_g == 3'h2; // @[InputUnit.scala 249:32]
  wire  vcalloc_vals_3 = states_3_g == 3'h2; // @[InputUnit.scala 249:32]
  wire  vcalloc_vals_2 = states_2_g == 3'h2; // @[InputUnit.scala 249:32]
  wire [3:0] _vcalloc_filter_T = {vcalloc_vals_3,vcalloc_vals_2,vcalloc_vals_1,vcalloc_vals_0}; // @[InputUnit.scala 236:59]
  wire [3:0] _vcalloc_filter_T_2 = ~mask; // @[InputUnit.scala 236:89]
  wire [3:0] _vcalloc_filter_T_3 = _vcalloc_filter_T & _vcalloc_filter_T_2; // @[InputUnit.scala 236:87]
  wire [7:0] _vcalloc_filter_T_4 = {vcalloc_vals_3,vcalloc_vals_2,vcalloc_vals_1,vcalloc_vals_0,_vcalloc_filter_T_3}; // @[Cat.scala 33:92]
  wire [7:0] _vcalloc_filter_T_13 = _vcalloc_filter_T_4[7] ? 8'h80 : 8'h0; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_14 = _vcalloc_filter_T_4[6] ? 8'h40 : _vcalloc_filter_T_13; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_15 = _vcalloc_filter_T_4[5] ? 8'h20 : _vcalloc_filter_T_14; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_16 = _vcalloc_filter_T_4[4] ? 8'h10 : _vcalloc_filter_T_15; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_17 = _vcalloc_filter_T_4[3] ? 8'h8 : _vcalloc_filter_T_16; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_18 = _vcalloc_filter_T_4[2] ? 8'h4 : _vcalloc_filter_T_17; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_19 = _vcalloc_filter_T_4[1] ? 8'h2 : _vcalloc_filter_T_18; // @[Mux.scala 47:70]
  wire [7:0] vcalloc_filter = _vcalloc_filter_T_4[0] ? 8'h1 : _vcalloc_filter_T_19; // @[Mux.scala 47:70]
  wire [3:0] vcalloc_sel = vcalloc_filter[3:0] | vcalloc_filter[7:4]; // @[InputUnit.scala 237:58]
  wire [3:0] _mask_T = 4'h1 << io_router_req_bits_src_virt_id; // @[InputUnit.scala 240:18]
  wire [3:0] _mask_T_2 = _mask_T - 4'h1; // @[InputUnit.scala 240:53]
  wire  _T_26 = vcalloc_vals_0 | vcalloc_vals_1 | vcalloc_vals_2 | vcalloc_vals_3; // @[package.scala 73:59]
  wire [1:0] _mask_T_12 = vcalloc_sel[1] ? 2'h3 : 2'h0; // @[Mux.scala 27:73]
  wire [2:0] _mask_T_13 = vcalloc_sel[2] ? 3'h7 : 3'h0; // @[Mux.scala 27:73]
  wire [3:0] _mask_T_14 = vcalloc_sel[3] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [1:0] _GEN_60 = {{1'd0}, vcalloc_sel[0]}; // @[Mux.scala 27:73]
  wire [1:0] _mask_T_15 = _GEN_60 | _mask_T_12; // @[Mux.scala 27:73]
  wire [2:0] _GEN_61 = {{1'd0}, _mask_T_15}; // @[Mux.scala 27:73]
  wire [2:0] _mask_T_16 = _GEN_61 | _mask_T_13; // @[Mux.scala 27:73]
  wire [3:0] _GEN_62 = {{1'd0}, _mask_T_16}; // @[Mux.scala 27:73]
  wire [3:0] _mask_T_17 = _GEN_62 | _mask_T_14; // @[Mux.scala 27:73]
  wire [2:0] _GEN_222 = vcalloc_vals_0 & vcalloc_sel[0] & io_vcalloc_req_ready ? 3'h3 : _GEN_180; // @[InputUnit.scala 253:{76,82}]
  wire [2:0] _GEN_223 = vcalloc_vals_1 & vcalloc_sel[1] & io_vcalloc_req_ready ? 3'h3 : _GEN_181; // @[InputUnit.scala 253:{76,82}]
  wire [2:0] _GEN_224 = vcalloc_vals_2 & vcalloc_sel[2] & io_vcalloc_req_ready ? 3'h3 : _GEN_182; // @[InputUnit.scala 253:{76,82}]
  wire [2:0] _GEN_225 = vcalloc_vals_3 & vcalloc_sel[3] & io_vcalloc_req_ready ? 3'h3 : _GEN_183; // @[InputUnit.scala 253:{76,82}]
  wire [1:0] _io_debug_va_stall_T = vcalloc_vals_0 + vcalloc_vals_1; // @[Bitwise.scala 51:90]
  wire [1:0] _io_debug_va_stall_T_2 = vcalloc_vals_2 + vcalloc_vals_3; // @[Bitwise.scala 51:90]
  wire [2:0] _io_debug_va_stall_T_4 = _io_debug_va_stall_T + _io_debug_va_stall_T_2; // @[Bitwise.scala 51:90]
  wire [2:0] _GEN_63 = {{2'd0}, io_vcalloc_req_ready}; // @[InputUnit.scala 266:47]
  wire [2:0] _io_debug_va_stall_T_7 = _io_debug_va_stall_T_4 - _GEN_63; // @[InputUnit.scala 266:47]
  wire  _T_39 = io_vcalloc_req_ready & io_vcalloc_req_valid; // @[Decoupled.scala 51:35]
  wire [8:0] _credit_available_T = {states_0_vc_sel_2_0,1'h0,1'h0,1'h0,states_0_vc_sel_1_0,2'h0,1'h0,states_0_vc_sel_0_0
    }; // @[InputUnit.scala 287:40]
  wire [8:0] _credit_available_T_1 = {io_out_credit_available_2_0,io_out_credit_available_1_3,
    io_out_credit_available_1_2,io_out_credit_available_1_1,io_out_credit_available_1_0,io_out_credit_available_0_3,
    io_out_credit_available_0_2,io_out_credit_available_0_1,io_out_credit_available_0_0}; // @[InputUnit.scala 287:73]
  wire [8:0] _credit_available_T_2 = _credit_available_T & _credit_available_T_1; // @[InputUnit.scala 287:47]
  wire  credit_available = _credit_available_T_2 != 9'h0; // @[InputUnit.scala 287:81]
  wire  _T_60 = salloc_arb_io_in_0_ready & salloc_arb_io_in_0_valid; // @[Decoupled.scala 51:35]
  wire [8:0] _credit_available_T_3 = {states_1_vc_sel_2_0,1'h0,1'h0,states_1_vc_sel_1_1,states_1_vc_sel_1_0,2'h0,1'h0,
    states_1_vc_sel_0_0}; // @[InputUnit.scala 287:40]
  wire [8:0] _credit_available_T_5 = _credit_available_T_3 & _credit_available_T_1; // @[InputUnit.scala 287:47]
  wire  credit_available_1 = _credit_available_T_5 != 9'h0; // @[InputUnit.scala 287:81]
  wire  _T_62 = salloc_arb_io_in_1_ready & salloc_arb_io_in_1_valid; // @[Decoupled.scala 51:35]
  wire [8:0] _credit_available_T_6 = {states_2_vc_sel_2_0,1'h0,states_2_vc_sel_1_2,states_2_vc_sel_1_1,
    states_2_vc_sel_1_0,2'h0,states_2_vc_sel_0_1,states_2_vc_sel_0_0}; // @[InputUnit.scala 287:40]
  wire [8:0] _credit_available_T_8 = _credit_available_T_6 & _credit_available_T_1; // @[InputUnit.scala 287:47]
  wire  credit_available_2 = _credit_available_T_8 != 9'h0; // @[InputUnit.scala 287:81]
  wire  _T_64 = salloc_arb_io_in_2_ready & salloc_arb_io_in_2_valid; // @[Decoupled.scala 51:35]
  wire [8:0] _credit_available_T_9 = {states_3_vc_sel_2_0,states_3_vc_sel_1_3,states_3_vc_sel_1_2,states_3_vc_sel_1_1,
    states_3_vc_sel_1_0,1'h0,states_3_vc_sel_0_2,states_3_vc_sel_0_1,states_3_vc_sel_0_0}; // @[InputUnit.scala 287:40]
  wire [8:0] _credit_available_T_11 = _credit_available_T_9 & _credit_available_T_1; // @[InputUnit.scala 287:47]
  wire  credit_available_3 = _credit_available_T_11 != 9'h0; // @[InputUnit.scala 287:81]
  wire  _T_66 = salloc_arb_io_in_3_ready & salloc_arb_io_in_3_valid; // @[Decoupled.scala 51:35]
  wire  _io_debug_sa_stall_T_1 = salloc_arb_io_in_0_valid & ~salloc_arb_io_in_0_ready; // @[InputUnit.scala 301:67]
  wire  _io_debug_sa_stall_T_3 = salloc_arb_io_in_1_valid & ~salloc_arb_io_in_1_ready; // @[InputUnit.scala 301:67]
  wire  _io_debug_sa_stall_T_5 = salloc_arb_io_in_2_valid & ~salloc_arb_io_in_2_ready; // @[InputUnit.scala 301:67]
  wire  _io_debug_sa_stall_T_7 = salloc_arb_io_in_3_valid & ~salloc_arb_io_in_3_ready; // @[InputUnit.scala 301:67]
  wire [1:0] _io_debug_sa_stall_T_8 = _io_debug_sa_stall_T_1 + _io_debug_sa_stall_T_3; // @[Bitwise.scala 51:90]
  wire [1:0] _io_debug_sa_stall_T_10 = _io_debug_sa_stall_T_5 + _io_debug_sa_stall_T_7; // @[Bitwise.scala 51:90]
  wire [2:0] _io_debug_sa_stall_T_12 = _io_debug_sa_stall_T_8 + _io_debug_sa_stall_T_10; // @[Bitwise.scala 51:90]
  reg  salloc_outs_0_valid; // @[InputUnit.scala 318:8]
  reg [1:0] salloc_outs_0_out_vid; // @[InputUnit.scala 318:8]
  reg  salloc_outs_0_flit_head; // @[InputUnit.scala 318:8]
  reg  salloc_outs_0_flit_tail; // @[InputUnit.scala 318:8]
  reg [63:0] salloc_outs_0_flit_payload; // @[InputUnit.scala 318:8]
  reg [1:0] salloc_outs_0_flit_flow_ingress_node; // @[InputUnit.scala 318:8]
  reg [1:0] salloc_outs_0_flit_flow_egress_node; // @[InputUnit.scala 318:8]
  wire  _io_in_credit_return_T = salloc_arb_io_out_0_ready & salloc_arb_io_out_0_valid; // @[Decoupled.scala 51:35]
  wire  _io_in_vc_free_T_11 = salloc_arb_io_chosen_oh_0[0] & input_buffer_io_deq_0_bits_tail | salloc_arb_io_chosen_oh_0
    [1] & input_buffer_io_deq_1_bits_tail | salloc_arb_io_chosen_oh_0[2] & input_buffer_io_deq_2_bits_tail |
    salloc_arb_io_chosen_oh_0[3] & input_buffer_io_deq_3_bits_tail; // @[Mux.scala 27:73]
  wire  vc_sel_0_0 = salloc_arb_io_chosen_oh_0[0] & states_0_vc_sel_0_0 | salloc_arb_io_chosen_oh_0[1] &
    states_1_vc_sel_0_0 | salloc_arb_io_chosen_oh_0[2] & states_2_vc_sel_0_0 | salloc_arb_io_chosen_oh_0[3] &
    states_3_vc_sel_0_0; // @[Mux.scala 27:73]
  wire  vc_sel_0_1 = salloc_arb_io_chosen_oh_0[2] & states_2_vc_sel_0_1 | salloc_arb_io_chosen_oh_0[3] &
    states_3_vc_sel_0_1; // @[Mux.scala 27:73]
  wire  vc_sel_0_2 = salloc_arb_io_chosen_oh_0[3] & states_3_vc_sel_0_2; // @[Mux.scala 27:73]
  wire  vc_sel_1_0 = salloc_arb_io_chosen_oh_0[0] & states_0_vc_sel_1_0 | salloc_arb_io_chosen_oh_0[1] &
    states_1_vc_sel_1_0 | salloc_arb_io_chosen_oh_0[2] & states_2_vc_sel_1_0 | salloc_arb_io_chosen_oh_0[3] &
    states_3_vc_sel_1_0; // @[Mux.scala 27:73]
  wire  vc_sel_1_1 = salloc_arb_io_chosen_oh_0[1] & states_1_vc_sel_1_1 | salloc_arb_io_chosen_oh_0[2] &
    states_2_vc_sel_1_1 | salloc_arb_io_chosen_oh_0[3] & states_3_vc_sel_1_1; // @[Mux.scala 27:73]
  wire  vc_sel_1_2 = salloc_arb_io_chosen_oh_0[2] & states_2_vc_sel_1_2 | salloc_arb_io_chosen_oh_0[3] &
    states_3_vc_sel_1_2; // @[Mux.scala 27:73]
  wire  vc_sel_1_3 = salloc_arb_io_chosen_oh_0[3] & states_3_vc_sel_1_3; // @[Mux.scala 27:73]
  wire  channel_oh_0 = vc_sel_0_0 | vc_sel_0_1 | vc_sel_0_2; // @[InputUnit.scala 334:43]
  wire  channel_oh_1 = vc_sel_1_0 | vc_sel_1_1 | vc_sel_1_2 | vc_sel_1_3; // @[InputUnit.scala 334:43]
  wire [3:0] _virt_channel_T = {1'h0,vc_sel_0_2,vc_sel_0_1,vc_sel_0_0}; // @[OneHot.scala 22:45]
  wire [1:0] virt_channel_hi_1 = _virt_channel_T[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] virt_channel_lo_1 = _virt_channel_T[1:0]; // @[OneHot.scala 31:18]
  wire  _virt_channel_T_1 = |virt_channel_hi_1; // @[OneHot.scala 32:14]
  wire [1:0] _virt_channel_T_2 = virt_channel_hi_1 | virt_channel_lo_1; // @[OneHot.scala 32:28]
  wire [1:0] _virt_channel_T_4 = {_virt_channel_T_1,_virt_channel_T_2[1]}; // @[Cat.scala 33:92]
  wire [3:0] _virt_channel_T_5 = {vc_sel_1_3,vc_sel_1_2,vc_sel_1_1,vc_sel_1_0}; // @[OneHot.scala 22:45]
  wire [1:0] virt_channel_hi_3 = _virt_channel_T_5[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] virt_channel_lo_3 = _virt_channel_T_5[1:0]; // @[OneHot.scala 31:18]
  wire  _virt_channel_T_6 = |virt_channel_hi_3; // @[OneHot.scala 32:14]
  wire [1:0] _virt_channel_T_7 = virt_channel_hi_3 | virt_channel_lo_3; // @[OneHot.scala 32:28]
  wire [1:0] _virt_channel_T_9 = {_virt_channel_T_6,_virt_channel_T_7[1]}; // @[Cat.scala 33:92]
  wire [1:0] _virt_channel_T_10 = channel_oh_0 ? _virt_channel_T_4 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _virt_channel_T_11 = channel_oh_1 ? _virt_channel_T_9 : 2'h0; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_4 = salloc_arb_io_chosen_oh_0[0] ? input_buffer_io_deq_0_bits_payload : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_5 = salloc_arb_io_chosen_oh_0[1] ? input_buffer_io_deq_1_bits_payload : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_6 = salloc_arb_io_chosen_oh_0[2] ? input_buffer_io_deq_2_bits_payload : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_7 = salloc_arb_io_chosen_oh_0[3] ? input_buffer_io_deq_3_bits_payload : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_8 = _salloc_outs_0_flit_payload_T_4 | _salloc_outs_0_flit_payload_T_5; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_9 = _salloc_outs_0_flit_payload_T_8 | _salloc_outs_0_flit_payload_T_6; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_11 = salloc_arb_io_chosen_oh_0[0] ? states_0_flow_egress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_12 = salloc_arb_io_chosen_oh_0[1] ? states_1_flow_egress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_13 = salloc_arb_io_chosen_oh_0[2] ? states_2_flow_egress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_14 = salloc_arb_io_chosen_oh_0[3] ? states_3_flow_egress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_15 = _salloc_outs_0_flit_flow_T_11 | _salloc_outs_0_flit_flow_T_12; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_16 = _salloc_outs_0_flit_flow_T_15 | _salloc_outs_0_flit_flow_T_13; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_25 = salloc_arb_io_chosen_oh_0[0] ? states_0_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_26 = salloc_arb_io_chosen_oh_0[1] ? states_1_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_27 = salloc_arb_io_chosen_oh_0[2] ? states_2_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_28 = salloc_arb_io_chosen_oh_0[3] ? states_3_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_29 = _salloc_outs_0_flit_flow_T_25 | _salloc_outs_0_flit_flow_T_26; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_30 = _salloc_outs_0_flit_flow_T_29 | _salloc_outs_0_flit_flow_T_27; // @[Mux.scala 27:73]
  InputBuffer input_buffer ( // @[InputUnit.scala 180:28]
    .clock(input_buffer_clock),
    .reset(input_buffer_reset),
    .io_enq_0_valid(input_buffer_io_enq_0_valid),
    .io_enq_0_bits_head(input_buffer_io_enq_0_bits_head),
    .io_enq_0_bits_tail(input_buffer_io_enq_0_bits_tail),
    .io_enq_0_bits_payload(input_buffer_io_enq_0_bits_payload),
    .io_enq_0_bits_virt_channel_id(input_buffer_io_enq_0_bits_virt_channel_id),
    .io_deq_0_ready(input_buffer_io_deq_0_ready),
    .io_deq_0_valid(input_buffer_io_deq_0_valid),
    .io_deq_0_bits_head(input_buffer_io_deq_0_bits_head),
    .io_deq_0_bits_tail(input_buffer_io_deq_0_bits_tail),
    .io_deq_0_bits_payload(input_buffer_io_deq_0_bits_payload),
    .io_deq_1_ready(input_buffer_io_deq_1_ready),
    .io_deq_1_valid(input_buffer_io_deq_1_valid),
    .io_deq_1_bits_head(input_buffer_io_deq_1_bits_head),
    .io_deq_1_bits_tail(input_buffer_io_deq_1_bits_tail),
    .io_deq_1_bits_payload(input_buffer_io_deq_1_bits_payload),
    .io_deq_2_ready(input_buffer_io_deq_2_ready),
    .io_deq_2_valid(input_buffer_io_deq_2_valid),
    .io_deq_2_bits_head(input_buffer_io_deq_2_bits_head),
    .io_deq_2_bits_tail(input_buffer_io_deq_2_bits_tail),
    .io_deq_2_bits_payload(input_buffer_io_deq_2_bits_payload),
    .io_deq_3_ready(input_buffer_io_deq_3_ready),
    .io_deq_3_valid(input_buffer_io_deq_3_valid),
    .io_deq_3_bits_head(input_buffer_io_deq_3_bits_head),
    .io_deq_3_bits_tail(input_buffer_io_deq_3_bits_tail),
    .io_deq_3_bits_payload(input_buffer_io_deq_3_bits_payload)
  );
  Arbiter route_arbiter ( // @[InputUnit.scala 186:29]
    .io_in_0_valid(route_arbiter_io_in_0_valid),
    .io_in_0_bits_flow_ingress_node(route_arbiter_io_in_0_bits_flow_ingress_node),
    .io_in_0_bits_flow_egress_node(route_arbiter_io_in_0_bits_flow_egress_node),
    .io_in_1_ready(route_arbiter_io_in_1_ready),
    .io_in_1_valid(route_arbiter_io_in_1_valid),
    .io_in_1_bits_flow_ingress_node(route_arbiter_io_in_1_bits_flow_ingress_node),
    .io_in_1_bits_flow_egress_node(route_arbiter_io_in_1_bits_flow_egress_node),
    .io_in_2_ready(route_arbiter_io_in_2_ready),
    .io_in_2_valid(route_arbiter_io_in_2_valid),
    .io_in_2_bits_flow_ingress_node(route_arbiter_io_in_2_bits_flow_ingress_node),
    .io_in_2_bits_flow_egress_node(route_arbiter_io_in_2_bits_flow_egress_node),
    .io_in_3_ready(route_arbiter_io_in_3_ready),
    .io_in_3_valid(route_arbiter_io_in_3_valid),
    .io_in_3_bits_flow_ingress_node(route_arbiter_io_in_3_bits_flow_ingress_node),
    .io_in_3_bits_flow_egress_node(route_arbiter_io_in_3_bits_flow_egress_node),
    .io_out_valid(route_arbiter_io_out_valid),
    .io_out_bits_src_virt_id(route_arbiter_io_out_bits_src_virt_id),
    .io_out_bits_flow_ingress_node(route_arbiter_io_out_bits_flow_ingress_node),
    .io_out_bits_flow_egress_node(route_arbiter_io_out_bits_flow_egress_node)
  );
  SwitchArbiter salloc_arb ( // @[InputUnit.scala 279:26]
    .clock(salloc_arb_clock),
    .reset(salloc_arb_reset),
    .io_in_0_ready(salloc_arb_io_in_0_ready),
    .io_in_0_valid(salloc_arb_io_in_0_valid),
    .io_in_0_bits_vc_sel_2_0(salloc_arb_io_in_0_bits_vc_sel_2_0),
    .io_in_0_bits_vc_sel_1_0(salloc_arb_io_in_0_bits_vc_sel_1_0),
    .io_in_0_bits_vc_sel_0_0(salloc_arb_io_in_0_bits_vc_sel_0_0),
    .io_in_0_bits_tail(salloc_arb_io_in_0_bits_tail),
    .io_in_1_ready(salloc_arb_io_in_1_ready),
    .io_in_1_valid(salloc_arb_io_in_1_valid),
    .io_in_1_bits_vc_sel_2_0(salloc_arb_io_in_1_bits_vc_sel_2_0),
    .io_in_1_bits_vc_sel_1_0(salloc_arb_io_in_1_bits_vc_sel_1_0),
    .io_in_1_bits_vc_sel_1_1(salloc_arb_io_in_1_bits_vc_sel_1_1),
    .io_in_1_bits_vc_sel_0_0(salloc_arb_io_in_1_bits_vc_sel_0_0),
    .io_in_1_bits_vc_sel_0_1(salloc_arb_io_in_1_bits_vc_sel_0_1),
    .io_in_1_bits_tail(salloc_arb_io_in_1_bits_tail),
    .io_in_2_ready(salloc_arb_io_in_2_ready),
    .io_in_2_valid(salloc_arb_io_in_2_valid),
    .io_in_2_bits_vc_sel_2_0(salloc_arb_io_in_2_bits_vc_sel_2_0),
    .io_in_2_bits_vc_sel_1_0(salloc_arb_io_in_2_bits_vc_sel_1_0),
    .io_in_2_bits_vc_sel_1_1(salloc_arb_io_in_2_bits_vc_sel_1_1),
    .io_in_2_bits_vc_sel_1_2(salloc_arb_io_in_2_bits_vc_sel_1_2),
    .io_in_2_bits_vc_sel_0_0(salloc_arb_io_in_2_bits_vc_sel_0_0),
    .io_in_2_bits_vc_sel_0_1(salloc_arb_io_in_2_bits_vc_sel_0_1),
    .io_in_2_bits_vc_sel_0_2(salloc_arb_io_in_2_bits_vc_sel_0_2),
    .io_in_2_bits_tail(salloc_arb_io_in_2_bits_tail),
    .io_in_3_ready(salloc_arb_io_in_3_ready),
    .io_in_3_valid(salloc_arb_io_in_3_valid),
    .io_in_3_bits_vc_sel_2_0(salloc_arb_io_in_3_bits_vc_sel_2_0),
    .io_in_3_bits_vc_sel_1_0(salloc_arb_io_in_3_bits_vc_sel_1_0),
    .io_in_3_bits_vc_sel_1_1(salloc_arb_io_in_3_bits_vc_sel_1_1),
    .io_in_3_bits_vc_sel_1_2(salloc_arb_io_in_3_bits_vc_sel_1_2),
    .io_in_3_bits_vc_sel_1_3(salloc_arb_io_in_3_bits_vc_sel_1_3),
    .io_in_3_bits_vc_sel_0_0(salloc_arb_io_in_3_bits_vc_sel_0_0),
    .io_in_3_bits_vc_sel_0_1(salloc_arb_io_in_3_bits_vc_sel_0_1),
    .io_in_3_bits_vc_sel_0_2(salloc_arb_io_in_3_bits_vc_sel_0_2),
    .io_in_3_bits_vc_sel_0_3(salloc_arb_io_in_3_bits_vc_sel_0_3),
    .io_in_3_bits_tail(salloc_arb_io_in_3_bits_tail),
    .io_out_0_ready(salloc_arb_io_out_0_ready),
    .io_out_0_valid(salloc_arb_io_out_0_valid),
    .io_out_0_bits_vc_sel_2_0(salloc_arb_io_out_0_bits_vc_sel_2_0),
    .io_out_0_bits_vc_sel_1_0(salloc_arb_io_out_0_bits_vc_sel_1_0),
    .io_out_0_bits_vc_sel_1_1(salloc_arb_io_out_0_bits_vc_sel_1_1),
    .io_out_0_bits_vc_sel_1_2(salloc_arb_io_out_0_bits_vc_sel_1_2),
    .io_out_0_bits_vc_sel_1_3(salloc_arb_io_out_0_bits_vc_sel_1_3),
    .io_out_0_bits_vc_sel_0_0(salloc_arb_io_out_0_bits_vc_sel_0_0),
    .io_out_0_bits_vc_sel_0_1(salloc_arb_io_out_0_bits_vc_sel_0_1),
    .io_out_0_bits_vc_sel_0_2(salloc_arb_io_out_0_bits_vc_sel_0_2),
    .io_out_0_bits_vc_sel_0_3(salloc_arb_io_out_0_bits_vc_sel_0_3),
    .io_out_0_bits_tail(salloc_arb_io_out_0_bits_tail),
    .io_chosen_oh_0(salloc_arb_io_chosen_oh_0)
  );
  assign io_router_req_valid = route_arbiter_io_out_valid; // @[InputUnit.scala 189:17]
  assign io_router_req_bits_src_virt_id = route_arbiter_io_out_bits_src_virt_id; // @[InputUnit.scala 189:17]
  assign io_router_req_bits_flow_ingress_node = route_arbiter_io_out_bits_flow_ingress_node; // @[InputUnit.scala 189:17]
  assign io_router_req_bits_flow_egress_node = route_arbiter_io_out_bits_flow_egress_node; // @[InputUnit.scala 189:17]
  assign io_vcalloc_req_valid = vcalloc_vals_0 | vcalloc_vals_1 | vcalloc_vals_2 | vcalloc_vals_3; // @[package.scala 73:59]
  assign io_vcalloc_req_bits_vc_sel_2_0 = vcalloc_sel[0] & states_0_vc_sel_2_0 | vcalloc_sel[1] & states_1_vc_sel_2_0 |
    vcalloc_sel[2] & states_2_vc_sel_2_0 | vcalloc_sel[3] & states_3_vc_sel_2_0; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_1_0 = vcalloc_sel[0] & states_0_vc_sel_1_0 | vcalloc_sel[1] & states_1_vc_sel_1_0 |
    vcalloc_sel[2] & states_2_vc_sel_1_0 | vcalloc_sel[3] & states_3_vc_sel_1_0; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_1_1 = vcalloc_sel[1] & states_1_vc_sel_1_1 | vcalloc_sel[2] & states_2_vc_sel_1_1 |
    vcalloc_sel[3] & states_3_vc_sel_1_1; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_1_2 = vcalloc_sel[2] & states_2_vc_sel_1_2 | vcalloc_sel[3] & states_3_vc_sel_1_2; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_1_3 = vcalloc_sel[3] & states_3_vc_sel_1_3; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_0_0 = vcalloc_sel[0] & states_0_vc_sel_0_0 | vcalloc_sel[1] & states_1_vc_sel_0_0 |
    vcalloc_sel[2] & states_2_vc_sel_0_0 | vcalloc_sel[3] & states_3_vc_sel_0_0; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_0_1 = vcalloc_sel[2] & states_2_vc_sel_0_1 | vcalloc_sel[3] & states_3_vc_sel_0_1; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_0_2 = vcalloc_sel[3] & states_3_vc_sel_0_2; // @[Mux.scala 27:73]
  assign io_salloc_req_0_valid = salloc_arb_io_out_0_valid; // @[InputUnit.scala 302:17 303:19 305:35]
  assign io_salloc_req_0_bits_vc_sel_2_0 = salloc_arb_io_out_0_bits_vc_sel_2_0; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_1_0 = salloc_arb_io_out_0_bits_vc_sel_1_0; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_1_1 = salloc_arb_io_out_0_bits_vc_sel_1_1; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_1_2 = salloc_arb_io_out_0_bits_vc_sel_1_2; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_1_3 = salloc_arb_io_out_0_bits_vc_sel_1_3; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_0_0 = salloc_arb_io_out_0_bits_vc_sel_0_0; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_0_1 = salloc_arb_io_out_0_bits_vc_sel_0_1; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_0_2 = salloc_arb_io_out_0_bits_vc_sel_0_2; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_0_3 = salloc_arb_io_out_0_bits_vc_sel_0_3; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_tail = salloc_arb_io_out_0_bits_tail; // @[InputUnit.scala 302:17]
  assign io_out_0_valid = salloc_outs_0_valid; // @[InputUnit.scala 349:21]
  assign io_out_0_bits_flit_head = salloc_outs_0_flit_head; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_flit_tail = salloc_outs_0_flit_tail; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_flit_payload = salloc_outs_0_flit_payload; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_flit_flow_ingress_node = salloc_outs_0_flit_flow_ingress_node; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_flit_flow_egress_node = salloc_outs_0_flit_flow_egress_node; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_out_virt_channel = salloc_outs_0_out_vid; // @[InputUnit.scala 351:37]
  assign io_debug_va_stall = _io_debug_va_stall_T_7[1:0]; // @[InputUnit.scala 266:21]
  assign io_debug_sa_stall = _io_debug_sa_stall_T_12[1:0]; // @[InputUnit.scala 301:21]
  assign io_in_credit_return = _io_in_credit_return_T ? salloc_arb_io_chosen_oh_0 : 4'h0; // @[InputUnit.scala 322:8]
  assign io_in_vc_free = _io_in_credit_return_T & _io_in_vc_free_T_11 ? salloc_arb_io_chosen_oh_0 : 4'h0; // @[InputUnit.scala 325:8]
  assign input_buffer_clock = clock;
  assign input_buffer_reset = reset;
  assign input_buffer_io_enq_0_valid = io_in_flit_0_valid; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_head = io_in_flit_0_bits_head; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_tail = io_in_flit_0_bits_tail; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_payload = io_in_flit_0_bits_payload; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_virt_channel_id = io_in_flit_0_bits_virt_channel_id; // @[InputUnit.scala 182:28]
  assign input_buffer_io_deq_0_ready = salloc_arb_io_in_0_ready; // @[InputUnit.scala 295:36]
  assign input_buffer_io_deq_1_ready = salloc_arb_io_in_1_ready; // @[InputUnit.scala 295:36]
  assign input_buffer_io_deq_2_ready = salloc_arb_io_in_2_ready; // @[InputUnit.scala 295:36]
  assign input_buffer_io_deq_3_ready = salloc_arb_io_in_3_ready; // @[InputUnit.scala 295:36]
  assign route_arbiter_io_in_0_valid = states_0_g == 3'h1; // @[InputUnit.scala 212:22]
  assign route_arbiter_io_in_0_bits_flow_ingress_node = states_0_flow_ingress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_0_bits_flow_egress_node = states_0_flow_egress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_1_valid = states_1_g == 3'h1; // @[InputUnit.scala 212:22]
  assign route_arbiter_io_in_1_bits_flow_ingress_node = states_1_flow_ingress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_1_bits_flow_egress_node = states_1_flow_egress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_2_valid = states_2_g == 3'h1; // @[InputUnit.scala 212:22]
  assign route_arbiter_io_in_2_bits_flow_ingress_node = states_2_flow_ingress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_2_bits_flow_egress_node = states_2_flow_egress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_3_valid = states_3_g == 3'h1; // @[InputUnit.scala 212:22]
  assign route_arbiter_io_in_3_bits_flow_ingress_node = states_3_flow_ingress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_3_bits_flow_egress_node = states_3_flow_egress_node; // @[InputUnit.scala 213:19]
  assign salloc_arb_clock = clock;
  assign salloc_arb_reset = reset;
  assign salloc_arb_io_in_0_valid = states_0_g == 3'h3 & credit_available & input_buffer_io_deq_0_valid; // @[InputUnit.scala 288:50]
  assign salloc_arb_io_in_0_bits_vc_sel_2_0 = states_0_vc_sel_2_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_0_bits_vc_sel_1_0 = states_0_vc_sel_1_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_0_bits_vc_sel_0_0 = states_0_vc_sel_0_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_0_bits_tail = input_buffer_io_deq_0_bits_tail; // @[InputUnit.scala 291:19]
  assign salloc_arb_io_in_1_valid = states_1_g == 3'h3 & credit_available_1 & input_buffer_io_deq_1_valid; // @[InputUnit.scala 288:50]
  assign salloc_arb_io_in_1_bits_vc_sel_2_0 = states_1_vc_sel_2_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_1_bits_vc_sel_1_0 = states_1_vc_sel_1_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_1_bits_vc_sel_1_1 = states_1_vc_sel_1_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_1_bits_vc_sel_0_0 = states_1_vc_sel_0_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_1_bits_vc_sel_0_1 = 1'h0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_1_bits_tail = input_buffer_io_deq_1_bits_tail; // @[InputUnit.scala 291:19]
  assign salloc_arb_io_in_2_valid = states_2_g == 3'h3 & credit_available_2 & input_buffer_io_deq_2_valid; // @[InputUnit.scala 288:50]
  assign salloc_arb_io_in_2_bits_vc_sel_2_0 = states_2_vc_sel_2_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_1_0 = states_2_vc_sel_1_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_1_1 = states_2_vc_sel_1_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_1_2 = states_2_vc_sel_1_2; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_0_0 = states_2_vc_sel_0_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_0_1 = states_2_vc_sel_0_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_0_2 = 1'h0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_tail = input_buffer_io_deq_2_bits_tail; // @[InputUnit.scala 291:19]
  assign salloc_arb_io_in_3_valid = states_3_g == 3'h3 & credit_available_3 & input_buffer_io_deq_3_valid; // @[InputUnit.scala 288:50]
  assign salloc_arb_io_in_3_bits_vc_sel_2_0 = states_3_vc_sel_2_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_1_0 = states_3_vc_sel_1_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_1_1 = states_3_vc_sel_1_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_1_2 = states_3_vc_sel_1_2; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_1_3 = states_3_vc_sel_1_3; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_0_0 = states_3_vc_sel_0_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_0_1 = states_3_vc_sel_0_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_0_2 = states_3_vc_sel_0_2; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_0_3 = 1'h0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_tail = input_buffer_io_deq_3_bits_tail; // @[InputUnit.scala 291:19]
  assign salloc_arb_io_out_0_ready = io_salloc_req_0_ready; // @[InputUnit.scala 302:17 303:19 304:39]
  always @(posedge clock) begin
    if (reset) begin // @[InputUnit.scala 377:23]
      states_0_g <= 3'h0; // @[InputUnit.scala 378:24]
    end else if (_T_60 & input_buffer_io_deq_0_bits_tail) begin // @[InputUnit.scala 292:35]
      states_0_g <= 3'h0; // @[InputUnit.scala 293:13]
    end else if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[0]) begin // @[InputUnit.scala 270:29]
        states_0_g <= 3'h3; // @[InputUnit.scala 272:21]
      end else begin
        states_0_g <= _GEN_222;
      end
    end else begin
      states_0_g <= _GEN_222;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[0]) begin // @[InputUnit.scala 270:29]
        states_0_vc_sel_2_0 <= io_vcalloc_resp_vc_sel_2_0; // @[InputUnit.scala 271:26]
      end else begin
        states_0_vc_sel_2_0 <= _GEN_184;
      end
    end else begin
      states_0_vc_sel_2_0 <= _GEN_184;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[0]) begin // @[InputUnit.scala 270:29]
        states_0_vc_sel_1_0 <= io_vcalloc_resp_vc_sel_1_0; // @[InputUnit.scala 271:26]
      end else begin
        states_0_vc_sel_1_0 <= _GEN_185;
      end
    end else begin
      states_0_vc_sel_1_0 <= _GEN_185;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[0]) begin // @[InputUnit.scala 270:29]
        states_0_vc_sel_0_0 <= io_vcalloc_resp_vc_sel_0_0; // @[InputUnit.scala 271:26]
      end else begin
        states_0_vc_sel_0_0 <= _GEN_189;
      end
    end else begin
      states_0_vc_sel_0_0 <= _GEN_189;
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h0 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_0_flow_ingress_node <= io_in_flit_0_bits_flow_ingress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h0 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_0_flow_egress_node <= io_in_flit_0_bits_flow_egress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (reset) begin // @[InputUnit.scala 377:23]
      states_1_g <= 3'h0; // @[InputUnit.scala 378:24]
    end else if (_T_62 & input_buffer_io_deq_1_bits_tail) begin // @[InputUnit.scala 292:35]
      states_1_g <= 3'h0; // @[InputUnit.scala 293:13]
    end else if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_g <= 3'h3; // @[InputUnit.scala 272:21]
      end else begin
        states_1_g <= _GEN_223;
      end
    end else begin
      states_1_g <= _GEN_223;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_vc_sel_2_0 <= io_vcalloc_resp_vc_sel_2_0; // @[InputUnit.scala 271:26]
      end else begin
        states_1_vc_sel_2_0 <= _GEN_193;
      end
    end else begin
      states_1_vc_sel_2_0 <= _GEN_193;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_vc_sel_1_0 <= io_vcalloc_resp_vc_sel_1_0; // @[InputUnit.scala 271:26]
      end else begin
        states_1_vc_sel_1_0 <= _GEN_194;
      end
    end else begin
      states_1_vc_sel_1_0 <= _GEN_194;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_vc_sel_1_1 <= io_vcalloc_resp_vc_sel_1_1; // @[InputUnit.scala 271:26]
      end else begin
        states_1_vc_sel_1_1 <= _GEN_195;
      end
    end else begin
      states_1_vc_sel_1_1 <= _GEN_195;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_vc_sel_0_0 <= io_vcalloc_resp_vc_sel_0_0; // @[InputUnit.scala 271:26]
      end else begin
        states_1_vc_sel_0_0 <= _GEN_198;
      end
    end else begin
      states_1_vc_sel_0_0 <= _GEN_198;
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h1 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_1_flow_ingress_node <= io_in_flit_0_bits_flow_ingress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h1 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_1_flow_egress_node <= io_in_flit_0_bits_flow_egress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (reset) begin // @[InputUnit.scala 377:23]
      states_2_g <= 3'h0; // @[InputUnit.scala 378:24]
    end else if (_T_64 & input_buffer_io_deq_2_bits_tail) begin // @[InputUnit.scala 292:35]
      states_2_g <= 3'h0; // @[InputUnit.scala 293:13]
    end else if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_g <= 3'h3; // @[InputUnit.scala 272:21]
      end else begin
        states_2_g <= _GEN_224;
      end
    end else begin
      states_2_g <= _GEN_224;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_2_0 <= io_vcalloc_resp_vc_sel_2_0; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_2_0 <= _GEN_202;
      end
    end else begin
      states_2_vc_sel_2_0 <= _GEN_202;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_1_0 <= io_vcalloc_resp_vc_sel_1_0; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_1_0 <= _GEN_203;
      end
    end else begin
      states_2_vc_sel_1_0 <= _GEN_203;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_1_1 <= io_vcalloc_resp_vc_sel_1_1; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_1_1 <= _GEN_204;
      end
    end else begin
      states_2_vc_sel_1_1 <= _GEN_204;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_1_2 <= io_vcalloc_resp_vc_sel_1_2; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_1_2 <= _GEN_205;
      end
    end else begin
      states_2_vc_sel_1_2 <= _GEN_205;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_0_0 <= io_vcalloc_resp_vc_sel_0_0; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_0_0 <= _GEN_207;
      end
    end else begin
      states_2_vc_sel_0_0 <= _GEN_207;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_0_1 <= io_vcalloc_resp_vc_sel_0_1; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_0_1 <= _GEN_208;
      end
    end else begin
      states_2_vc_sel_0_1 <= _GEN_208;
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h2 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_2_flow_ingress_node <= io_in_flit_0_bits_flow_ingress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h2 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_2_flow_egress_node <= io_in_flit_0_bits_flow_egress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (reset) begin // @[InputUnit.scala 377:23]
      states_3_g <= 3'h0; // @[InputUnit.scala 378:24]
    end else if (_T_66 & input_buffer_io_deq_3_bits_tail) begin // @[InputUnit.scala 292:35]
      states_3_g <= 3'h0; // @[InputUnit.scala 293:13]
    end else if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_g <= 3'h3; // @[InputUnit.scala 272:21]
      end else begin
        states_3_g <= _GEN_225;
      end
    end else begin
      states_3_g <= _GEN_225;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_2_0 <= io_vcalloc_resp_vc_sel_2_0; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_2_0 <= _GEN_211;
      end
    end else begin
      states_3_vc_sel_2_0 <= _GEN_211;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_1_0 <= io_vcalloc_resp_vc_sel_1_0; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_1_0 <= _GEN_212;
      end
    end else begin
      states_3_vc_sel_1_0 <= _GEN_212;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_1_1 <= io_vcalloc_resp_vc_sel_1_1; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_1_1 <= _GEN_213;
      end
    end else begin
      states_3_vc_sel_1_1 <= _GEN_213;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_1_2 <= io_vcalloc_resp_vc_sel_1_2; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_1_2 <= _GEN_214;
      end
    end else begin
      states_3_vc_sel_1_2 <= _GEN_214;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_1_3 <= io_vcalloc_resp_vc_sel_1_3; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_1_3 <= _GEN_215;
      end
    end else begin
      states_3_vc_sel_1_3 <= _GEN_215;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_0_0 <= io_vcalloc_resp_vc_sel_0_0; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_0_0 <= _GEN_216;
      end
    end else begin
      states_3_vc_sel_0_0 <= _GEN_216;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_0_1 <= io_vcalloc_resp_vc_sel_0_1; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_0_1 <= _GEN_217;
      end
    end else begin
      states_3_vc_sel_0_1 <= _GEN_217;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_0_2 <= io_vcalloc_resp_vc_sel_0_2; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_0_2 <= _GEN_218;
      end
    end else begin
      states_3_vc_sel_0_2 <= _GEN_218;
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h3 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_3_flow_ingress_node <= io_in_flit_0_bits_flow_ingress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h3 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_3_flow_egress_node <= io_in_flit_0_bits_flow_egress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (reset) begin // @[InputUnit.scala 233:21]
      mask <= 4'h0; // @[InputUnit.scala 233:21]
    end else if (io_router_req_valid) begin // @[InputUnit.scala 239:31]
      mask <= _mask_T_2; // @[InputUnit.scala 240:10]
    end else if (_T_26) begin // @[InputUnit.scala 241:34]
      mask <= _mask_T_17; // @[InputUnit.scala 242:10]
    end
    salloc_outs_0_valid <= salloc_arb_io_out_0_ready & salloc_arb_io_out_0_valid; // @[Decoupled.scala 51:35]
    salloc_outs_0_out_vid <= _virt_channel_T_10 | _virt_channel_T_11; // @[Mux.scala 27:73]
    salloc_outs_0_flit_head <= salloc_arb_io_chosen_oh_0[0] & input_buffer_io_deq_0_bits_head |
      salloc_arb_io_chosen_oh_0[1] & input_buffer_io_deq_1_bits_head | salloc_arb_io_chosen_oh_0[2] &
      input_buffer_io_deq_2_bits_head | salloc_arb_io_chosen_oh_0[3] & input_buffer_io_deq_3_bits_head; // @[Mux.scala 27:73]
    salloc_outs_0_flit_tail <= salloc_arb_io_chosen_oh_0[0] & input_buffer_io_deq_0_bits_tail |
      salloc_arb_io_chosen_oh_0[1] & input_buffer_io_deq_1_bits_tail | salloc_arb_io_chosen_oh_0[2] &
      input_buffer_io_deq_2_bits_tail | salloc_arb_io_chosen_oh_0[3] & input_buffer_io_deq_3_bits_tail; // @[Mux.scala 27:73]
    salloc_outs_0_flit_payload <= _salloc_outs_0_flit_payload_T_9 | _salloc_outs_0_flit_payload_T_7; // @[Mux.scala 27:73]
    salloc_outs_0_flit_flow_ingress_node <= _salloc_outs_0_flit_flow_T_30 | _salloc_outs_0_flit_flow_T_28; // @[Mux.scala 27:73]
    salloc_outs_0_flit_flow_egress_node <= _salloc_outs_0_flit_flow_T_16 | _salloc_outs_0_flit_flow_T_14; // @[Mux.scala 27:73]
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T & _T_3 & ~(_GEN_3 == 3'h0)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:197 assert(states(id).g === g_i)\n"); // @[InputUnit.scala 197:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_router_req_valid & _T_3 & ~(_GEN_139 == 3'h1)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:224 assert(states(id).g === g_r)\n"); // @[InputUnit.scala 224:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_39 & vcalloc_sel[0] & _T_3 & ~vcalloc_vals_0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:274 assert(states(i).g === g_v)\n"); // @[InputUnit.scala 274:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_39 & vcalloc_sel[1] & _T_3 & ~vcalloc_vals_1) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:274 assert(states(i).g === g_v)\n"); // @[InputUnit.scala 274:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_39 & vcalloc_sel[2] & _T_3 & ~vcalloc_vals_2) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:274 assert(states(i).g === g_v)\n"); // @[InputUnit.scala 274:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_39 & vcalloc_sel[3] & _T_3 & ~vcalloc_vals_3) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:274 assert(states(i).g === g_v)\n"); // @[InputUnit.scala 274:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  states_0_g = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  states_0_vc_sel_2_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  states_0_vc_sel_1_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  states_0_vc_sel_0_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  states_0_flow_ingress_node = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  states_0_flow_egress_node = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  states_1_g = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  states_1_vc_sel_2_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  states_1_vc_sel_1_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  states_1_vc_sel_1_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  states_1_vc_sel_0_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  states_1_flow_ingress_node = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  states_1_flow_egress_node = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  states_2_g = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  states_2_vc_sel_2_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  states_2_vc_sel_1_0 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  states_2_vc_sel_1_1 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  states_2_vc_sel_1_2 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  states_2_vc_sel_0_0 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  states_2_vc_sel_0_1 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  states_2_flow_ingress_node = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  states_2_flow_egress_node = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  states_3_g = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  states_3_vc_sel_2_0 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  states_3_vc_sel_1_0 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  states_3_vc_sel_1_1 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  states_3_vc_sel_1_2 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  states_3_vc_sel_1_3 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  states_3_vc_sel_0_0 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  states_3_vc_sel_0_1 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  states_3_vc_sel_0_2 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  states_3_flow_ingress_node = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  states_3_flow_egress_node = _RAND_32[1:0];
  _RAND_33 = {1{`RANDOM}};
  mask = _RAND_33[3:0];
  _RAND_34 = {1{`RANDOM}};
  salloc_outs_0_valid = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  salloc_outs_0_out_vid = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  salloc_outs_0_flit_head = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  salloc_outs_0_flit_tail = _RAND_37[0:0];
  _RAND_38 = {2{`RANDOM}};
  salloc_outs_0_flit_payload = _RAND_38[63:0];
  _RAND_39 = {1{`RANDOM}};
  salloc_outs_0_flit_flow_ingress_node = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  salloc_outs_0_flit_flow_egress_node = _RAND_40[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (_T & ~reset) begin
      assert(1'h1); // @[InputUnit.scala 196:13]
    end
    //
    if (_T & _T_3) begin
      assert(_GEN_3 == 3'h0); // @[InputUnit.scala 197:13]
    end
    //
    if (io_router_req_valid & _T_3) begin
      assert(_GEN_139 == 3'h1); // @[InputUnit.scala 224:11]
    end
    //
    if (_T_39 & vcalloc_sel[0] & _T_3) begin
      assert(vcalloc_vals_0); // @[InputUnit.scala 274:17]
    end
    //
    if (_T_39 & vcalloc_sel[1] & _T_3) begin
      assert(vcalloc_vals_1); // @[InputUnit.scala 274:17]
    end
    //
    if (_T_39 & vcalloc_sel[2] & _T_3) begin
      assert(vcalloc_vals_2); // @[InputUnit.scala 274:17]
    end
    //
    if (_T_39 & vcalloc_sel[3] & _T_3) begin
      assert(vcalloc_vals_3); // @[InputUnit.scala 274:17]
    end
  end
endmodule
module InputUnit_7(
  input         clock,
  input         reset,
  output        io_router_req_valid,
  output [1:0]  io_router_req_bits_src_virt_id,
  output [1:0]  io_router_req_bits_flow_ingress_node,
  output [1:0]  io_router_req_bits_flow_egress_node,
  input         io_router_resp_vc_sel_1_0,
  input         io_router_resp_vc_sel_1_1,
  input         io_router_resp_vc_sel_1_2,
  input         io_router_resp_vc_sel_1_3,
  input         io_router_resp_vc_sel_0_0,
  input         io_router_resp_vc_sel_0_1,
  input         io_router_resp_vc_sel_0_2,
  input         io_vcalloc_req_ready,
  output        io_vcalloc_req_valid,
  output        io_vcalloc_req_bits_vc_sel_2_0,
  output        io_vcalloc_req_bits_vc_sel_1_0,
  output        io_vcalloc_req_bits_vc_sel_1_1,
  output        io_vcalloc_req_bits_vc_sel_1_2,
  output        io_vcalloc_req_bits_vc_sel_1_3,
  output        io_vcalloc_req_bits_vc_sel_0_0,
  output        io_vcalloc_req_bits_vc_sel_0_1,
  output        io_vcalloc_req_bits_vc_sel_0_2,
  input         io_vcalloc_resp_vc_sel_2_0,
  input         io_vcalloc_resp_vc_sel_1_0,
  input         io_vcalloc_resp_vc_sel_1_1,
  input         io_vcalloc_resp_vc_sel_1_2,
  input         io_vcalloc_resp_vc_sel_1_3,
  input         io_vcalloc_resp_vc_sel_0_0,
  input         io_vcalloc_resp_vc_sel_0_1,
  input         io_vcalloc_resp_vc_sel_0_2,
  input         io_out_credit_available_2_0,
  input         io_out_credit_available_1_0,
  input         io_out_credit_available_1_1,
  input         io_out_credit_available_1_2,
  input         io_out_credit_available_1_3,
  input         io_out_credit_available_0_0,
  input         io_out_credit_available_0_1,
  input         io_out_credit_available_0_2,
  input         io_out_credit_available_0_3,
  input         io_salloc_req_0_ready,
  output        io_salloc_req_0_valid,
  output        io_salloc_req_0_bits_vc_sel_2_0,
  output        io_salloc_req_0_bits_vc_sel_1_0,
  output        io_salloc_req_0_bits_vc_sel_1_1,
  output        io_salloc_req_0_bits_vc_sel_1_2,
  output        io_salloc_req_0_bits_vc_sel_1_3,
  output        io_salloc_req_0_bits_vc_sel_0_0,
  output        io_salloc_req_0_bits_vc_sel_0_1,
  output        io_salloc_req_0_bits_vc_sel_0_2,
  output        io_salloc_req_0_bits_vc_sel_0_3,
  output        io_salloc_req_0_bits_tail,
  output        io_out_0_valid,
  output        io_out_0_bits_flit_head,
  output        io_out_0_bits_flit_tail,
  output [63:0] io_out_0_bits_flit_payload,
  output [1:0]  io_out_0_bits_flit_flow_ingress_node,
  output [1:0]  io_out_0_bits_flit_flow_egress_node,
  output [1:0]  io_out_0_bits_out_virt_channel,
  output [1:0]  io_debug_va_stall,
  output [1:0]  io_debug_sa_stall,
  input         io_in_flit_0_valid,
  input         io_in_flit_0_bits_head,
  input         io_in_flit_0_bits_tail,
  input  [63:0] io_in_flit_0_bits_payload,
  input  [1:0]  io_in_flit_0_bits_flow_ingress_node,
  input  [1:0]  io_in_flit_0_bits_flow_egress_node,
  input  [1:0]  io_in_flit_0_bits_virt_channel_id,
  output [3:0]  io_in_credit_return,
  output [3:0]  io_in_vc_free
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
`endif // RANDOMIZE_REG_INIT
  wire  input_buffer_clock; // @[InputUnit.scala 180:28]
  wire  input_buffer_reset; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_enq_0_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_enq_0_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_enq_0_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_enq_0_bits_payload; // @[InputUnit.scala 180:28]
  wire [1:0] input_buffer_io_enq_0_bits_virt_channel_id; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_0_ready; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_0_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_0_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_0_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_deq_0_bits_payload; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_ready; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_deq_1_bits_payload; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_ready; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_deq_2_bits_payload; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_3_ready; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_3_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_3_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_3_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_deq_3_bits_payload; // @[InputUnit.scala 180:28]
  wire  route_arbiter_io_in_0_valid; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_0_bits_flow_ingress_node; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_0_bits_flow_egress_node; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_1_ready; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_1_valid; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_1_bits_flow_ingress_node; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_1_bits_flow_egress_node; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_2_ready; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_2_valid; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_2_bits_flow_ingress_node; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_2_bits_flow_egress_node; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_3_ready; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_3_valid; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_3_bits_flow_ingress_node; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_in_3_bits_flow_egress_node; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_out_valid; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_out_bits_src_virt_id; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_out_bits_flow_ingress_node; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_out_bits_flow_egress_node; // @[InputUnit.scala 186:29]
  wire  salloc_arb_clock; // @[InputUnit.scala 279:26]
  wire  salloc_arb_reset; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_bits_vc_sel_2_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_bits_vc_sel_1_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_bits_tail; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_vc_sel_2_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_vc_sel_1_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_vc_sel_1_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_vc_sel_0_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_tail; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_2_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_1_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_1_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_1_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_0_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_0_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_tail; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_2_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_1_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_1_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_1_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_1_3; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_0_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_0_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_0_3; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_tail; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_2_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_1_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_1_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_1_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_1_3; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_0_1; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_0_2; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_0_3; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_tail; // @[InputUnit.scala 279:26]
  wire [3:0] salloc_arb_io_chosen_oh_0; // @[InputUnit.scala 279:26]
  reg [2:0] states_0_g; // @[InputUnit.scala 191:19]
  reg  states_0_vc_sel_2_0; // @[InputUnit.scala 191:19]
  reg  states_0_vc_sel_1_0; // @[InputUnit.scala 191:19]
  reg  states_0_vc_sel_0_0; // @[InputUnit.scala 191:19]
  reg [1:0] states_0_flow_ingress_node; // @[InputUnit.scala 191:19]
  reg [1:0] states_0_flow_egress_node; // @[InputUnit.scala 191:19]
  reg [2:0] states_1_g; // @[InputUnit.scala 191:19]
  reg  states_1_vc_sel_2_0; // @[InputUnit.scala 191:19]
  reg  states_1_vc_sel_1_1; // @[InputUnit.scala 191:19]
  reg  states_1_vc_sel_0_0; // @[InputUnit.scala 191:19]
  reg [1:0] states_1_flow_ingress_node; // @[InputUnit.scala 191:19]
  reg [1:0] states_1_flow_egress_node; // @[InputUnit.scala 191:19]
  reg [2:0] states_2_g; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_2_0; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_1_1; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_1_2; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_0_0; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_0_1; // @[InputUnit.scala 191:19]
  reg [1:0] states_2_flow_ingress_node; // @[InputUnit.scala 191:19]
  reg [1:0] states_2_flow_egress_node; // @[InputUnit.scala 191:19]
  reg [2:0] states_3_g; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_2_0; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_1_1; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_1_2; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_1_3; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_0_0; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_0_1; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_0_2; // @[InputUnit.scala 191:19]
  reg [1:0] states_3_flow_ingress_node; // @[InputUnit.scala 191:19]
  reg [1:0] states_3_flow_egress_node; // @[InputUnit.scala 191:19]
  wire  _T = io_in_flit_0_valid & io_in_flit_0_bits_head; // @[InputUnit.scala 194:32]
  wire  _T_3 = ~reset; // @[InputUnit.scala 196:13]
  wire [2:0] _GEN_1 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? states_1_g : states_0_g; // @[InputUnit.scala 197:{27,27}]
  wire [2:0] _GEN_2 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? states_2_g : _GEN_1; // @[InputUnit.scala 197:{27,27}]
  wire [2:0] _GEN_3 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? states_3_g : _GEN_2; // @[InputUnit.scala 197:{27,27}]
  wire  at_dest = io_in_flit_0_bits_flow_egress_node == 2'h3; // @[InputUnit.scala 198:57]
  wire [2:0] _states_g_T = at_dest ? 3'h2 : 3'h1; // @[InputUnit.scala 199:26]
  wire [2:0] _GEN_4 = 2'h0 == io_in_flit_0_bits_virt_channel_id ? _states_g_T : states_0_g; // @[InputUnit.scala 191:19 199:{20,20}]
  wire [2:0] _GEN_5 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? _states_g_T : states_1_g; // @[InputUnit.scala 191:19 199:{20,20}]
  wire [2:0] _GEN_6 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? _states_g_T : states_2_g; // @[InputUnit.scala 191:19 199:{20,20}]
  wire [2:0] _GEN_7 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? _states_g_T : states_3_g; // @[InputUnit.scala 191:19 199:{20,20}]
  wire  _GEN_8 = 2'h0 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_0_vc_sel_0_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_9 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_1_vc_sel_0_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_10 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_0_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_11 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_0_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_14 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_0_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_15 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_0_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_19 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_0_2; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_24 = 2'h0 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_0_vc_sel_1_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_29 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_1_vc_sel_1_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_30 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_1_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_31 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_1_1; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_34 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_1_2; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_35 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_1_2; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_39 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_1_3; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_40 = 2'h0 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_0_vc_sel_2_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_41 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_1_vc_sel_2_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_42 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_2_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_43 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_2_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_44 = 2'h0 == io_in_flit_0_bits_virt_channel_id | _GEN_40; // @[InputUnit.scala 203:{44,44}]
  wire  _GEN_45 = 2'h1 == io_in_flit_0_bits_virt_channel_id | _GEN_41; // @[InputUnit.scala 203:{44,44}]
  wire  _GEN_46 = 2'h2 == io_in_flit_0_bits_virt_channel_id | _GEN_42; // @[InputUnit.scala 203:{44,44}]
  wire  _GEN_47 = 2'h3 == io_in_flit_0_bits_virt_channel_id | _GEN_43; // @[InputUnit.scala 203:{44,44}]
  wire [2:0] _GEN_72 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_4 : states_0_g; // @[InputUnit.scala 191:19 194:60]
  wire [2:0] _GEN_73 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_5 : states_1_g; // @[InputUnit.scala 191:19 194:60]
  wire [2:0] _GEN_74 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_6 : states_2_g; // @[InputUnit.scala 191:19 194:60]
  wire [2:0] _GEN_75 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_7 : states_3_g; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_76 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_8 : states_0_vc_sel_0_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_77 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_9 : states_1_vc_sel_0_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_78 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_10 : states_2_vc_sel_0_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_79 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_11 : states_3_vc_sel_0_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_82 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_14 : states_2_vc_sel_0_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_83 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_15 : states_3_vc_sel_0_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_87 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_19 : states_3_vc_sel_0_2; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_92 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_24 : states_0_vc_sel_1_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_97 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_29 : states_1_vc_sel_1_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_98 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_30 : states_2_vc_sel_1_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_99 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_31 : states_3_vc_sel_1_1; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_102 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_34 : states_2_vc_sel_1_2; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_103 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_35 : states_3_vc_sel_1_2; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_107 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_39 : states_3_vc_sel_1_3; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_108 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_44 : states_0_vc_sel_2_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_109 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_45 : states_1_vc_sel_2_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_110 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_46 : states_2_vc_sel_2_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_111 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_47 : states_3_vc_sel_2_0; // @[InputUnit.scala 191:19 194:60]
  wire  _T_10 = route_arbiter_io_in_0_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_132 = _T_10 ? 3'h2 : _GEN_72; // @[InputUnit.scala 215:{23,29}]
  wire  _T_11 = route_arbiter_io_in_1_ready & route_arbiter_io_in_1_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_133 = _T_11 ? 3'h2 : _GEN_73; // @[InputUnit.scala 215:{23,29}]
  wire  _T_12 = route_arbiter_io_in_2_ready & route_arbiter_io_in_2_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_134 = _T_12 ? 3'h2 : _GEN_74; // @[InputUnit.scala 215:{23,29}]
  wire  _T_13 = route_arbiter_io_in_3_ready & route_arbiter_io_in_3_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_135 = _T_13 ? 3'h2 : _GEN_75; // @[InputUnit.scala 215:{23,29}]
  wire [2:0] _GEN_137 = 2'h1 == io_router_req_bits_src_virt_id ? states_1_g : states_0_g; // @[InputUnit.scala 224:{25,25}]
  wire [2:0] _GEN_138 = 2'h2 == io_router_req_bits_src_virt_id ? states_2_g : _GEN_137; // @[InputUnit.scala 224:{25,25}]
  wire [2:0] _GEN_139 = 2'h3 == io_router_req_bits_src_virt_id ? states_3_g : _GEN_138; // @[InputUnit.scala 224:{25,25}]
  wire [2:0] _GEN_140 = 2'h0 == io_router_req_bits_src_virt_id ? 3'h2 : _GEN_132; // @[InputUnit.scala 225:{18,18}]
  wire [2:0] _GEN_141 = 2'h1 == io_router_req_bits_src_virt_id ? 3'h2 : _GEN_133; // @[InputUnit.scala 225:{18,18}]
  wire [2:0] _GEN_142 = 2'h2 == io_router_req_bits_src_virt_id ? 3'h2 : _GEN_134; // @[InputUnit.scala 225:{18,18}]
  wire [2:0] _GEN_143 = 2'h3 == io_router_req_bits_src_virt_id ? 3'h2 : _GEN_135; // @[InputUnit.scala 225:{18,18}]
  wire  _GEN_144 = 2'h0 == io_router_req_bits_src_virt_id ? 1'h0 : _GEN_108; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_145 = 2'h0 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_0 : _GEN_92; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_149 = 2'h0 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_0 : _GEN_76; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_153 = 2'h1 == io_router_req_bits_src_virt_id ? 1'h0 : _GEN_109; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_155 = 2'h1 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_1 : _GEN_97; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_158 = 2'h1 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_0 : _GEN_77; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_162 = 2'h2 == io_router_req_bits_src_virt_id ? 1'h0 : _GEN_110; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_164 = 2'h2 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_1 : _GEN_98; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_165 = 2'h2 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_2 : _GEN_102; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_167 = 2'h2 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_0 : _GEN_78; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_168 = 2'h2 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_1 : _GEN_82; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_171 = 2'h3 == io_router_req_bits_src_virt_id ? 1'h0 : _GEN_111; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_173 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_1 : _GEN_99; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_174 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_2 : _GEN_103; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_175 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_1_3 : _GEN_107; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_176 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_0 : _GEN_79; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_177 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_1 : _GEN_83; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_178 = 2'h3 == io_router_req_bits_src_virt_id ? io_router_resp_vc_sel_0_2 : _GEN_87; // @[InputUnit.scala 227:25 228:26]
  wire [2:0] _GEN_180 = io_router_req_valid ? _GEN_140 : _GEN_132; // @[InputUnit.scala 222:31]
  wire [2:0] _GEN_181 = io_router_req_valid ? _GEN_141 : _GEN_133; // @[InputUnit.scala 222:31]
  wire [2:0] _GEN_182 = io_router_req_valid ? _GEN_142 : _GEN_134; // @[InputUnit.scala 222:31]
  wire [2:0] _GEN_183 = io_router_req_valid ? _GEN_143 : _GEN_135; // @[InputUnit.scala 222:31]
  wire  _GEN_184 = io_router_req_valid ? _GEN_144 : _GEN_108; // @[InputUnit.scala 222:31]
  wire  _GEN_185 = io_router_req_valid ? _GEN_145 : _GEN_92; // @[InputUnit.scala 222:31]
  wire  _GEN_189 = io_router_req_valid ? _GEN_149 : _GEN_76; // @[InputUnit.scala 222:31]
  wire  _GEN_193 = io_router_req_valid ? _GEN_153 : _GEN_109; // @[InputUnit.scala 222:31]
  wire  _GEN_195 = io_router_req_valid ? _GEN_155 : _GEN_97; // @[InputUnit.scala 222:31]
  wire  _GEN_198 = io_router_req_valid ? _GEN_158 : _GEN_77; // @[InputUnit.scala 222:31]
  wire  _GEN_202 = io_router_req_valid ? _GEN_162 : _GEN_110; // @[InputUnit.scala 222:31]
  wire  _GEN_204 = io_router_req_valid ? _GEN_164 : _GEN_98; // @[InputUnit.scala 222:31]
  wire  _GEN_205 = io_router_req_valid ? _GEN_165 : _GEN_102; // @[InputUnit.scala 222:31]
  wire  _GEN_207 = io_router_req_valid ? _GEN_167 : _GEN_78; // @[InputUnit.scala 222:31]
  wire  _GEN_208 = io_router_req_valid ? _GEN_168 : _GEN_82; // @[InputUnit.scala 222:31]
  wire  _GEN_211 = io_router_req_valid ? _GEN_171 : _GEN_111; // @[InputUnit.scala 222:31]
  wire  _GEN_213 = io_router_req_valid ? _GEN_173 : _GEN_99; // @[InputUnit.scala 222:31]
  wire  _GEN_214 = io_router_req_valid ? _GEN_174 : _GEN_103; // @[InputUnit.scala 222:31]
  wire  _GEN_215 = io_router_req_valid ? _GEN_175 : _GEN_107; // @[InputUnit.scala 222:31]
  wire  _GEN_216 = io_router_req_valid ? _GEN_176 : _GEN_79; // @[InputUnit.scala 222:31]
  wire  _GEN_217 = io_router_req_valid ? _GEN_177 : _GEN_83; // @[InputUnit.scala 222:31]
  wire  _GEN_218 = io_router_req_valid ? _GEN_178 : _GEN_87; // @[InputUnit.scala 222:31]
  reg [3:0] mask; // @[InputUnit.scala 233:21]
  wire  vcalloc_vals_1 = states_1_g == 3'h2; // @[InputUnit.scala 249:32]
  wire  vcalloc_vals_0 = states_0_g == 3'h2; // @[InputUnit.scala 249:32]
  wire  vcalloc_vals_3 = states_3_g == 3'h2; // @[InputUnit.scala 249:32]
  wire  vcalloc_vals_2 = states_2_g == 3'h2; // @[InputUnit.scala 249:32]
  wire [3:0] _vcalloc_filter_T = {vcalloc_vals_3,vcalloc_vals_2,vcalloc_vals_1,vcalloc_vals_0}; // @[InputUnit.scala 236:59]
  wire [3:0] _vcalloc_filter_T_2 = ~mask; // @[InputUnit.scala 236:89]
  wire [3:0] _vcalloc_filter_T_3 = _vcalloc_filter_T & _vcalloc_filter_T_2; // @[InputUnit.scala 236:87]
  wire [7:0] _vcalloc_filter_T_4 = {vcalloc_vals_3,vcalloc_vals_2,vcalloc_vals_1,vcalloc_vals_0,_vcalloc_filter_T_3}; // @[Cat.scala 33:92]
  wire [7:0] _vcalloc_filter_T_13 = _vcalloc_filter_T_4[7] ? 8'h80 : 8'h0; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_14 = _vcalloc_filter_T_4[6] ? 8'h40 : _vcalloc_filter_T_13; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_15 = _vcalloc_filter_T_4[5] ? 8'h20 : _vcalloc_filter_T_14; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_16 = _vcalloc_filter_T_4[4] ? 8'h10 : _vcalloc_filter_T_15; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_17 = _vcalloc_filter_T_4[3] ? 8'h8 : _vcalloc_filter_T_16; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_18 = _vcalloc_filter_T_4[2] ? 8'h4 : _vcalloc_filter_T_17; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_19 = _vcalloc_filter_T_4[1] ? 8'h2 : _vcalloc_filter_T_18; // @[Mux.scala 47:70]
  wire [7:0] vcalloc_filter = _vcalloc_filter_T_4[0] ? 8'h1 : _vcalloc_filter_T_19; // @[Mux.scala 47:70]
  wire [3:0] vcalloc_sel = vcalloc_filter[3:0] | vcalloc_filter[7:4]; // @[InputUnit.scala 237:58]
  wire [3:0] _mask_T = 4'h1 << io_router_req_bits_src_virt_id; // @[InputUnit.scala 240:18]
  wire [3:0] _mask_T_2 = _mask_T - 4'h1; // @[InputUnit.scala 240:53]
  wire  _T_26 = vcalloc_vals_0 | vcalloc_vals_1 | vcalloc_vals_2 | vcalloc_vals_3; // @[package.scala 73:59]
  wire [1:0] _mask_T_12 = vcalloc_sel[1] ? 2'h3 : 2'h0; // @[Mux.scala 27:73]
  wire [2:0] _mask_T_13 = vcalloc_sel[2] ? 3'h7 : 3'h0; // @[Mux.scala 27:73]
  wire [3:0] _mask_T_14 = vcalloc_sel[3] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [1:0] _GEN_60 = {{1'd0}, vcalloc_sel[0]}; // @[Mux.scala 27:73]
  wire [1:0] _mask_T_15 = _GEN_60 | _mask_T_12; // @[Mux.scala 27:73]
  wire [2:0] _GEN_61 = {{1'd0}, _mask_T_15}; // @[Mux.scala 27:73]
  wire [2:0] _mask_T_16 = _GEN_61 | _mask_T_13; // @[Mux.scala 27:73]
  wire [3:0] _GEN_62 = {{1'd0}, _mask_T_16}; // @[Mux.scala 27:73]
  wire [3:0] _mask_T_17 = _GEN_62 | _mask_T_14; // @[Mux.scala 27:73]
  wire [2:0] _GEN_222 = vcalloc_vals_0 & vcalloc_sel[0] & io_vcalloc_req_ready ? 3'h3 : _GEN_180; // @[InputUnit.scala 253:{76,82}]
  wire [2:0] _GEN_223 = vcalloc_vals_1 & vcalloc_sel[1] & io_vcalloc_req_ready ? 3'h3 : _GEN_181; // @[InputUnit.scala 253:{76,82}]
  wire [2:0] _GEN_224 = vcalloc_vals_2 & vcalloc_sel[2] & io_vcalloc_req_ready ? 3'h3 : _GEN_182; // @[InputUnit.scala 253:{76,82}]
  wire [2:0] _GEN_225 = vcalloc_vals_3 & vcalloc_sel[3] & io_vcalloc_req_ready ? 3'h3 : _GEN_183; // @[InputUnit.scala 253:{76,82}]
  wire [1:0] _io_debug_va_stall_T = vcalloc_vals_0 + vcalloc_vals_1; // @[Bitwise.scala 51:90]
  wire [1:0] _io_debug_va_stall_T_2 = vcalloc_vals_2 + vcalloc_vals_3; // @[Bitwise.scala 51:90]
  wire [2:0] _io_debug_va_stall_T_4 = _io_debug_va_stall_T + _io_debug_va_stall_T_2; // @[Bitwise.scala 51:90]
  wire [2:0] _GEN_63 = {{2'd0}, io_vcalloc_req_ready}; // @[InputUnit.scala 266:47]
  wire [2:0] _io_debug_va_stall_T_7 = _io_debug_va_stall_T_4 - _GEN_63; // @[InputUnit.scala 266:47]
  wire  _T_39 = io_vcalloc_req_ready & io_vcalloc_req_valid; // @[Decoupled.scala 51:35]
  wire [8:0] _credit_available_T = {states_0_vc_sel_2_0,1'h0,1'h0,1'h0,states_0_vc_sel_1_0,2'h0,1'h0,states_0_vc_sel_0_0
    }; // @[InputUnit.scala 287:40]
  wire [8:0] _credit_available_T_1 = {io_out_credit_available_2_0,io_out_credit_available_1_3,
    io_out_credit_available_1_2,io_out_credit_available_1_1,io_out_credit_available_1_0,io_out_credit_available_0_3,
    io_out_credit_available_0_2,io_out_credit_available_0_1,io_out_credit_available_0_0}; // @[InputUnit.scala 287:73]
  wire [8:0] _credit_available_T_2 = _credit_available_T & _credit_available_T_1; // @[InputUnit.scala 287:47]
  wire  credit_available = _credit_available_T_2 != 9'h0; // @[InputUnit.scala 287:81]
  wire  _T_60 = salloc_arb_io_in_0_ready & salloc_arb_io_in_0_valid; // @[Decoupled.scala 51:35]
  wire [8:0] _credit_available_T_3 = {states_1_vc_sel_2_0,1'h0,1'h0,states_1_vc_sel_1_1,1'h0,2'h0,1'h0,
    states_1_vc_sel_0_0}; // @[InputUnit.scala 287:40]
  wire [8:0] _credit_available_T_5 = _credit_available_T_3 & _credit_available_T_1; // @[InputUnit.scala 287:47]
  wire  credit_available_1 = _credit_available_T_5 != 9'h0; // @[InputUnit.scala 287:81]
  wire  _T_62 = salloc_arb_io_in_1_ready & salloc_arb_io_in_1_valid; // @[Decoupled.scala 51:35]
  wire [8:0] _credit_available_T_6 = {states_2_vc_sel_2_0,1'h0,states_2_vc_sel_1_2,states_2_vc_sel_1_1,1'h0,2'h0,
    states_2_vc_sel_0_1,states_2_vc_sel_0_0}; // @[InputUnit.scala 287:40]
  wire [8:0] _credit_available_T_8 = _credit_available_T_6 & _credit_available_T_1; // @[InputUnit.scala 287:47]
  wire  credit_available_2 = _credit_available_T_8 != 9'h0; // @[InputUnit.scala 287:81]
  wire  _T_64 = salloc_arb_io_in_2_ready & salloc_arb_io_in_2_valid; // @[Decoupled.scala 51:35]
  wire [8:0] _credit_available_T_9 = {states_3_vc_sel_2_0,states_3_vc_sel_1_3,states_3_vc_sel_1_2,states_3_vc_sel_1_1,1'h0
    ,1'h0,states_3_vc_sel_0_2,states_3_vc_sel_0_1,states_3_vc_sel_0_0}; // @[InputUnit.scala 287:40]
  wire [8:0] _credit_available_T_11 = _credit_available_T_9 & _credit_available_T_1; // @[InputUnit.scala 287:47]
  wire  credit_available_3 = _credit_available_T_11 != 9'h0; // @[InputUnit.scala 287:81]
  wire  _T_66 = salloc_arb_io_in_3_ready & salloc_arb_io_in_3_valid; // @[Decoupled.scala 51:35]
  wire  _io_debug_sa_stall_T_1 = salloc_arb_io_in_0_valid & ~salloc_arb_io_in_0_ready; // @[InputUnit.scala 301:67]
  wire  _io_debug_sa_stall_T_3 = salloc_arb_io_in_1_valid & ~salloc_arb_io_in_1_ready; // @[InputUnit.scala 301:67]
  wire  _io_debug_sa_stall_T_5 = salloc_arb_io_in_2_valid & ~salloc_arb_io_in_2_ready; // @[InputUnit.scala 301:67]
  wire  _io_debug_sa_stall_T_7 = salloc_arb_io_in_3_valid & ~salloc_arb_io_in_3_ready; // @[InputUnit.scala 301:67]
  wire [1:0] _io_debug_sa_stall_T_8 = _io_debug_sa_stall_T_1 + _io_debug_sa_stall_T_3; // @[Bitwise.scala 51:90]
  wire [1:0] _io_debug_sa_stall_T_10 = _io_debug_sa_stall_T_5 + _io_debug_sa_stall_T_7; // @[Bitwise.scala 51:90]
  wire [2:0] _io_debug_sa_stall_T_12 = _io_debug_sa_stall_T_8 + _io_debug_sa_stall_T_10; // @[Bitwise.scala 51:90]
  reg  salloc_outs_0_valid; // @[InputUnit.scala 318:8]
  reg [1:0] salloc_outs_0_out_vid; // @[InputUnit.scala 318:8]
  reg  salloc_outs_0_flit_head; // @[InputUnit.scala 318:8]
  reg  salloc_outs_0_flit_tail; // @[InputUnit.scala 318:8]
  reg [63:0] salloc_outs_0_flit_payload; // @[InputUnit.scala 318:8]
  reg [1:0] salloc_outs_0_flit_flow_ingress_node; // @[InputUnit.scala 318:8]
  reg [1:0] salloc_outs_0_flit_flow_egress_node; // @[InputUnit.scala 318:8]
  wire  _io_in_credit_return_T = salloc_arb_io_out_0_ready & salloc_arb_io_out_0_valid; // @[Decoupled.scala 51:35]
  wire  _io_in_vc_free_T_11 = salloc_arb_io_chosen_oh_0[0] & input_buffer_io_deq_0_bits_tail | salloc_arb_io_chosen_oh_0
    [1] & input_buffer_io_deq_1_bits_tail | salloc_arb_io_chosen_oh_0[2] & input_buffer_io_deq_2_bits_tail |
    salloc_arb_io_chosen_oh_0[3] & input_buffer_io_deq_3_bits_tail; // @[Mux.scala 27:73]
  wire  vc_sel_0_0 = salloc_arb_io_chosen_oh_0[0] & states_0_vc_sel_0_0 | salloc_arb_io_chosen_oh_0[1] &
    states_1_vc_sel_0_0 | salloc_arb_io_chosen_oh_0[2] & states_2_vc_sel_0_0 | salloc_arb_io_chosen_oh_0[3] &
    states_3_vc_sel_0_0; // @[Mux.scala 27:73]
  wire  vc_sel_0_1 = salloc_arb_io_chosen_oh_0[2] & states_2_vc_sel_0_1 | salloc_arb_io_chosen_oh_0[3] &
    states_3_vc_sel_0_1; // @[Mux.scala 27:73]
  wire  vc_sel_0_2 = salloc_arb_io_chosen_oh_0[3] & states_3_vc_sel_0_2; // @[Mux.scala 27:73]
  wire  vc_sel_1_0 = salloc_arb_io_chosen_oh_0[0] & states_0_vc_sel_1_0; // @[Mux.scala 27:73]
  wire  vc_sel_1_1 = salloc_arb_io_chosen_oh_0[1] & states_1_vc_sel_1_1 | salloc_arb_io_chosen_oh_0[2] &
    states_2_vc_sel_1_1 | salloc_arb_io_chosen_oh_0[3] & states_3_vc_sel_1_1; // @[Mux.scala 27:73]
  wire  vc_sel_1_2 = salloc_arb_io_chosen_oh_0[2] & states_2_vc_sel_1_2 | salloc_arb_io_chosen_oh_0[3] &
    states_3_vc_sel_1_2; // @[Mux.scala 27:73]
  wire  vc_sel_1_3 = salloc_arb_io_chosen_oh_0[3] & states_3_vc_sel_1_3; // @[Mux.scala 27:73]
  wire  channel_oh_0 = vc_sel_0_0 | vc_sel_0_1 | vc_sel_0_2; // @[InputUnit.scala 334:43]
  wire  channel_oh_1 = vc_sel_1_0 | vc_sel_1_1 | vc_sel_1_2 | vc_sel_1_3; // @[InputUnit.scala 334:43]
  wire [3:0] _virt_channel_T = {1'h0,vc_sel_0_2,vc_sel_0_1,vc_sel_0_0}; // @[OneHot.scala 22:45]
  wire [1:0] virt_channel_hi_1 = _virt_channel_T[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] virt_channel_lo_1 = _virt_channel_T[1:0]; // @[OneHot.scala 31:18]
  wire  _virt_channel_T_1 = |virt_channel_hi_1; // @[OneHot.scala 32:14]
  wire [1:0] _virt_channel_T_2 = virt_channel_hi_1 | virt_channel_lo_1; // @[OneHot.scala 32:28]
  wire [1:0] _virt_channel_T_4 = {_virt_channel_T_1,_virt_channel_T_2[1]}; // @[Cat.scala 33:92]
  wire [3:0] _virt_channel_T_5 = {vc_sel_1_3,vc_sel_1_2,vc_sel_1_1,vc_sel_1_0}; // @[OneHot.scala 22:45]
  wire [1:0] virt_channel_hi_3 = _virt_channel_T_5[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] virt_channel_lo_3 = _virt_channel_T_5[1:0]; // @[OneHot.scala 31:18]
  wire  _virt_channel_T_6 = |virt_channel_hi_3; // @[OneHot.scala 32:14]
  wire [1:0] _virt_channel_T_7 = virt_channel_hi_3 | virt_channel_lo_3; // @[OneHot.scala 32:28]
  wire [1:0] _virt_channel_T_9 = {_virt_channel_T_6,_virt_channel_T_7[1]}; // @[Cat.scala 33:92]
  wire [1:0] _virt_channel_T_10 = channel_oh_0 ? _virt_channel_T_4 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _virt_channel_T_11 = channel_oh_1 ? _virt_channel_T_9 : 2'h0; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_4 = salloc_arb_io_chosen_oh_0[0] ? input_buffer_io_deq_0_bits_payload : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_5 = salloc_arb_io_chosen_oh_0[1] ? input_buffer_io_deq_1_bits_payload : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_6 = salloc_arb_io_chosen_oh_0[2] ? input_buffer_io_deq_2_bits_payload : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_7 = salloc_arb_io_chosen_oh_0[3] ? input_buffer_io_deq_3_bits_payload : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_8 = _salloc_outs_0_flit_payload_T_4 | _salloc_outs_0_flit_payload_T_5; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_9 = _salloc_outs_0_flit_payload_T_8 | _salloc_outs_0_flit_payload_T_6; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_11 = salloc_arb_io_chosen_oh_0[0] ? states_0_flow_egress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_12 = salloc_arb_io_chosen_oh_0[1] ? states_1_flow_egress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_13 = salloc_arb_io_chosen_oh_0[2] ? states_2_flow_egress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_14 = salloc_arb_io_chosen_oh_0[3] ? states_3_flow_egress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_15 = _salloc_outs_0_flit_flow_T_11 | _salloc_outs_0_flit_flow_T_12; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_16 = _salloc_outs_0_flit_flow_T_15 | _salloc_outs_0_flit_flow_T_13; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_25 = salloc_arb_io_chosen_oh_0[0] ? states_0_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_26 = salloc_arb_io_chosen_oh_0[1] ? states_1_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_27 = salloc_arb_io_chosen_oh_0[2] ? states_2_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_28 = salloc_arb_io_chosen_oh_0[3] ? states_3_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_29 = _salloc_outs_0_flit_flow_T_25 | _salloc_outs_0_flit_flow_T_26; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_30 = _salloc_outs_0_flit_flow_T_29 | _salloc_outs_0_flit_flow_T_27; // @[Mux.scala 27:73]
  InputBuffer input_buffer ( // @[InputUnit.scala 180:28]
    .clock(input_buffer_clock),
    .reset(input_buffer_reset),
    .io_enq_0_valid(input_buffer_io_enq_0_valid),
    .io_enq_0_bits_head(input_buffer_io_enq_0_bits_head),
    .io_enq_0_bits_tail(input_buffer_io_enq_0_bits_tail),
    .io_enq_0_bits_payload(input_buffer_io_enq_0_bits_payload),
    .io_enq_0_bits_virt_channel_id(input_buffer_io_enq_0_bits_virt_channel_id),
    .io_deq_0_ready(input_buffer_io_deq_0_ready),
    .io_deq_0_valid(input_buffer_io_deq_0_valid),
    .io_deq_0_bits_head(input_buffer_io_deq_0_bits_head),
    .io_deq_0_bits_tail(input_buffer_io_deq_0_bits_tail),
    .io_deq_0_bits_payload(input_buffer_io_deq_0_bits_payload),
    .io_deq_1_ready(input_buffer_io_deq_1_ready),
    .io_deq_1_valid(input_buffer_io_deq_1_valid),
    .io_deq_1_bits_head(input_buffer_io_deq_1_bits_head),
    .io_deq_1_bits_tail(input_buffer_io_deq_1_bits_tail),
    .io_deq_1_bits_payload(input_buffer_io_deq_1_bits_payload),
    .io_deq_2_ready(input_buffer_io_deq_2_ready),
    .io_deq_2_valid(input_buffer_io_deq_2_valid),
    .io_deq_2_bits_head(input_buffer_io_deq_2_bits_head),
    .io_deq_2_bits_tail(input_buffer_io_deq_2_bits_tail),
    .io_deq_2_bits_payload(input_buffer_io_deq_2_bits_payload),
    .io_deq_3_ready(input_buffer_io_deq_3_ready),
    .io_deq_3_valid(input_buffer_io_deq_3_valid),
    .io_deq_3_bits_head(input_buffer_io_deq_3_bits_head),
    .io_deq_3_bits_tail(input_buffer_io_deq_3_bits_tail),
    .io_deq_3_bits_payload(input_buffer_io_deq_3_bits_payload)
  );
  Arbiter route_arbiter ( // @[InputUnit.scala 186:29]
    .io_in_0_valid(route_arbiter_io_in_0_valid),
    .io_in_0_bits_flow_ingress_node(route_arbiter_io_in_0_bits_flow_ingress_node),
    .io_in_0_bits_flow_egress_node(route_arbiter_io_in_0_bits_flow_egress_node),
    .io_in_1_ready(route_arbiter_io_in_1_ready),
    .io_in_1_valid(route_arbiter_io_in_1_valid),
    .io_in_1_bits_flow_ingress_node(route_arbiter_io_in_1_bits_flow_ingress_node),
    .io_in_1_bits_flow_egress_node(route_arbiter_io_in_1_bits_flow_egress_node),
    .io_in_2_ready(route_arbiter_io_in_2_ready),
    .io_in_2_valid(route_arbiter_io_in_2_valid),
    .io_in_2_bits_flow_ingress_node(route_arbiter_io_in_2_bits_flow_ingress_node),
    .io_in_2_bits_flow_egress_node(route_arbiter_io_in_2_bits_flow_egress_node),
    .io_in_3_ready(route_arbiter_io_in_3_ready),
    .io_in_3_valid(route_arbiter_io_in_3_valid),
    .io_in_3_bits_flow_ingress_node(route_arbiter_io_in_3_bits_flow_ingress_node),
    .io_in_3_bits_flow_egress_node(route_arbiter_io_in_3_bits_flow_egress_node),
    .io_out_valid(route_arbiter_io_out_valid),
    .io_out_bits_src_virt_id(route_arbiter_io_out_bits_src_virt_id),
    .io_out_bits_flow_ingress_node(route_arbiter_io_out_bits_flow_ingress_node),
    .io_out_bits_flow_egress_node(route_arbiter_io_out_bits_flow_egress_node)
  );
  SwitchArbiter salloc_arb ( // @[InputUnit.scala 279:26]
    .clock(salloc_arb_clock),
    .reset(salloc_arb_reset),
    .io_in_0_ready(salloc_arb_io_in_0_ready),
    .io_in_0_valid(salloc_arb_io_in_0_valid),
    .io_in_0_bits_vc_sel_2_0(salloc_arb_io_in_0_bits_vc_sel_2_0),
    .io_in_0_bits_vc_sel_1_0(salloc_arb_io_in_0_bits_vc_sel_1_0),
    .io_in_0_bits_vc_sel_0_0(salloc_arb_io_in_0_bits_vc_sel_0_0),
    .io_in_0_bits_tail(salloc_arb_io_in_0_bits_tail),
    .io_in_1_ready(salloc_arb_io_in_1_ready),
    .io_in_1_valid(salloc_arb_io_in_1_valid),
    .io_in_1_bits_vc_sel_2_0(salloc_arb_io_in_1_bits_vc_sel_2_0),
    .io_in_1_bits_vc_sel_1_0(salloc_arb_io_in_1_bits_vc_sel_1_0),
    .io_in_1_bits_vc_sel_1_1(salloc_arb_io_in_1_bits_vc_sel_1_1),
    .io_in_1_bits_vc_sel_0_0(salloc_arb_io_in_1_bits_vc_sel_0_0),
    .io_in_1_bits_vc_sel_0_1(salloc_arb_io_in_1_bits_vc_sel_0_1),
    .io_in_1_bits_tail(salloc_arb_io_in_1_bits_tail),
    .io_in_2_ready(salloc_arb_io_in_2_ready),
    .io_in_2_valid(salloc_arb_io_in_2_valid),
    .io_in_2_bits_vc_sel_2_0(salloc_arb_io_in_2_bits_vc_sel_2_0),
    .io_in_2_bits_vc_sel_1_0(salloc_arb_io_in_2_bits_vc_sel_1_0),
    .io_in_2_bits_vc_sel_1_1(salloc_arb_io_in_2_bits_vc_sel_1_1),
    .io_in_2_bits_vc_sel_1_2(salloc_arb_io_in_2_bits_vc_sel_1_2),
    .io_in_2_bits_vc_sel_0_0(salloc_arb_io_in_2_bits_vc_sel_0_0),
    .io_in_2_bits_vc_sel_0_1(salloc_arb_io_in_2_bits_vc_sel_0_1),
    .io_in_2_bits_vc_sel_0_2(salloc_arb_io_in_2_bits_vc_sel_0_2),
    .io_in_2_bits_tail(salloc_arb_io_in_2_bits_tail),
    .io_in_3_ready(salloc_arb_io_in_3_ready),
    .io_in_3_valid(salloc_arb_io_in_3_valid),
    .io_in_3_bits_vc_sel_2_0(salloc_arb_io_in_3_bits_vc_sel_2_0),
    .io_in_3_bits_vc_sel_1_0(salloc_arb_io_in_3_bits_vc_sel_1_0),
    .io_in_3_bits_vc_sel_1_1(salloc_arb_io_in_3_bits_vc_sel_1_1),
    .io_in_3_bits_vc_sel_1_2(salloc_arb_io_in_3_bits_vc_sel_1_2),
    .io_in_3_bits_vc_sel_1_3(salloc_arb_io_in_3_bits_vc_sel_1_3),
    .io_in_3_bits_vc_sel_0_0(salloc_arb_io_in_3_bits_vc_sel_0_0),
    .io_in_3_bits_vc_sel_0_1(salloc_arb_io_in_3_bits_vc_sel_0_1),
    .io_in_3_bits_vc_sel_0_2(salloc_arb_io_in_3_bits_vc_sel_0_2),
    .io_in_3_bits_vc_sel_0_3(salloc_arb_io_in_3_bits_vc_sel_0_3),
    .io_in_3_bits_tail(salloc_arb_io_in_3_bits_tail),
    .io_out_0_ready(salloc_arb_io_out_0_ready),
    .io_out_0_valid(salloc_arb_io_out_0_valid),
    .io_out_0_bits_vc_sel_2_0(salloc_arb_io_out_0_bits_vc_sel_2_0),
    .io_out_0_bits_vc_sel_1_0(salloc_arb_io_out_0_bits_vc_sel_1_0),
    .io_out_0_bits_vc_sel_1_1(salloc_arb_io_out_0_bits_vc_sel_1_1),
    .io_out_0_bits_vc_sel_1_2(salloc_arb_io_out_0_bits_vc_sel_1_2),
    .io_out_0_bits_vc_sel_1_3(salloc_arb_io_out_0_bits_vc_sel_1_3),
    .io_out_0_bits_vc_sel_0_0(salloc_arb_io_out_0_bits_vc_sel_0_0),
    .io_out_0_bits_vc_sel_0_1(salloc_arb_io_out_0_bits_vc_sel_0_1),
    .io_out_0_bits_vc_sel_0_2(salloc_arb_io_out_0_bits_vc_sel_0_2),
    .io_out_0_bits_vc_sel_0_3(salloc_arb_io_out_0_bits_vc_sel_0_3),
    .io_out_0_bits_tail(salloc_arb_io_out_0_bits_tail),
    .io_chosen_oh_0(salloc_arb_io_chosen_oh_0)
  );
  assign io_router_req_valid = route_arbiter_io_out_valid; // @[InputUnit.scala 189:17]
  assign io_router_req_bits_src_virt_id = route_arbiter_io_out_bits_src_virt_id; // @[InputUnit.scala 189:17]
  assign io_router_req_bits_flow_ingress_node = route_arbiter_io_out_bits_flow_ingress_node; // @[InputUnit.scala 189:17]
  assign io_router_req_bits_flow_egress_node = route_arbiter_io_out_bits_flow_egress_node; // @[InputUnit.scala 189:17]
  assign io_vcalloc_req_valid = vcalloc_vals_0 | vcalloc_vals_1 | vcalloc_vals_2 | vcalloc_vals_3; // @[package.scala 73:59]
  assign io_vcalloc_req_bits_vc_sel_2_0 = vcalloc_sel[0] & states_0_vc_sel_2_0 | vcalloc_sel[1] & states_1_vc_sel_2_0 |
    vcalloc_sel[2] & states_2_vc_sel_2_0 | vcalloc_sel[3] & states_3_vc_sel_2_0; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_1_0 = vcalloc_sel[0] & states_0_vc_sel_1_0; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_1_1 = vcalloc_sel[1] & states_1_vc_sel_1_1 | vcalloc_sel[2] & states_2_vc_sel_1_1 |
    vcalloc_sel[3] & states_3_vc_sel_1_1; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_1_2 = vcalloc_sel[2] & states_2_vc_sel_1_2 | vcalloc_sel[3] & states_3_vc_sel_1_2; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_1_3 = vcalloc_sel[3] & states_3_vc_sel_1_3; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_0_0 = vcalloc_sel[0] & states_0_vc_sel_0_0 | vcalloc_sel[1] & states_1_vc_sel_0_0 |
    vcalloc_sel[2] & states_2_vc_sel_0_0 | vcalloc_sel[3] & states_3_vc_sel_0_0; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_0_1 = vcalloc_sel[2] & states_2_vc_sel_0_1 | vcalloc_sel[3] & states_3_vc_sel_0_1; // @[Mux.scala 27:73]
  assign io_vcalloc_req_bits_vc_sel_0_2 = vcalloc_sel[3] & states_3_vc_sel_0_2; // @[Mux.scala 27:73]
  assign io_salloc_req_0_valid = salloc_arb_io_out_0_valid; // @[InputUnit.scala 302:17 303:19 305:35]
  assign io_salloc_req_0_bits_vc_sel_2_0 = salloc_arb_io_out_0_bits_vc_sel_2_0; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_1_0 = salloc_arb_io_out_0_bits_vc_sel_1_0; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_1_1 = salloc_arb_io_out_0_bits_vc_sel_1_1; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_1_2 = salloc_arb_io_out_0_bits_vc_sel_1_2; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_1_3 = salloc_arb_io_out_0_bits_vc_sel_1_3; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_0_0 = salloc_arb_io_out_0_bits_vc_sel_0_0; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_0_1 = salloc_arb_io_out_0_bits_vc_sel_0_1; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_0_2 = salloc_arb_io_out_0_bits_vc_sel_0_2; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_vc_sel_0_3 = salloc_arb_io_out_0_bits_vc_sel_0_3; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_tail = salloc_arb_io_out_0_bits_tail; // @[InputUnit.scala 302:17]
  assign io_out_0_valid = salloc_outs_0_valid; // @[InputUnit.scala 349:21]
  assign io_out_0_bits_flit_head = salloc_outs_0_flit_head; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_flit_tail = salloc_outs_0_flit_tail; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_flit_payload = salloc_outs_0_flit_payload; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_flit_flow_ingress_node = salloc_outs_0_flit_flow_ingress_node; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_flit_flow_egress_node = salloc_outs_0_flit_flow_egress_node; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_out_virt_channel = salloc_outs_0_out_vid; // @[InputUnit.scala 351:37]
  assign io_debug_va_stall = _io_debug_va_stall_T_7[1:0]; // @[InputUnit.scala 266:21]
  assign io_debug_sa_stall = _io_debug_sa_stall_T_12[1:0]; // @[InputUnit.scala 301:21]
  assign io_in_credit_return = _io_in_credit_return_T ? salloc_arb_io_chosen_oh_0 : 4'h0; // @[InputUnit.scala 322:8]
  assign io_in_vc_free = _io_in_credit_return_T & _io_in_vc_free_T_11 ? salloc_arb_io_chosen_oh_0 : 4'h0; // @[InputUnit.scala 325:8]
  assign input_buffer_clock = clock;
  assign input_buffer_reset = reset;
  assign input_buffer_io_enq_0_valid = io_in_flit_0_valid; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_head = io_in_flit_0_bits_head; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_tail = io_in_flit_0_bits_tail; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_payload = io_in_flit_0_bits_payload; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_virt_channel_id = io_in_flit_0_bits_virt_channel_id; // @[InputUnit.scala 182:28]
  assign input_buffer_io_deq_0_ready = salloc_arb_io_in_0_ready; // @[InputUnit.scala 295:36]
  assign input_buffer_io_deq_1_ready = salloc_arb_io_in_1_ready; // @[InputUnit.scala 295:36]
  assign input_buffer_io_deq_2_ready = salloc_arb_io_in_2_ready; // @[InputUnit.scala 295:36]
  assign input_buffer_io_deq_3_ready = salloc_arb_io_in_3_ready; // @[InputUnit.scala 295:36]
  assign route_arbiter_io_in_0_valid = states_0_g == 3'h1; // @[InputUnit.scala 212:22]
  assign route_arbiter_io_in_0_bits_flow_ingress_node = states_0_flow_ingress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_0_bits_flow_egress_node = states_0_flow_egress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_1_valid = states_1_g == 3'h1; // @[InputUnit.scala 212:22]
  assign route_arbiter_io_in_1_bits_flow_ingress_node = states_1_flow_ingress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_1_bits_flow_egress_node = states_1_flow_egress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_2_valid = states_2_g == 3'h1; // @[InputUnit.scala 212:22]
  assign route_arbiter_io_in_2_bits_flow_ingress_node = states_2_flow_ingress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_2_bits_flow_egress_node = states_2_flow_egress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_3_valid = states_3_g == 3'h1; // @[InputUnit.scala 212:22]
  assign route_arbiter_io_in_3_bits_flow_ingress_node = states_3_flow_ingress_node; // @[InputUnit.scala 213:19]
  assign route_arbiter_io_in_3_bits_flow_egress_node = states_3_flow_egress_node; // @[InputUnit.scala 213:19]
  assign salloc_arb_clock = clock;
  assign salloc_arb_reset = reset;
  assign salloc_arb_io_in_0_valid = states_0_g == 3'h3 & credit_available & input_buffer_io_deq_0_valid; // @[InputUnit.scala 288:50]
  assign salloc_arb_io_in_0_bits_vc_sel_2_0 = states_0_vc_sel_2_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_0_bits_vc_sel_1_0 = states_0_vc_sel_1_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_0_bits_vc_sel_0_0 = states_0_vc_sel_0_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_0_bits_tail = input_buffer_io_deq_0_bits_tail; // @[InputUnit.scala 291:19]
  assign salloc_arb_io_in_1_valid = states_1_g == 3'h3 & credit_available_1 & input_buffer_io_deq_1_valid; // @[InputUnit.scala 288:50]
  assign salloc_arb_io_in_1_bits_vc_sel_2_0 = states_1_vc_sel_2_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_1_bits_vc_sel_1_0 = 1'h0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_1_bits_vc_sel_1_1 = states_1_vc_sel_1_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_1_bits_vc_sel_0_0 = states_1_vc_sel_0_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_1_bits_vc_sel_0_1 = 1'h0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_1_bits_tail = input_buffer_io_deq_1_bits_tail; // @[InputUnit.scala 291:19]
  assign salloc_arb_io_in_2_valid = states_2_g == 3'h3 & credit_available_2 & input_buffer_io_deq_2_valid; // @[InputUnit.scala 288:50]
  assign salloc_arb_io_in_2_bits_vc_sel_2_0 = states_2_vc_sel_2_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_1_0 = 1'h0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_1_1 = states_2_vc_sel_1_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_1_2 = states_2_vc_sel_1_2; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_0_0 = states_2_vc_sel_0_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_0_1 = states_2_vc_sel_0_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_vc_sel_0_2 = 1'h0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_tail = input_buffer_io_deq_2_bits_tail; // @[InputUnit.scala 291:19]
  assign salloc_arb_io_in_3_valid = states_3_g == 3'h3 & credit_available_3 & input_buffer_io_deq_3_valid; // @[InputUnit.scala 288:50]
  assign salloc_arb_io_in_3_bits_vc_sel_2_0 = states_3_vc_sel_2_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_1_0 = 1'h0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_1_1 = states_3_vc_sel_1_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_1_2 = states_3_vc_sel_1_2; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_1_3 = states_3_vc_sel_1_3; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_0_0 = states_3_vc_sel_0_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_0_1 = states_3_vc_sel_0_1; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_0_2 = states_3_vc_sel_0_2; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_vc_sel_0_3 = 1'h0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_tail = input_buffer_io_deq_3_bits_tail; // @[InputUnit.scala 291:19]
  assign salloc_arb_io_out_0_ready = io_salloc_req_0_ready; // @[InputUnit.scala 302:17 303:19 304:39]
  always @(posedge clock) begin
    if (reset) begin // @[InputUnit.scala 377:23]
      states_0_g <= 3'h0; // @[InputUnit.scala 378:24]
    end else if (_T_60 & input_buffer_io_deq_0_bits_tail) begin // @[InputUnit.scala 292:35]
      states_0_g <= 3'h0; // @[InputUnit.scala 293:13]
    end else if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[0]) begin // @[InputUnit.scala 270:29]
        states_0_g <= 3'h3; // @[InputUnit.scala 272:21]
      end else begin
        states_0_g <= _GEN_222;
      end
    end else begin
      states_0_g <= _GEN_222;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[0]) begin // @[InputUnit.scala 270:29]
        states_0_vc_sel_2_0 <= io_vcalloc_resp_vc_sel_2_0; // @[InputUnit.scala 271:26]
      end else begin
        states_0_vc_sel_2_0 <= _GEN_184;
      end
    end else begin
      states_0_vc_sel_2_0 <= _GEN_184;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[0]) begin // @[InputUnit.scala 270:29]
        states_0_vc_sel_1_0 <= io_vcalloc_resp_vc_sel_1_0; // @[InputUnit.scala 271:26]
      end else begin
        states_0_vc_sel_1_0 <= _GEN_185;
      end
    end else begin
      states_0_vc_sel_1_0 <= _GEN_185;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[0]) begin // @[InputUnit.scala 270:29]
        states_0_vc_sel_0_0 <= io_vcalloc_resp_vc_sel_0_0; // @[InputUnit.scala 271:26]
      end else begin
        states_0_vc_sel_0_0 <= _GEN_189;
      end
    end else begin
      states_0_vc_sel_0_0 <= _GEN_189;
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h0 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_0_flow_ingress_node <= io_in_flit_0_bits_flow_ingress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h0 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_0_flow_egress_node <= io_in_flit_0_bits_flow_egress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (reset) begin // @[InputUnit.scala 377:23]
      states_1_g <= 3'h0; // @[InputUnit.scala 378:24]
    end else if (_T_62 & input_buffer_io_deq_1_bits_tail) begin // @[InputUnit.scala 292:35]
      states_1_g <= 3'h0; // @[InputUnit.scala 293:13]
    end else if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_g <= 3'h3; // @[InputUnit.scala 272:21]
      end else begin
        states_1_g <= _GEN_223;
      end
    end else begin
      states_1_g <= _GEN_223;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_vc_sel_2_0 <= io_vcalloc_resp_vc_sel_2_0; // @[InputUnit.scala 271:26]
      end else begin
        states_1_vc_sel_2_0 <= _GEN_193;
      end
    end else begin
      states_1_vc_sel_2_0 <= _GEN_193;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_vc_sel_1_1 <= io_vcalloc_resp_vc_sel_1_1; // @[InputUnit.scala 271:26]
      end else begin
        states_1_vc_sel_1_1 <= _GEN_195;
      end
    end else begin
      states_1_vc_sel_1_1 <= _GEN_195;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_vc_sel_0_0 <= io_vcalloc_resp_vc_sel_0_0; // @[InputUnit.scala 271:26]
      end else begin
        states_1_vc_sel_0_0 <= _GEN_198;
      end
    end else begin
      states_1_vc_sel_0_0 <= _GEN_198;
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h1 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_1_flow_ingress_node <= io_in_flit_0_bits_flow_ingress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h1 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_1_flow_egress_node <= io_in_flit_0_bits_flow_egress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (reset) begin // @[InputUnit.scala 377:23]
      states_2_g <= 3'h0; // @[InputUnit.scala 378:24]
    end else if (_T_64 & input_buffer_io_deq_2_bits_tail) begin // @[InputUnit.scala 292:35]
      states_2_g <= 3'h0; // @[InputUnit.scala 293:13]
    end else if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_g <= 3'h3; // @[InputUnit.scala 272:21]
      end else begin
        states_2_g <= _GEN_224;
      end
    end else begin
      states_2_g <= _GEN_224;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_2_0 <= io_vcalloc_resp_vc_sel_2_0; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_2_0 <= _GEN_202;
      end
    end else begin
      states_2_vc_sel_2_0 <= _GEN_202;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_1_1 <= io_vcalloc_resp_vc_sel_1_1; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_1_1 <= _GEN_204;
      end
    end else begin
      states_2_vc_sel_1_1 <= _GEN_204;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_1_2 <= io_vcalloc_resp_vc_sel_1_2; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_1_2 <= _GEN_205;
      end
    end else begin
      states_2_vc_sel_1_2 <= _GEN_205;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_0_0 <= io_vcalloc_resp_vc_sel_0_0; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_0_0 <= _GEN_207;
      end
    end else begin
      states_2_vc_sel_0_0 <= _GEN_207;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_0_1 <= io_vcalloc_resp_vc_sel_0_1; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_0_1 <= _GEN_208;
      end
    end else begin
      states_2_vc_sel_0_1 <= _GEN_208;
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h2 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_2_flow_ingress_node <= io_in_flit_0_bits_flow_ingress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h2 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_2_flow_egress_node <= io_in_flit_0_bits_flow_egress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (reset) begin // @[InputUnit.scala 377:23]
      states_3_g <= 3'h0; // @[InputUnit.scala 378:24]
    end else if (_T_66 & input_buffer_io_deq_3_bits_tail) begin // @[InputUnit.scala 292:35]
      states_3_g <= 3'h0; // @[InputUnit.scala 293:13]
    end else if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_g <= 3'h3; // @[InputUnit.scala 272:21]
      end else begin
        states_3_g <= _GEN_225;
      end
    end else begin
      states_3_g <= _GEN_225;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_2_0 <= io_vcalloc_resp_vc_sel_2_0; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_2_0 <= _GEN_211;
      end
    end else begin
      states_3_vc_sel_2_0 <= _GEN_211;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_1_1 <= io_vcalloc_resp_vc_sel_1_1; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_1_1 <= _GEN_213;
      end
    end else begin
      states_3_vc_sel_1_1 <= _GEN_213;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_1_2 <= io_vcalloc_resp_vc_sel_1_2; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_1_2 <= _GEN_214;
      end
    end else begin
      states_3_vc_sel_1_2 <= _GEN_214;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_1_3 <= io_vcalloc_resp_vc_sel_1_3; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_1_3 <= _GEN_215;
      end
    end else begin
      states_3_vc_sel_1_3 <= _GEN_215;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_0_0 <= io_vcalloc_resp_vc_sel_0_0; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_0_0 <= _GEN_216;
      end
    end else begin
      states_3_vc_sel_0_0 <= _GEN_216;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_0_1 <= io_vcalloc_resp_vc_sel_0_1; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_0_1 <= _GEN_217;
      end
    end else begin
      states_3_vc_sel_0_1 <= _GEN_217;
    end
    if (_T_39) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_0_2 <= io_vcalloc_resp_vc_sel_0_2; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_0_2 <= _GEN_218;
      end
    end else begin
      states_3_vc_sel_0_2 <= _GEN_218;
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h3 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_3_flow_ingress_node <= io_in_flit_0_bits_flow_ingress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h3 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_3_flow_egress_node <= io_in_flit_0_bits_flow_egress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (reset) begin // @[InputUnit.scala 233:21]
      mask <= 4'h0; // @[InputUnit.scala 233:21]
    end else if (io_router_req_valid) begin // @[InputUnit.scala 239:31]
      mask <= _mask_T_2; // @[InputUnit.scala 240:10]
    end else if (_T_26) begin // @[InputUnit.scala 241:34]
      mask <= _mask_T_17; // @[InputUnit.scala 242:10]
    end
    salloc_outs_0_valid <= salloc_arb_io_out_0_ready & salloc_arb_io_out_0_valid; // @[Decoupled.scala 51:35]
    salloc_outs_0_out_vid <= _virt_channel_T_10 | _virt_channel_T_11; // @[Mux.scala 27:73]
    salloc_outs_0_flit_head <= salloc_arb_io_chosen_oh_0[0] & input_buffer_io_deq_0_bits_head |
      salloc_arb_io_chosen_oh_0[1] & input_buffer_io_deq_1_bits_head | salloc_arb_io_chosen_oh_0[2] &
      input_buffer_io_deq_2_bits_head | salloc_arb_io_chosen_oh_0[3] & input_buffer_io_deq_3_bits_head; // @[Mux.scala 27:73]
    salloc_outs_0_flit_tail <= salloc_arb_io_chosen_oh_0[0] & input_buffer_io_deq_0_bits_tail |
      salloc_arb_io_chosen_oh_0[1] & input_buffer_io_deq_1_bits_tail | salloc_arb_io_chosen_oh_0[2] &
      input_buffer_io_deq_2_bits_tail | salloc_arb_io_chosen_oh_0[3] & input_buffer_io_deq_3_bits_tail; // @[Mux.scala 27:73]
    salloc_outs_0_flit_payload <= _salloc_outs_0_flit_payload_T_9 | _salloc_outs_0_flit_payload_T_7; // @[Mux.scala 27:73]
    salloc_outs_0_flit_flow_ingress_node <= _salloc_outs_0_flit_flow_T_30 | _salloc_outs_0_flit_flow_T_28; // @[Mux.scala 27:73]
    salloc_outs_0_flit_flow_egress_node <= _salloc_outs_0_flit_flow_T_16 | _salloc_outs_0_flit_flow_T_14; // @[Mux.scala 27:73]
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T & _T_3 & ~(_GEN_3 == 3'h0)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:197 assert(states(id).g === g_i)\n"); // @[InputUnit.scala 197:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_router_req_valid & _T_3 & ~(_GEN_139 == 3'h1)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:224 assert(states(id).g === g_r)\n"); // @[InputUnit.scala 224:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_39 & vcalloc_sel[0] & _T_3 & ~vcalloc_vals_0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:274 assert(states(i).g === g_v)\n"); // @[InputUnit.scala 274:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_39 & vcalloc_sel[1] & _T_3 & ~vcalloc_vals_1) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:274 assert(states(i).g === g_v)\n"); // @[InputUnit.scala 274:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_39 & vcalloc_sel[2] & _T_3 & ~vcalloc_vals_2) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:274 assert(states(i).g === g_v)\n"); // @[InputUnit.scala 274:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_39 & vcalloc_sel[3] & _T_3 & ~vcalloc_vals_3) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:274 assert(states(i).g === g_v)\n"); // @[InputUnit.scala 274:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  states_0_g = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  states_0_vc_sel_2_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  states_0_vc_sel_1_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  states_0_vc_sel_0_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  states_0_flow_ingress_node = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  states_0_flow_egress_node = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  states_1_g = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  states_1_vc_sel_2_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  states_1_vc_sel_1_1 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  states_1_vc_sel_0_0 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  states_1_flow_ingress_node = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  states_1_flow_egress_node = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  states_2_g = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  states_2_vc_sel_2_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  states_2_vc_sel_1_1 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  states_2_vc_sel_1_2 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  states_2_vc_sel_0_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  states_2_vc_sel_0_1 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  states_2_flow_ingress_node = _RAND_18[1:0];
  _RAND_19 = {1{`RANDOM}};
  states_2_flow_egress_node = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  states_3_g = _RAND_20[2:0];
  _RAND_21 = {1{`RANDOM}};
  states_3_vc_sel_2_0 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  states_3_vc_sel_1_1 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  states_3_vc_sel_1_2 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  states_3_vc_sel_1_3 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  states_3_vc_sel_0_0 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  states_3_vc_sel_0_1 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  states_3_vc_sel_0_2 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  states_3_flow_ingress_node = _RAND_28[1:0];
  _RAND_29 = {1{`RANDOM}};
  states_3_flow_egress_node = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  mask = _RAND_30[3:0];
  _RAND_31 = {1{`RANDOM}};
  salloc_outs_0_valid = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  salloc_outs_0_out_vid = _RAND_32[1:0];
  _RAND_33 = {1{`RANDOM}};
  salloc_outs_0_flit_head = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  salloc_outs_0_flit_tail = _RAND_34[0:0];
  _RAND_35 = {2{`RANDOM}};
  salloc_outs_0_flit_payload = _RAND_35[63:0];
  _RAND_36 = {1{`RANDOM}};
  salloc_outs_0_flit_flow_ingress_node = _RAND_36[1:0];
  _RAND_37 = {1{`RANDOM}};
  salloc_outs_0_flit_flow_egress_node = _RAND_37[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (_T & ~reset) begin
      assert(1'h1); // @[InputUnit.scala 196:13]
    end
    //
    if (_T & _T_3) begin
      assert(_GEN_3 == 3'h0); // @[InputUnit.scala 197:13]
    end
    //
    if (io_router_req_valid & _T_3) begin
      assert(_GEN_139 == 3'h1); // @[InputUnit.scala 224:11]
    end
    //
    if (_T_39 & vcalloc_sel[0] & _T_3) begin
      assert(vcalloc_vals_0); // @[InputUnit.scala 274:17]
    end
    //
    if (_T_39 & vcalloc_sel[1] & _T_3) begin
      assert(vcalloc_vals_1); // @[InputUnit.scala 274:17]
    end
    //
    if (_T_39 & vcalloc_sel[2] & _T_3) begin
      assert(vcalloc_vals_2); // @[InputUnit.scala 274:17]
    end
    //
    if (_T_39 & vcalloc_sel[3] & _T_3) begin
      assert(vcalloc_vals_3); // @[InputUnit.scala 274:17]
    end
  end
endmodule
module IngressUnit_3(
  input         clock,
  input         reset,
  output        io_router_req_valid,
  output [1:0]  io_router_req_bits_flow_ingress_node,
  output [1:0]  io_router_req_bits_flow_egress_node,
  input         io_router_resp_vc_sel_1_0,
  input         io_router_resp_vc_sel_1_1,
  input         io_router_resp_vc_sel_1_2,
  input         io_router_resp_vc_sel_1_3,
  input         io_router_resp_vc_sel_0_0,
  input         io_router_resp_vc_sel_0_1,
  input         io_router_resp_vc_sel_0_2,
  input         io_router_resp_vc_sel_0_3,
  input         io_vcalloc_req_ready,
  output        io_vcalloc_req_valid,
  output        io_vcalloc_req_bits_vc_sel_2_0,
  output        io_vcalloc_req_bits_vc_sel_1_0,
  output        io_vcalloc_req_bits_vc_sel_1_1,
  output        io_vcalloc_req_bits_vc_sel_1_2,
  output        io_vcalloc_req_bits_vc_sel_1_3,
  output        io_vcalloc_req_bits_vc_sel_0_0,
  output        io_vcalloc_req_bits_vc_sel_0_1,
  output        io_vcalloc_req_bits_vc_sel_0_2,
  output        io_vcalloc_req_bits_vc_sel_0_3,
  input         io_vcalloc_resp_vc_sel_2_0,
  input         io_vcalloc_resp_vc_sel_1_0,
  input         io_vcalloc_resp_vc_sel_1_1,
  input         io_vcalloc_resp_vc_sel_1_2,
  input         io_vcalloc_resp_vc_sel_1_3,
  input         io_vcalloc_resp_vc_sel_0_0,
  input         io_vcalloc_resp_vc_sel_0_1,
  input         io_vcalloc_resp_vc_sel_0_2,
  input         io_vcalloc_resp_vc_sel_0_3,
  input         io_out_credit_available_2_0,
  input         io_out_credit_available_1_0,
  input         io_out_credit_available_1_1,
  input         io_out_credit_available_1_2,
  input         io_out_credit_available_1_3,
  input         io_out_credit_available_0_0,
  input         io_out_credit_available_0_1,
  input         io_out_credit_available_0_2,
  input         io_out_credit_available_0_3,
  input         io_salloc_req_0_ready,
  output        io_salloc_req_0_valid,
  output        io_salloc_req_0_bits_vc_sel_2_0,
  output        io_salloc_req_0_bits_vc_sel_1_0,
  output        io_salloc_req_0_bits_vc_sel_1_1,
  output        io_salloc_req_0_bits_vc_sel_1_2,
  output        io_salloc_req_0_bits_vc_sel_1_3,
  output        io_salloc_req_0_bits_vc_sel_0_0,
  output        io_salloc_req_0_bits_vc_sel_0_1,
  output        io_salloc_req_0_bits_vc_sel_0_2,
  output        io_salloc_req_0_bits_vc_sel_0_3,
  output        io_salloc_req_0_bits_tail,
  output        io_out_0_valid,
  output        io_out_0_bits_flit_head,
  output        io_out_0_bits_flit_tail,
  output [63:0] io_out_0_bits_flit_payload,
  output [1:0]  io_out_0_bits_flit_flow_ingress_node,
  output [1:0]  io_out_0_bits_flit_flow_egress_node,
  output [1:0]  io_out_0_bits_out_virt_channel,
  output        io_in_ready,
  input         io_in_valid,
  input         io_in_bits_head,
  input         io_in_bits_tail,
  input  [63:0] io_in_bits_payload,
  input  [1:0]  io_in_bits_egress_id
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  route_buffer_clock; // @[IngressUnit.scala 26:28]
  wire  route_buffer_reset; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_enq_ready; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_enq_valid; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_enq_bits_head; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_enq_bits_tail; // @[IngressUnit.scala 26:28]
  wire [63:0] route_buffer_io_enq_bits_payload; // @[IngressUnit.scala 26:28]
  wire [1:0] route_buffer_io_enq_bits_flow_ingress_node; // @[IngressUnit.scala 26:28]
  wire [1:0] route_buffer_io_enq_bits_flow_egress_node; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_deq_ready; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_deq_valid; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_deq_bits_head; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_deq_bits_tail; // @[IngressUnit.scala 26:28]
  wire [63:0] route_buffer_io_deq_bits_payload; // @[IngressUnit.scala 26:28]
  wire [1:0] route_buffer_io_deq_bits_flow_ingress_node; // @[IngressUnit.scala 26:28]
  wire [1:0] route_buffer_io_deq_bits_flow_egress_node; // @[IngressUnit.scala 26:28]
  wire  route_q_clock; // @[IngressUnit.scala 27:23]
  wire  route_q_reset; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_ready; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_valid; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_2_0; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_1_0; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_1_1; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_1_2; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_1_3; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_0_0; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_0_1; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_0_2; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_0_3; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_ready; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_valid; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_2_0; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_1_0; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_1_1; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_1_2; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_1_3; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_0_0; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_0_1; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_0_2; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_0_3; // @[IngressUnit.scala 27:23]
  wire  vcalloc_buffer_clock; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_reset; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_enq_ready; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_enq_valid; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_enq_bits_head; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_enq_bits_tail; // @[IngressUnit.scala 75:30]
  wire [63:0] vcalloc_buffer_io_enq_bits_payload; // @[IngressUnit.scala 75:30]
  wire [1:0] vcalloc_buffer_io_enq_bits_flow_ingress_node; // @[IngressUnit.scala 75:30]
  wire [1:0] vcalloc_buffer_io_enq_bits_flow_egress_node; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_deq_ready; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_deq_valid; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_deq_bits_head; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_deq_bits_tail; // @[IngressUnit.scala 75:30]
  wire [63:0] vcalloc_buffer_io_deq_bits_payload; // @[IngressUnit.scala 75:30]
  wire [1:0] vcalloc_buffer_io_deq_bits_flow_ingress_node; // @[IngressUnit.scala 75:30]
  wire [1:0] vcalloc_buffer_io_deq_bits_flow_egress_node; // @[IngressUnit.scala 75:30]
  wire  vcalloc_q_clock; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_reset; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_ready; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_valid; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_2_0; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_1_0; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_1_1; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_1_2; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_1_3; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_0_0; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_0_1; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_0_2; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_0_3; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_ready; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_valid; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_2_0; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_1_0; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_1_1; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_1_2; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_1_3; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_0_0; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_0_1; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_0_2; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_0_3; // @[IngressUnit.scala 76:25]
  wire  _T = 2'h0 == io_in_bits_egress_id; // @[IngressUnit.scala 30:72]
  wire  _T_1 = 2'h1 == io_in_bits_egress_id; // @[IngressUnit.scala 30:72]
  wire  _T_2 = 2'h2 == io_in_bits_egress_id; // @[IngressUnit.scala 30:72]
  wire  _T_3 = 2'h3 == io_in_bits_egress_id; // @[IngressUnit.scala 30:72]
  wire  _T_6 = _T | _T_1 | _T_2 | _T_3; // @[package.scala 73:59]
  wire  _T_11 = ~reset; // @[IngressUnit.scala 30:9]
  wire [1:0] _route_buffer_io_enq_bits_flow_egress_node_T_6 = _T_2 ? 2'h2 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _route_buffer_io_enq_bits_flow_egress_node_T_7 = _T_3 ? 2'h3 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _GEN_11 = {{1'd0}, _T_1}; // @[Mux.scala 27:73]
  wire [1:0] _route_buffer_io_enq_bits_flow_egress_node_T_9 = _GEN_11 | _route_buffer_io_enq_bits_flow_egress_node_T_6; // @[Mux.scala 27:73]
  wire  at_dest = route_buffer_io_enq_bits_flow_egress_node == 2'h3; // @[IngressUnit.scala 55:59]
  wire  _T_13 = io_in_ready & io_in_valid; // @[Decoupled.scala 51:35]
  wire  _vcalloc_buffer_io_enq_valid_T = ~route_buffer_io_deq_bits_head; // @[IngressUnit.scala 88:30]
  wire  _vcalloc_buffer_io_enq_valid_T_1 = route_q_io_deq_valid | ~route_buffer_io_deq_bits_head; // @[IngressUnit.scala 88:27]
  wire  _vcalloc_buffer_io_enq_valid_T_2 = route_buffer_io_deq_valid & _vcalloc_buffer_io_enq_valid_T_1; // @[IngressUnit.scala 87:61]
  wire  _vcalloc_buffer_io_enq_valid_T_4 = io_vcalloc_req_ready | _vcalloc_buffer_io_enq_valid_T; // @[IngressUnit.scala 89:27]
  wire  _io_vcalloc_req_valid_T_1 = route_buffer_io_deq_valid & route_q_io_deq_valid & route_buffer_io_deq_bits_head; // @[IngressUnit.scala 91:78]
  wire  _route_buffer_io_deq_ready_T_2 = vcalloc_buffer_io_enq_ready & _vcalloc_buffer_io_enq_valid_T_1; // @[IngressUnit.scala 93:61]
  wire  _route_buffer_io_deq_ready_T_5 = _route_buffer_io_deq_ready_T_2 & _vcalloc_buffer_io_enq_valid_T_4; // @[IngressUnit.scala 94:37]
  wire  _route_buffer_io_deq_ready_T_7 = vcalloc_q_io_enq_ready | _vcalloc_buffer_io_enq_valid_T; // @[IngressUnit.scala 96:29]
  wire  _route_q_io_deq_ready_T = route_buffer_io_deq_ready & route_buffer_io_deq_valid; // @[Decoupled.scala 51:35]
  wire [3:0] c_lo = {vcalloc_q_io_deq_bits_vc_sel_0_3,vcalloc_q_io_deq_bits_vc_sel_0_2,vcalloc_q_io_deq_bits_vc_sel_0_1,
    vcalloc_q_io_deq_bits_vc_sel_0_0}; // @[IngressUnit.scala 107:41]
  wire [8:0] _c_T = {vcalloc_q_io_deq_bits_vc_sel_2_0,vcalloc_q_io_deq_bits_vc_sel_1_3,vcalloc_q_io_deq_bits_vc_sel_1_2,
    vcalloc_q_io_deq_bits_vc_sel_1_1,vcalloc_q_io_deq_bits_vc_sel_1_0,vcalloc_q_io_deq_bits_vc_sel_0_3,
    vcalloc_q_io_deq_bits_vc_sel_0_2,vcalloc_q_io_deq_bits_vc_sel_0_1,vcalloc_q_io_deq_bits_vc_sel_0_0}; // @[IngressUnit.scala 107:41]
  wire [8:0] _c_T_1 = {io_out_credit_available_2_0,io_out_credit_available_1_3,io_out_credit_available_1_2,
    io_out_credit_available_1_1,io_out_credit_available_1_0,io_out_credit_available_0_3,io_out_credit_available_0_2,
    io_out_credit_available_0_1,io_out_credit_available_0_0}; // @[IngressUnit.scala 107:74]
  wire [8:0] _c_T_2 = _c_T & _c_T_1; // @[IngressUnit.scala 107:48]
  wire  c = _c_T_2 != 9'h0; // @[IngressUnit.scala 107:82]
  wire  _vcalloc_q_io_deq_ready_T = vcalloc_buffer_io_deq_ready & vcalloc_buffer_io_deq_valid; // @[Decoupled.scala 51:35]
  reg  out_bundle_valid; // @[IngressUnit.scala 116:8]
  reg  out_bundle_bits_flit_head; // @[IngressUnit.scala 116:8]
  reg  out_bundle_bits_flit_tail; // @[IngressUnit.scala 116:8]
  reg [63:0] out_bundle_bits_flit_payload; // @[IngressUnit.scala 116:8]
  reg [1:0] out_bundle_bits_flit_flow_ingress_node; // @[IngressUnit.scala 116:8]
  reg [1:0] out_bundle_bits_flit_flow_egress_node; // @[IngressUnit.scala 116:8]
  reg [1:0] out_bundle_bits_out_virt_channel; // @[IngressUnit.scala 116:8]
  wire  out_channel_oh_0 = vcalloc_q_io_deq_bits_vc_sel_0_0 | vcalloc_q_io_deq_bits_vc_sel_0_1 |
    vcalloc_q_io_deq_bits_vc_sel_0_2 | vcalloc_q_io_deq_bits_vc_sel_0_3; // @[IngressUnit.scala 123:67]
  wire  out_channel_oh_1 = vcalloc_q_io_deq_bits_vc_sel_1_0 | vcalloc_q_io_deq_bits_vc_sel_1_1 |
    vcalloc_q_io_deq_bits_vc_sel_1_2 | vcalloc_q_io_deq_bits_vc_sel_1_3; // @[IngressUnit.scala 123:67]
  wire [1:0] out_bundle_bits_out_virt_channel_hi_1 = c_lo[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] out_bundle_bits_out_virt_channel_lo_1 = c_lo[1:0]; // @[OneHot.scala 31:18]
  wire  _out_bundle_bits_out_virt_channel_T_1 = |out_bundle_bits_out_virt_channel_hi_1; // @[OneHot.scala 32:14]
  wire [1:0] _out_bundle_bits_out_virt_channel_T_2 = out_bundle_bits_out_virt_channel_hi_1 |
    out_bundle_bits_out_virt_channel_lo_1; // @[OneHot.scala 32:28]
  wire [1:0] _out_bundle_bits_out_virt_channel_T_4 = {_out_bundle_bits_out_virt_channel_T_1,
    _out_bundle_bits_out_virt_channel_T_2[1]}; // @[Cat.scala 33:92]
  wire [3:0] _out_bundle_bits_out_virt_channel_T_5 = {vcalloc_q_io_deq_bits_vc_sel_1_3,vcalloc_q_io_deq_bits_vc_sel_1_2,
    vcalloc_q_io_deq_bits_vc_sel_1_1,vcalloc_q_io_deq_bits_vc_sel_1_0}; // @[OneHot.scala 22:45]
  wire [1:0] out_bundle_bits_out_virt_channel_hi_3 = _out_bundle_bits_out_virt_channel_T_5[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] out_bundle_bits_out_virt_channel_lo_3 = _out_bundle_bits_out_virt_channel_T_5[1:0]; // @[OneHot.scala 31:18]
  wire  _out_bundle_bits_out_virt_channel_T_6 = |out_bundle_bits_out_virt_channel_hi_3; // @[OneHot.scala 32:14]
  wire [1:0] _out_bundle_bits_out_virt_channel_T_7 = out_bundle_bits_out_virt_channel_hi_3 |
    out_bundle_bits_out_virt_channel_lo_3; // @[OneHot.scala 32:28]
  wire [1:0] _out_bundle_bits_out_virt_channel_T_9 = {_out_bundle_bits_out_virt_channel_T_6,
    _out_bundle_bits_out_virt_channel_T_7[1]}; // @[Cat.scala 33:92]
  wire [1:0] _out_bundle_bits_out_virt_channel_T_10 = out_channel_oh_0 ? _out_bundle_bits_out_virt_channel_T_4 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _out_bundle_bits_out_virt_channel_T_11 = out_channel_oh_1 ? _out_bundle_bits_out_virt_channel_T_9 : 2'h0; // @[Mux.scala 27:73]
  Queue_8 route_buffer ( // @[IngressUnit.scala 26:28]
    .clock(route_buffer_clock),
    .reset(route_buffer_reset),
    .io_enq_ready(route_buffer_io_enq_ready),
    .io_enq_valid(route_buffer_io_enq_valid),
    .io_enq_bits_head(route_buffer_io_enq_bits_head),
    .io_enq_bits_tail(route_buffer_io_enq_bits_tail),
    .io_enq_bits_payload(route_buffer_io_enq_bits_payload),
    .io_enq_bits_flow_ingress_node(route_buffer_io_enq_bits_flow_ingress_node),
    .io_enq_bits_flow_egress_node(route_buffer_io_enq_bits_flow_egress_node),
    .io_deq_ready(route_buffer_io_deq_ready),
    .io_deq_valid(route_buffer_io_deq_valid),
    .io_deq_bits_head(route_buffer_io_deq_bits_head),
    .io_deq_bits_tail(route_buffer_io_deq_bits_tail),
    .io_deq_bits_payload(route_buffer_io_deq_bits_payload),
    .io_deq_bits_flow_ingress_node(route_buffer_io_deq_bits_flow_ingress_node),
    .io_deq_bits_flow_egress_node(route_buffer_io_deq_bits_flow_egress_node)
  );
  Queue_9 route_q ( // @[IngressUnit.scala 27:23]
    .clock(route_q_clock),
    .reset(route_q_reset),
    .io_enq_ready(route_q_io_enq_ready),
    .io_enq_valid(route_q_io_enq_valid),
    .io_enq_bits_vc_sel_2_0(route_q_io_enq_bits_vc_sel_2_0),
    .io_enq_bits_vc_sel_1_0(route_q_io_enq_bits_vc_sel_1_0),
    .io_enq_bits_vc_sel_1_1(route_q_io_enq_bits_vc_sel_1_1),
    .io_enq_bits_vc_sel_1_2(route_q_io_enq_bits_vc_sel_1_2),
    .io_enq_bits_vc_sel_1_3(route_q_io_enq_bits_vc_sel_1_3),
    .io_enq_bits_vc_sel_0_0(route_q_io_enq_bits_vc_sel_0_0),
    .io_enq_bits_vc_sel_0_1(route_q_io_enq_bits_vc_sel_0_1),
    .io_enq_bits_vc_sel_0_2(route_q_io_enq_bits_vc_sel_0_2),
    .io_enq_bits_vc_sel_0_3(route_q_io_enq_bits_vc_sel_0_3),
    .io_deq_ready(route_q_io_deq_ready),
    .io_deq_valid(route_q_io_deq_valid),
    .io_deq_bits_vc_sel_2_0(route_q_io_deq_bits_vc_sel_2_0),
    .io_deq_bits_vc_sel_1_0(route_q_io_deq_bits_vc_sel_1_0),
    .io_deq_bits_vc_sel_1_1(route_q_io_deq_bits_vc_sel_1_1),
    .io_deq_bits_vc_sel_1_2(route_q_io_deq_bits_vc_sel_1_2),
    .io_deq_bits_vc_sel_1_3(route_q_io_deq_bits_vc_sel_1_3),
    .io_deq_bits_vc_sel_0_0(route_q_io_deq_bits_vc_sel_0_0),
    .io_deq_bits_vc_sel_0_1(route_q_io_deq_bits_vc_sel_0_1),
    .io_deq_bits_vc_sel_0_2(route_q_io_deq_bits_vc_sel_0_2),
    .io_deq_bits_vc_sel_0_3(route_q_io_deq_bits_vc_sel_0_3)
  );
  Queue_8 vcalloc_buffer ( // @[IngressUnit.scala 75:30]
    .clock(vcalloc_buffer_clock),
    .reset(vcalloc_buffer_reset),
    .io_enq_ready(vcalloc_buffer_io_enq_ready),
    .io_enq_valid(vcalloc_buffer_io_enq_valid),
    .io_enq_bits_head(vcalloc_buffer_io_enq_bits_head),
    .io_enq_bits_tail(vcalloc_buffer_io_enq_bits_tail),
    .io_enq_bits_payload(vcalloc_buffer_io_enq_bits_payload),
    .io_enq_bits_flow_ingress_node(vcalloc_buffer_io_enq_bits_flow_ingress_node),
    .io_enq_bits_flow_egress_node(vcalloc_buffer_io_enq_bits_flow_egress_node),
    .io_deq_ready(vcalloc_buffer_io_deq_ready),
    .io_deq_valid(vcalloc_buffer_io_deq_valid),
    .io_deq_bits_head(vcalloc_buffer_io_deq_bits_head),
    .io_deq_bits_tail(vcalloc_buffer_io_deq_bits_tail),
    .io_deq_bits_payload(vcalloc_buffer_io_deq_bits_payload),
    .io_deq_bits_flow_ingress_node(vcalloc_buffer_io_deq_bits_flow_ingress_node),
    .io_deq_bits_flow_egress_node(vcalloc_buffer_io_deq_bits_flow_egress_node)
  );
  Queue_11 vcalloc_q ( // @[IngressUnit.scala 76:25]
    .clock(vcalloc_q_clock),
    .reset(vcalloc_q_reset),
    .io_enq_ready(vcalloc_q_io_enq_ready),
    .io_enq_valid(vcalloc_q_io_enq_valid),
    .io_enq_bits_vc_sel_2_0(vcalloc_q_io_enq_bits_vc_sel_2_0),
    .io_enq_bits_vc_sel_1_0(vcalloc_q_io_enq_bits_vc_sel_1_0),
    .io_enq_bits_vc_sel_1_1(vcalloc_q_io_enq_bits_vc_sel_1_1),
    .io_enq_bits_vc_sel_1_2(vcalloc_q_io_enq_bits_vc_sel_1_2),
    .io_enq_bits_vc_sel_1_3(vcalloc_q_io_enq_bits_vc_sel_1_3),
    .io_enq_bits_vc_sel_0_0(vcalloc_q_io_enq_bits_vc_sel_0_0),
    .io_enq_bits_vc_sel_0_1(vcalloc_q_io_enq_bits_vc_sel_0_1),
    .io_enq_bits_vc_sel_0_2(vcalloc_q_io_enq_bits_vc_sel_0_2),
    .io_enq_bits_vc_sel_0_3(vcalloc_q_io_enq_bits_vc_sel_0_3),
    .io_deq_ready(vcalloc_q_io_deq_ready),
    .io_deq_valid(vcalloc_q_io_deq_valid),
    .io_deq_bits_vc_sel_2_0(vcalloc_q_io_deq_bits_vc_sel_2_0),
    .io_deq_bits_vc_sel_1_0(vcalloc_q_io_deq_bits_vc_sel_1_0),
    .io_deq_bits_vc_sel_1_1(vcalloc_q_io_deq_bits_vc_sel_1_1),
    .io_deq_bits_vc_sel_1_2(vcalloc_q_io_deq_bits_vc_sel_1_2),
    .io_deq_bits_vc_sel_1_3(vcalloc_q_io_deq_bits_vc_sel_1_3),
    .io_deq_bits_vc_sel_0_0(vcalloc_q_io_deq_bits_vc_sel_0_0),
    .io_deq_bits_vc_sel_0_1(vcalloc_q_io_deq_bits_vc_sel_0_1),
    .io_deq_bits_vc_sel_0_2(vcalloc_q_io_deq_bits_vc_sel_0_2),
    .io_deq_bits_vc_sel_0_3(vcalloc_q_io_deq_bits_vc_sel_0_3)
  );
  assign io_router_req_valid = io_in_valid & route_buffer_io_enq_ready & io_in_bits_head & ~at_dest; // @[IngressUnit.scala 58:86]
  assign io_router_req_bits_flow_ingress_node = route_buffer_io_enq_bits_flow_ingress_node; // @[IngressUnit.scala 53:27]
  assign io_router_req_bits_flow_egress_node = route_buffer_io_enq_bits_flow_egress_node; // @[IngressUnit.scala 53:27]
  assign io_vcalloc_req_valid = _io_vcalloc_req_valid_T_1 & vcalloc_buffer_io_enq_ready & vcalloc_q_io_enq_ready; // @[IngressUnit.scala 92:41]
  assign io_vcalloc_req_bits_vc_sel_2_0 = route_q_io_deq_bits_vc_sel_2_0; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_1_0 = route_q_io_deq_bits_vc_sel_1_0; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_1_1 = route_q_io_deq_bits_vc_sel_1_1; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_1_2 = route_q_io_deq_bits_vc_sel_1_2; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_1_3 = route_q_io_deq_bits_vc_sel_1_3; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_0_0 = route_q_io_deq_bits_vc_sel_0_0; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_0_1 = route_q_io_deq_bits_vc_sel_0_1; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_0_2 = route_q_io_deq_bits_vc_sel_0_2; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_0_3 = route_q_io_deq_bits_vc_sel_0_3; // @[IngressUnit.scala 81:30]
  assign io_salloc_req_0_valid = vcalloc_buffer_io_deq_valid & vcalloc_q_io_deq_valid & c; // @[IngressUnit.scala 109:83]
  assign io_salloc_req_0_bits_vc_sel_2_0 = vcalloc_q_io_deq_bits_vc_sel_2_0; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_1_0 = vcalloc_q_io_deq_bits_vc_sel_1_0; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_1_1 = vcalloc_q_io_deq_bits_vc_sel_1_1; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_1_2 = vcalloc_q_io_deq_bits_vc_sel_1_2; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_1_3 = vcalloc_q_io_deq_bits_vc_sel_1_3; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_0_0 = vcalloc_q_io_deq_bits_vc_sel_0_0; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_0_1 = vcalloc_q_io_deq_bits_vc_sel_0_1; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_0_2 = vcalloc_q_io_deq_bits_vc_sel_0_2; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_0_3 = vcalloc_q_io_deq_bits_vc_sel_0_3; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_tail = vcalloc_buffer_io_deq_bits_tail; // @[IngressUnit.scala 105:30]
  assign io_out_0_valid = out_bundle_valid; // @[IngressUnit.scala 118:13]
  assign io_out_0_bits_flit_head = out_bundle_bits_flit_head; // @[IngressUnit.scala 118:13]
  assign io_out_0_bits_flit_tail = out_bundle_bits_flit_tail; // @[IngressUnit.scala 118:13]
  assign io_out_0_bits_flit_payload = out_bundle_bits_flit_payload; // @[IngressUnit.scala 118:13]
  assign io_out_0_bits_flit_flow_ingress_node = out_bundle_bits_flit_flow_ingress_node; // @[IngressUnit.scala 118:13]
  assign io_out_0_bits_flit_flow_egress_node = out_bundle_bits_flit_flow_egress_node; // @[IngressUnit.scala 118:13]
  assign io_out_0_bits_out_virt_channel = out_bundle_bits_out_virt_channel; // @[IngressUnit.scala 118:13]
  assign io_in_ready = route_buffer_io_enq_ready; // @[IngressUnit.scala 59:44]
  assign route_buffer_clock = clock;
  assign route_buffer_reset = reset;
  assign route_buffer_io_enq_valid = io_in_valid; // @[IngressUnit.scala 56:44]
  assign route_buffer_io_enq_bits_head = io_in_bits_head; // @[IngressUnit.scala 32:33]
  assign route_buffer_io_enq_bits_tail = io_in_bits_tail; // @[IngressUnit.scala 33:33]
  assign route_buffer_io_enq_bits_payload = io_in_bits_payload; // @[IngressUnit.scala 50:36]
  assign route_buffer_io_enq_bits_flow_ingress_node = 2'h3; // @[IngressUnit.scala 38:51]
  assign route_buffer_io_enq_bits_flow_egress_node = _route_buffer_io_enq_bits_flow_egress_node_T_9 |
    _route_buffer_io_enq_bits_flow_egress_node_T_7; // @[Mux.scala 27:73]
  assign route_buffer_io_deq_ready = _route_buffer_io_deq_ready_T_5 & _route_buffer_io_deq_ready_T_7; // @[IngressUnit.scala 95:37]
  assign route_q_clock = clock;
  assign route_q_reset = reset;
  assign route_q_io_enq_valid = _T_13 & io_in_bits_head & at_dest | io_router_req_valid; // @[IngressUnit.scala 62:24 64:53 65:26]
  assign route_q_io_enq_bits_vc_sel_2_0 = _T_13 & io_in_bits_head & at_dest & _T_3; // @[IngressUnit.scala 63:23 64:53]
  assign route_q_io_enq_bits_vc_sel_1_0 = _T_13 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_1_0; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_1_1 = _T_13 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_1_1; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_1_2 = _T_13 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_1_2; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_1_3 = _T_13 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_1_3; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_0_0 = _T_13 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_0_0; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_0_1 = _T_13 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_0_1; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_0_2 = _T_13 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_0_2; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_0_3 = _T_13 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_0_3; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_deq_ready = _route_q_io_deq_ready_T & route_buffer_io_deq_bits_tail; // @[IngressUnit.scala 97:55]
  assign vcalloc_buffer_clock = clock;
  assign vcalloc_buffer_reset = reset;
  assign vcalloc_buffer_io_enq_valid = _vcalloc_buffer_io_enq_valid_T_2 & _vcalloc_buffer_io_enq_valid_T_4; // @[IngressUnit.scala 88:37]
  assign vcalloc_buffer_io_enq_bits_head = route_buffer_io_deq_bits_head; // @[IngressUnit.scala 79:30]
  assign vcalloc_buffer_io_enq_bits_tail = route_buffer_io_deq_bits_tail; // @[IngressUnit.scala 79:30]
  assign vcalloc_buffer_io_enq_bits_payload = route_buffer_io_deq_bits_payload; // @[IngressUnit.scala 79:30]
  assign vcalloc_buffer_io_enq_bits_flow_ingress_node = route_buffer_io_deq_bits_flow_ingress_node; // @[IngressUnit.scala 79:30]
  assign vcalloc_buffer_io_enq_bits_flow_egress_node = route_buffer_io_deq_bits_flow_egress_node; // @[IngressUnit.scala 79:30]
  assign vcalloc_buffer_io_deq_ready = io_salloc_req_0_ready & vcalloc_q_io_deq_valid & c; // @[IngressUnit.scala 110:83]
  assign vcalloc_q_clock = clock;
  assign vcalloc_q_reset = reset;
  assign vcalloc_q_io_enq_valid = io_vcalloc_req_ready & io_vcalloc_req_valid; // @[Decoupled.scala 51:35]
  assign vcalloc_q_io_enq_bits_vc_sel_2_0 = io_vcalloc_resp_vc_sel_2_0; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_1_0 = io_vcalloc_resp_vc_sel_1_0; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_1_1 = io_vcalloc_resp_vc_sel_1_1; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_1_2 = io_vcalloc_resp_vc_sel_1_2; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_1_3 = io_vcalloc_resp_vc_sel_1_3; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_0_0 = io_vcalloc_resp_vc_sel_0_0; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_0_1 = io_vcalloc_resp_vc_sel_0_1; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_0_2 = io_vcalloc_resp_vc_sel_0_2; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_0_3 = io_vcalloc_resp_vc_sel_0_3; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_deq_ready = vcalloc_buffer_io_deq_bits_tail & _vcalloc_q_io_deq_ready_T; // @[IngressUnit.scala 111:42]
  always @(posedge clock) begin
    out_bundle_valid <= vcalloc_buffer_io_deq_ready & vcalloc_buffer_io_deq_valid; // @[Decoupled.scala 51:35]
    out_bundle_bits_flit_head <= vcalloc_buffer_io_deq_bits_head; // @[IngressUnit.scala 121:24]
    out_bundle_bits_flit_tail <= vcalloc_buffer_io_deq_bits_tail; // @[IngressUnit.scala 121:24]
    out_bundle_bits_flit_payload <= vcalloc_buffer_io_deq_bits_payload; // @[IngressUnit.scala 121:24]
    out_bundle_bits_flit_flow_ingress_node <= vcalloc_buffer_io_deq_bits_flow_ingress_node; // @[IngressUnit.scala 121:24]
    out_bundle_bits_flit_flow_egress_node <= vcalloc_buffer_io_deq_bits_flow_egress_node; // @[IngressUnit.scala 121:24]
    out_bundle_bits_out_virt_channel <= _out_bundle_bits_out_virt_channel_T_10 | _out_bundle_bits_out_virt_channel_T_11; // @[Mux.scala 27:73]
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~(io_in_valid & ~_T_6))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at IngressUnit.scala:30 assert(!(io.in.valid && !cParam.possibleFlows.toSeq.map(_.egressId.U === io.in.bits.egress_id).orR))\n"
            ); // @[IngressUnit.scala 30:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_11 & ~(~(route_q_io_enq_valid & ~route_q_io_enq_ready))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at IngressUnit.scala:73 assert(!(route_q.io.enq.valid && !route_q.io.enq.ready))\n"); // @[IngressUnit.scala 73:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_11 & ~(~(vcalloc_q_io_enq_valid & ~vcalloc_q_io_enq_ready))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at IngressUnit.scala:102 assert(!(vcalloc_q.io.enq.valid && !vcalloc_q.io.enq.ready))\n"
            ); // @[IngressUnit.scala 102:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  out_bundle_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  out_bundle_bits_flit_head = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  out_bundle_bits_flit_tail = _RAND_2[0:0];
  _RAND_3 = {2{`RANDOM}};
  out_bundle_bits_flit_payload = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  out_bundle_bits_flit_flow_ingress_node = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  out_bundle_bits_flit_flow_egress_node = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  out_bundle_bits_out_virt_channel = _RAND_6[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(~(io_in_valid & ~_T_6)); // @[IngressUnit.scala 30:9]
    end
    //
    if (_T_11) begin
      assert(~(route_q_io_enq_valid & ~route_q_io_enq_ready)); // @[IngressUnit.scala 73:9]
    end
    //
    if (_T_11) begin
      assert(~(vcalloc_q_io_enq_valid & ~vcalloc_q_io_enq_ready)); // @[IngressUnit.scala 102:9]
    end
  end
endmodule
module RouteComputer_3(
  input  [1:0] io_req_2_bits_flow_ingress_node,
  input  [1:0] io_req_2_bits_flow_egress_node,
  input  [1:0] io_req_1_bits_src_virt_id,
  input  [1:0] io_req_1_bits_flow_ingress_node,
  input  [1:0] io_req_1_bits_flow_egress_node,
  input  [1:0] io_req_0_bits_src_virt_id,
  input  [1:0] io_req_0_bits_flow_ingress_node,
  input  [1:0] io_req_0_bits_flow_egress_node,
  output       io_resp_2_vc_sel_1_0,
  output       io_resp_2_vc_sel_1_1,
  output       io_resp_2_vc_sel_1_2,
  output       io_resp_2_vc_sel_1_3,
  output       io_resp_2_vc_sel_0_0,
  output       io_resp_2_vc_sel_0_1,
  output       io_resp_2_vc_sel_0_2,
  output       io_resp_2_vc_sel_0_3,
  output       io_resp_1_vc_sel_1_0,
  output       io_resp_1_vc_sel_1_1,
  output       io_resp_1_vc_sel_1_2,
  output       io_resp_1_vc_sel_1_3,
  output       io_resp_1_vc_sel_0_0,
  output       io_resp_1_vc_sel_0_1,
  output       io_resp_1_vc_sel_0_2,
  output       io_resp_0_vc_sel_1_0,
  output       io_resp_0_vc_sel_1_1,
  output       io_resp_0_vc_sel_1_2,
  output       io_resp_0_vc_sel_1_3,
  output       io_resp_0_vc_sel_0_0,
  output       io_resp_0_vc_sel_0_1,
  output       io_resp_0_vc_sel_0_2
);
  wire [5:0] addr = {io_req_0_bits_src_virt_id,io_req_0_bits_flow_ingress_node,io_req_0_bits_flow_egress_node}; // @[RouteComputer.scala 74:27]
  wire [5:0] decoded_invInputs = ~addr; // @[pla.scala 78:21]
  wire  decoded_andMatrixInput_0 = decoded_invInputs[4]; // @[pla.scala 91:29]
  wire  decoded_andMatrixInput_1 = decoded_invInputs[5]; // @[pla.scala 91:29]
  wire [1:0] _decoded_T = {decoded_andMatrixInput_0,decoded_andMatrixInput_1}; // @[Cat.scala 33:92]
  wire  _decoded_T_1 = &_decoded_T; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_0_1 = decoded_invInputs[0]; // @[pla.scala 91:29]
  wire  decoded_andMatrixInput_1_1 = addr[1]; // @[pla.scala 90:45]
  wire [1:0] _decoded_T_2 = {decoded_andMatrixInput_0_1,decoded_andMatrixInput_1_1}; // @[Cat.scala 33:92]
  wire  _decoded_T_3 = &_decoded_T_2; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_0_2 = addr[0]; // @[pla.scala 90:45]
  wire [1:0] _decoded_T_4 = {decoded_andMatrixInput_0_2,decoded_andMatrixInput_1_1}; // @[Cat.scala 33:92]
  wire  _decoded_T_5 = &_decoded_T_4; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_1_3 = addr[4]; // @[pla.scala 90:45]
  wire [1:0] _decoded_T_6 = {decoded_andMatrixInput_1_1,decoded_andMatrixInput_1_3}; // @[Cat.scala 33:92]
  wire  _decoded_T_7 = &_decoded_T_6; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_1_4 = addr[5]; // @[pla.scala 90:45]
  wire [1:0] _decoded_T_8 = {decoded_andMatrixInput_1_1,decoded_andMatrixInput_1_4}; // @[Cat.scala 33:92]
  wire  _decoded_T_9 = &_decoded_T_8; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_2 = decoded_invInputs[3]; // @[pla.scala 91:29]
  wire [3:0] _decoded_T_10 = {decoded_andMatrixInput_0_2,decoded_andMatrixInput_1_1,decoded_andMatrixInput_2,
    decoded_andMatrixInput_1_4}; // @[Cat.scala 33:92]
  wire  _decoded_T_11 = &_decoded_T_10; // @[pla.scala 98:74]
  wire [1:0] _decoded_T_12 = {decoded_andMatrixInput_1_3,decoded_andMatrixInput_1_4}; // @[Cat.scala 33:92]
  wire  _decoded_T_13 = &_decoded_T_12; // @[pla.scala 98:74]
  wire [3:0] _decoded_T_14 = {decoded_andMatrixInput_0_2,decoded_andMatrixInput_2,decoded_andMatrixInput_1_3,
    decoded_andMatrixInput_1_4}; // @[Cat.scala 33:92]
  wire  _decoded_T_15 = &_decoded_T_14; // @[pla.scala 98:74]
  wire  _decoded_orMatrixOutputs_T = |_decoded_T_13; // @[pla.scala 114:39]
  wire  _decoded_orMatrixOutputs_T_1 = |_decoded_T_9; // @[pla.scala 114:39]
  wire [1:0] _decoded_orMatrixOutputs_T_2 = {_decoded_T_7,_decoded_T_9}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_3 = |_decoded_orMatrixOutputs_T_2; // @[pla.scala 114:39]
  wire [1:0] _decoded_orMatrixOutputs_T_4 = {_decoded_T_1,_decoded_T_3}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_5 = |_decoded_orMatrixOutputs_T_4; // @[pla.scala 114:39]
  wire  _decoded_orMatrixOutputs_T_6 = |_decoded_T_15; // @[pla.scala 114:39]
  wire  _decoded_orMatrixOutputs_T_7 = |_decoded_T_11; // @[pla.scala 114:39]
  wire  _decoded_orMatrixOutputs_T_8 = |_decoded_T_5; // @[pla.scala 114:39]
  wire [7:0] decoded_orMatrixOutputs = {_decoded_orMatrixOutputs_T_8,_decoded_orMatrixOutputs_T_7,
    _decoded_orMatrixOutputs_T_6,1'h0,_decoded_orMatrixOutputs_T_5,_decoded_orMatrixOutputs_T_3,
    _decoded_orMatrixOutputs_T_1,_decoded_orMatrixOutputs_T}; // @[Cat.scala 33:92]
  wire [7:0] decoded_invMatrixOutputs = {decoded_orMatrixOutputs[7],decoded_orMatrixOutputs[6],decoded_orMatrixOutputs[5
    ],decoded_orMatrixOutputs[4],decoded_orMatrixOutputs[3],decoded_orMatrixOutputs[2],decoded_orMatrixOutputs[1],
    decoded_orMatrixOutputs[0]}; // @[Cat.scala 33:92]
  wire [7:0] _GEN_0 = {{4'd0}, decoded_invMatrixOutputs[7:4]}; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_19 = _GEN_0 & 8'hf; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_21 = {decoded_invMatrixOutputs[3:0], 4'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _decoded_T_23 = _decoded_T_21 & 8'hf0; // @[Bitwise.scala 108:80]
  wire [7:0] _decoded_T_24 = _decoded_T_19 | _decoded_T_23; // @[Bitwise.scala 108:39]
  wire [7:0] _GEN_1 = {{2'd0}, _decoded_T_24[7:2]}; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_29 = _GEN_1 & 8'h33; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_31 = {_decoded_T_24[5:0], 2'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _decoded_T_33 = _decoded_T_31 & 8'hcc; // @[Bitwise.scala 108:80]
  wire [7:0] _decoded_T_34 = _decoded_T_29 | _decoded_T_33; // @[Bitwise.scala 108:39]
  wire [7:0] _GEN_2 = {{1'd0}, _decoded_T_34[7:1]}; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_39 = _GEN_2 & 8'h55; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_41 = {_decoded_T_34[6:0], 1'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _decoded_T_43 = _decoded_T_41 & 8'haa; // @[Bitwise.scala 108:80]
  wire [7:0] decoded = _decoded_T_39 | _decoded_T_43; // @[Bitwise.scala 108:39]
  wire [5:0] addr_1 = {io_req_1_bits_src_virt_id,io_req_1_bits_flow_ingress_node,io_req_1_bits_flow_egress_node}; // @[RouteComputer.scala 74:27]
  wire [5:0] decoded_invInputs_1 = ~addr_1; // @[pla.scala 78:21]
  wire  decoded_andMatrixInput_0_8 = decoded_invInputs_1[0]; // @[pla.scala 91:29]
  wire  decoded_andMatrixInput_1_8 = decoded_invInputs_1[1]; // @[pla.scala 91:29]
  wire [1:0] _decoded_T_44 = {decoded_andMatrixInput_0_8,decoded_andMatrixInput_1_8}; // @[Cat.scala 33:92]
  wire  _decoded_T_45 = &_decoded_T_44; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_0_9 = decoded_invInputs_1[3]; // @[pla.scala 91:29]
  wire  decoded_andMatrixInput_1_9 = decoded_invInputs_1[4]; // @[pla.scala 91:29]
  wire  decoded_andMatrixInput_2_2 = decoded_invInputs_1[5]; // @[pla.scala 91:29]
  wire [2:0] _decoded_T_46 = {decoded_andMatrixInput_0_9,decoded_andMatrixInput_1_9,decoded_andMatrixInput_2_2}; // @[Cat.scala 33:92]
  wire  _decoded_T_47 = &_decoded_T_46; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_0_10 = addr_1[0]; // @[pla.scala 90:45]
  wire  decoded_andMatrixInput_1_10 = addr_1[1]; // @[pla.scala 90:45]
  wire [1:0] _decoded_T_48 = {decoded_andMatrixInput_0_10,decoded_andMatrixInput_1_10}; // @[Cat.scala 33:92]
  wire  _decoded_T_49 = &_decoded_T_48; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_1_11 = decoded_invInputs_1[2]; // @[pla.scala 91:29]
  wire  decoded_andMatrixInput_2_3 = addr_1[3]; // @[pla.scala 90:45]
  wire [4:0] _decoded_T_50 = {decoded_andMatrixInput_1_10,decoded_andMatrixInput_1_11,decoded_andMatrixInput_2_3,
    decoded_andMatrixInput_1_9,decoded_andMatrixInput_2_2}; // @[Cat.scala 33:92]
  wire  _decoded_T_51 = &_decoded_T_50; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_1_12 = addr_1[4]; // @[pla.scala 90:45]
  wire [1:0] _decoded_T_52 = {decoded_andMatrixInput_0_10,decoded_andMatrixInput_1_12}; // @[Cat.scala 33:92]
  wire  _decoded_T_53 = &_decoded_T_52; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_1_13 = addr_1[5]; // @[pla.scala 90:45]
  wire [1:0] _decoded_T_54 = {decoded_andMatrixInput_1_11,decoded_andMatrixInput_1_13}; // @[Cat.scala 33:92]
  wire  _decoded_T_55 = &_decoded_T_54; // @[pla.scala 98:74]
  wire [1:0] _decoded_T_56 = {decoded_andMatrixInput_0_10,decoded_andMatrixInput_1_13}; // @[Cat.scala 33:92]
  wire  _decoded_T_57 = &_decoded_T_56; // @[pla.scala 98:74]
  wire [1:0] _decoded_T_58 = {decoded_andMatrixInput_1_12,decoded_andMatrixInput_1_13}; // @[Cat.scala 33:92]
  wire  _decoded_T_59 = &_decoded_T_58; // @[pla.scala 98:74]
  wire [2:0] _decoded_T_60 = {decoded_andMatrixInput_0_9,decoded_andMatrixInput_1_12,decoded_andMatrixInput_1_13}; // @[Cat.scala 33:92]
  wire  _decoded_T_61 = &_decoded_T_60; // @[pla.scala 98:74]
  wire [4:0] _decoded_T_62 = {decoded_andMatrixInput_1_10,decoded_andMatrixInput_1_11,decoded_andMatrixInput_2_3,
    decoded_andMatrixInput_1_12,decoded_andMatrixInput_1_13}; // @[Cat.scala 33:92]
  wire  _decoded_T_63 = &_decoded_T_62; // @[pla.scala 98:74]
  wire [1:0] _decoded_orMatrixOutputs_T_9 = {_decoded_T_61,_decoded_T_63}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_10 = |_decoded_orMatrixOutputs_T_9; // @[pla.scala 114:39]
  wire  _decoded_orMatrixOutputs_T_11 = |_decoded_T_57; // @[pla.scala 114:39]
  wire [1:0] _decoded_orMatrixOutputs_T_12 = {_decoded_T_53,_decoded_T_57}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_13 = |_decoded_orMatrixOutputs_T_12; // @[pla.scala 114:39]
  wire [1:0] _decoded_orMatrixOutputs_T_14 = {_decoded_T_47,_decoded_T_51}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_15 = |_decoded_orMatrixOutputs_T_14; // @[pla.scala 114:39]
  wire  _decoded_orMatrixOutputs_T_16 = |_decoded_T_59; // @[pla.scala 114:39]
  wire [1:0] _decoded_orMatrixOutputs_T_17 = {_decoded_T_55,_decoded_T_57}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_18 = |_decoded_orMatrixOutputs_T_17; // @[pla.scala 114:39]
  wire [1:0] _decoded_orMatrixOutputs_T_19 = {_decoded_T_45,_decoded_T_49}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_20 = |_decoded_orMatrixOutputs_T_19; // @[pla.scala 114:39]
  wire [7:0] decoded_orMatrixOutputs_1 = {_decoded_orMatrixOutputs_T_20,_decoded_orMatrixOutputs_T_18,
    _decoded_orMatrixOutputs_T_16,1'h0,_decoded_orMatrixOutputs_T_15,_decoded_orMatrixOutputs_T_13,
    _decoded_orMatrixOutputs_T_11,_decoded_orMatrixOutputs_T_10}; // @[Cat.scala 33:92]
  wire [7:0] decoded_invMatrixOutputs_1 = {decoded_orMatrixOutputs_1[7],decoded_orMatrixOutputs_1[6],
    decoded_orMatrixOutputs_1[5],decoded_orMatrixOutputs_1[4],decoded_orMatrixOutputs_1[3],decoded_orMatrixOutputs_1[2],
    decoded_orMatrixOutputs_1[1],decoded_orMatrixOutputs_1[0]}; // @[Cat.scala 33:92]
  wire [7:0] _GEN_3 = {{4'd0}, decoded_invMatrixOutputs_1[7:4]}; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_67 = _GEN_3 & 8'hf; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_69 = {decoded_invMatrixOutputs_1[3:0], 4'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _decoded_T_71 = _decoded_T_69 & 8'hf0; // @[Bitwise.scala 108:80]
  wire [7:0] _decoded_T_72 = _decoded_T_67 | _decoded_T_71; // @[Bitwise.scala 108:39]
  wire [7:0] _GEN_4 = {{2'd0}, _decoded_T_72[7:2]}; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_77 = _GEN_4 & 8'h33; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_79 = {_decoded_T_72[5:0], 2'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _decoded_T_81 = _decoded_T_79 & 8'hcc; // @[Bitwise.scala 108:80]
  wire [7:0] _decoded_T_82 = _decoded_T_77 | _decoded_T_81; // @[Bitwise.scala 108:39]
  wire [7:0] _GEN_5 = {{1'd0}, _decoded_T_82[7:1]}; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_87 = _GEN_5 & 8'h55; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_89 = {_decoded_T_82[6:0], 1'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _decoded_T_91 = _decoded_T_89 & 8'haa; // @[Bitwise.scala 108:80]
  wire [7:0] decoded_1 = _decoded_T_87 | _decoded_T_91; // @[Bitwise.scala 108:39]
  wire [5:0] addr_2 = {2'h0,io_req_2_bits_flow_ingress_node,io_req_2_bits_flow_egress_node}; // @[RouteComputer.scala 74:27]
  wire [5:0] decoded_invInputs_2 = ~addr_2; // @[pla.scala 78:21]
  wire  decoded_andMatrixInput_0_18 = decoded_invInputs_2[1]; // @[pla.scala 91:29]
  wire  decoded_andMatrixInput_1_18 = addr_2[2]; // @[pla.scala 90:45]
  wire  decoded_andMatrixInput_2_6 = addr_2[3]; // @[pla.scala 90:45]
  wire  decoded_andMatrixInput_3_4 = decoded_invInputs_2[4]; // @[pla.scala 91:29]
  wire  decoded_andMatrixInput_4_2 = decoded_invInputs_2[5]; // @[pla.scala 91:29]
  wire [4:0] _decoded_T_92 = {decoded_andMatrixInput_0_18,decoded_andMatrixInput_1_18,decoded_andMatrixInput_2_6,
    decoded_andMatrixInput_3_4,decoded_andMatrixInput_4_2}; // @[Cat.scala 33:92]
  wire  _decoded_T_93 = &_decoded_T_92; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_0_19 = addr_2[0]; // @[pla.scala 90:45]
  wire [4:0] _decoded_T_94 = {decoded_andMatrixInput_0_19,decoded_andMatrixInput_1_18,decoded_andMatrixInput_2_6,
    decoded_andMatrixInput_3_4,decoded_andMatrixInput_4_2}; // @[Cat.scala 33:92]
  wire  _decoded_T_95 = &_decoded_T_94; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_0_20 = addr_2[1]; // @[pla.scala 90:45]
  wire [4:0] _decoded_T_96 = {decoded_andMatrixInput_0_20,decoded_andMatrixInput_1_18,decoded_andMatrixInput_2_6,
    decoded_andMatrixInput_3_4,decoded_andMatrixInput_4_2}; // @[Cat.scala 33:92]
  wire  _decoded_T_97 = &_decoded_T_96; // @[pla.scala 98:74]
  wire [1:0] _decoded_orMatrixOutputs_T_21 = {_decoded_T_95,_decoded_T_97}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_22 = |_decoded_orMatrixOutputs_T_21; // @[pla.scala 114:39]
  wire [1:0] _decoded_orMatrixOutputs_T_27 = {_decoded_T_93,_decoded_T_95}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_28 = |_decoded_orMatrixOutputs_T_27; // @[pla.scala 114:39]
  wire [7:0] decoded_orMatrixOutputs_2 = {1'h0,_decoded_orMatrixOutputs_T_28,_decoded_orMatrixOutputs_T_28,
    _decoded_orMatrixOutputs_T_28,1'h0,_decoded_orMatrixOutputs_T_22,_decoded_orMatrixOutputs_T_22,
    _decoded_orMatrixOutputs_T_22}; // @[Cat.scala 33:92]
  wire [7:0] decoded_invMatrixOutputs_2 = {decoded_orMatrixOutputs_2[7],decoded_orMatrixOutputs_2[6],
    decoded_orMatrixOutputs_2[5],decoded_orMatrixOutputs_2[4],decoded_orMatrixOutputs_2[3],decoded_orMatrixOutputs_2[2],
    decoded_orMatrixOutputs_2[1],decoded_orMatrixOutputs_2[0]}; // @[Cat.scala 33:92]
  wire [7:0] _GEN_6 = {{4'd0}, decoded_invMatrixOutputs_2[7:4]}; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_101 = _GEN_6 & 8'hf; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_103 = {decoded_invMatrixOutputs_2[3:0], 4'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _decoded_T_105 = _decoded_T_103 & 8'hf0; // @[Bitwise.scala 108:80]
  wire [7:0] _decoded_T_106 = _decoded_T_101 | _decoded_T_105; // @[Bitwise.scala 108:39]
  wire [7:0] _GEN_7 = {{2'd0}, _decoded_T_106[7:2]}; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_111 = _GEN_7 & 8'h33; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_113 = {_decoded_T_106[5:0], 2'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _decoded_T_115 = _decoded_T_113 & 8'hcc; // @[Bitwise.scala 108:80]
  wire [7:0] _decoded_T_116 = _decoded_T_111 | _decoded_T_115; // @[Bitwise.scala 108:39]
  wire [7:0] _GEN_8 = {{1'd0}, _decoded_T_116[7:1]}; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_121 = _GEN_8 & 8'h55; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_123 = {_decoded_T_116[6:0], 1'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _decoded_T_125 = _decoded_T_123 & 8'haa; // @[Bitwise.scala 108:80]
  wire [7:0] decoded_2 = _decoded_T_121 | _decoded_T_125; // @[Bitwise.scala 108:39]
  assign io_resp_2_vc_sel_1_0 = decoded_2[4]; // @[RouteComputer.scala 90:46]
  assign io_resp_2_vc_sel_1_1 = decoded_2[5]; // @[RouteComputer.scala 90:46]
  assign io_resp_2_vc_sel_1_2 = decoded_2[6]; // @[RouteComputer.scala 90:46]
  assign io_resp_2_vc_sel_1_3 = decoded_2[7]; // @[RouteComputer.scala 90:46]
  assign io_resp_2_vc_sel_0_0 = decoded_2[0]; // @[RouteComputer.scala 90:46]
  assign io_resp_2_vc_sel_0_1 = decoded_2[1]; // @[RouteComputer.scala 90:46]
  assign io_resp_2_vc_sel_0_2 = decoded_2[2]; // @[RouteComputer.scala 90:46]
  assign io_resp_2_vc_sel_0_3 = decoded_2[3]; // @[RouteComputer.scala 90:46]
  assign io_resp_1_vc_sel_1_0 = decoded_1[4]; // @[RouteComputer.scala 90:46]
  assign io_resp_1_vc_sel_1_1 = decoded_1[5]; // @[RouteComputer.scala 90:46]
  assign io_resp_1_vc_sel_1_2 = decoded_1[6]; // @[RouteComputer.scala 90:46]
  assign io_resp_1_vc_sel_1_3 = decoded_1[7]; // @[RouteComputer.scala 90:46]
  assign io_resp_1_vc_sel_0_0 = decoded_1[0]; // @[RouteComputer.scala 90:46]
  assign io_resp_1_vc_sel_0_1 = decoded_1[1]; // @[RouteComputer.scala 90:46]
  assign io_resp_1_vc_sel_0_2 = decoded_1[2]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_1_0 = decoded[4]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_1_1 = decoded[5]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_1_2 = decoded[6]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_1_3 = decoded[7]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_0_0 = decoded[0]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_0_1 = decoded[1]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_0_2 = decoded[2]; // @[RouteComputer.scala 90:46]
endmodule
module Router_3(
  input         clock,
  input         reset,
  output [1:0]  auto_debug_out_va_stall_0,
  output [1:0]  auto_debug_out_va_stall_1,
  output [1:0]  auto_debug_out_sa_stall_0,
  output [1:0]  auto_debug_out_sa_stall_1,
  output        auto_egress_nodes_out_flit_valid,
  output        auto_egress_nodes_out_flit_bits_head,
  output        auto_egress_nodes_out_flit_bits_tail,
  output [63:0] auto_egress_nodes_out_flit_bits_payload,
  output [1:0]  auto_egress_nodes_out_flit_bits_ingress_id,
  output        auto_ingress_nodes_in_flit_ready,
  input         auto_ingress_nodes_in_flit_valid,
  input         auto_ingress_nodes_in_flit_bits_head,
  input         auto_ingress_nodes_in_flit_bits_tail,
  input  [63:0] auto_ingress_nodes_in_flit_bits_payload,
  input  [1:0]  auto_ingress_nodes_in_flit_bits_egress_id,
  output        auto_source_nodes_out_1_flit_0_valid,
  output        auto_source_nodes_out_1_flit_0_bits_head,
  output        auto_source_nodes_out_1_flit_0_bits_tail,
  output [63:0] auto_source_nodes_out_1_flit_0_bits_payload,
  output [1:0]  auto_source_nodes_out_1_flit_0_bits_flow_ingress_node,
  output [1:0]  auto_source_nodes_out_1_flit_0_bits_flow_egress_node,
  output [1:0]  auto_source_nodes_out_1_flit_0_bits_virt_channel_id,
  input  [3:0]  auto_source_nodes_out_1_credit_return,
  input  [3:0]  auto_source_nodes_out_1_vc_free,
  output        auto_source_nodes_out_0_flit_0_valid,
  output        auto_source_nodes_out_0_flit_0_bits_head,
  output        auto_source_nodes_out_0_flit_0_bits_tail,
  output [63:0] auto_source_nodes_out_0_flit_0_bits_payload,
  output [1:0]  auto_source_nodes_out_0_flit_0_bits_flow_ingress_node,
  output [1:0]  auto_source_nodes_out_0_flit_0_bits_flow_egress_node,
  output [1:0]  auto_source_nodes_out_0_flit_0_bits_virt_channel_id,
  input  [3:0]  auto_source_nodes_out_0_credit_return,
  input  [3:0]  auto_source_nodes_out_0_vc_free,
  input         auto_dest_nodes_in_1_flit_0_valid,
  input         auto_dest_nodes_in_1_flit_0_bits_head,
  input         auto_dest_nodes_in_1_flit_0_bits_tail,
  input  [63:0] auto_dest_nodes_in_1_flit_0_bits_payload,
  input  [1:0]  auto_dest_nodes_in_1_flit_0_bits_flow_ingress_node,
  input  [1:0]  auto_dest_nodes_in_1_flit_0_bits_flow_egress_node,
  input  [1:0]  auto_dest_nodes_in_1_flit_0_bits_virt_channel_id,
  output [3:0]  auto_dest_nodes_in_1_credit_return,
  output [3:0]  auto_dest_nodes_in_1_vc_free,
  input         auto_dest_nodes_in_0_flit_0_valid,
  input         auto_dest_nodes_in_0_flit_0_bits_head,
  input         auto_dest_nodes_in_0_flit_0_bits_tail,
  input  [63:0] auto_dest_nodes_in_0_flit_0_bits_payload,
  input  [1:0]  auto_dest_nodes_in_0_flit_0_bits_flow_ingress_node,
  input  [1:0]  auto_dest_nodes_in_0_flit_0_bits_flow_egress_node,
  input  [1:0]  auto_dest_nodes_in_0_flit_0_bits_virt_channel_id,
  output [3:0]  auto_dest_nodes_in_0_credit_return,
  output [3:0]  auto_dest_nodes_in_0_vc_free
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_REG_INIT
  wire  monitor_clock; // @[Nodes.scala 24:25]
  wire  monitor_reset; // @[Nodes.scala 24:25]
  wire  monitor_io_in_flit_0_valid; // @[Nodes.scala 24:25]
  wire  monitor_io_in_flit_0_bits_head; // @[Nodes.scala 24:25]
  wire  monitor_io_in_flit_0_bits_tail; // @[Nodes.scala 24:25]
  wire [1:0] monitor_io_in_flit_0_bits_flow_ingress_node; // @[Nodes.scala 24:25]
  wire [1:0] monitor_io_in_flit_0_bits_flow_egress_node; // @[Nodes.scala 24:25]
  wire [1:0] monitor_io_in_flit_0_bits_virt_channel_id; // @[Nodes.scala 24:25]
  wire  monitor_1_clock; // @[Nodes.scala 24:25]
  wire  monitor_1_reset; // @[Nodes.scala 24:25]
  wire  monitor_1_io_in_flit_0_valid; // @[Nodes.scala 24:25]
  wire  monitor_1_io_in_flit_0_bits_head; // @[Nodes.scala 24:25]
  wire  monitor_1_io_in_flit_0_bits_tail; // @[Nodes.scala 24:25]
  wire [1:0] monitor_1_io_in_flit_0_bits_flow_ingress_node; // @[Nodes.scala 24:25]
  wire [1:0] monitor_1_io_in_flit_0_bits_flow_egress_node; // @[Nodes.scala 24:25]
  wire [1:0] monitor_1_io_in_flit_0_bits_virt_channel_id; // @[Nodes.scala 24:25]
  wire  input_unit_0_from_0_clock; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_reset; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_router_req_valid; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_0_io_router_req_bits_src_virt_id; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_0_io_router_req_bits_flow_ingress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_0_io_router_req_bits_flow_egress_node; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_router_resp_vc_sel_1_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_router_resp_vc_sel_1_1; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_router_resp_vc_sel_1_2; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_router_resp_vc_sel_1_3; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_router_resp_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_router_resp_vc_sel_0_1; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_router_resp_vc_sel_0_2; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_req_ready; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_req_valid; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_2_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_1_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_1_1; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_1_2; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_1_3; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_1; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_2; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_resp_vc_sel_2_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_resp_vc_sel_1_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_resp_vc_sel_1_1; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_resp_vc_sel_1_2; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_resp_vc_sel_1_3; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_resp_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_resp_vc_sel_0_1; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_resp_vc_sel_0_2; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_out_credit_available_2_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_out_credit_available_1_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_out_credit_available_1_1; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_out_credit_available_1_2; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_out_credit_available_1_3; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_out_credit_available_0_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_out_credit_available_0_1; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_out_credit_available_0_2; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_out_credit_available_0_3; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_salloc_req_0_ready; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_salloc_req_0_valid; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_2_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_1_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_1_1; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_1_2; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_1_3; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_1; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_2; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_3; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_salloc_req_0_bits_tail; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_out_0_valid; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_out_0_bits_flit_head; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_out_0_bits_flit_tail; // @[Router.scala 112:13]
  wire [63:0] input_unit_0_from_0_io_out_0_bits_flit_payload; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_0_io_out_0_bits_flit_flow_ingress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_0_io_out_0_bits_flit_flow_egress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_0_io_out_0_bits_out_virt_channel; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_0_io_debug_va_stall; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_0_io_debug_sa_stall; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_in_flit_0_valid; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_in_flit_0_bits_head; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_in_flit_0_bits_tail; // @[Router.scala 112:13]
  wire [63:0] input_unit_0_from_0_io_in_flit_0_bits_payload; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_0_io_in_flit_0_bits_flow_ingress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_0_io_in_flit_0_bits_flow_egress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_0_io_in_flit_0_bits_virt_channel_id; // @[Router.scala 112:13]
  wire [3:0] input_unit_0_from_0_io_in_credit_return; // @[Router.scala 112:13]
  wire [3:0] input_unit_0_from_0_io_in_vc_free; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_clock; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_reset; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_router_req_valid; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_2_io_router_req_bits_src_virt_id; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_2_io_router_req_bits_flow_ingress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_2_io_router_req_bits_flow_egress_node; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_router_resp_vc_sel_1_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_router_resp_vc_sel_1_1; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_router_resp_vc_sel_1_2; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_router_resp_vc_sel_1_3; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_router_resp_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_router_resp_vc_sel_0_1; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_router_resp_vc_sel_0_2; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_req_ready; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_req_valid; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_2_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_1_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_1_1; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_1_2; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_1_3; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_0_1; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_0_2; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_resp_vc_sel_2_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_resp_vc_sel_1_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_resp_vc_sel_1_1; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_resp_vc_sel_1_2; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_resp_vc_sel_1_3; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_resp_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_resp_vc_sel_0_1; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_resp_vc_sel_0_2; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_out_credit_available_2_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_out_credit_available_1_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_out_credit_available_1_1; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_out_credit_available_1_2; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_out_credit_available_1_3; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_out_credit_available_0_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_out_credit_available_0_1; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_out_credit_available_0_2; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_out_credit_available_0_3; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_salloc_req_0_ready; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_salloc_req_0_valid; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_2_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_1_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_1_1; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_1_2; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_1_3; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_0_1; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_0_2; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_0_3; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_salloc_req_0_bits_tail; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_out_0_valid; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_out_0_bits_flit_head; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_out_0_bits_flit_tail; // @[Router.scala 112:13]
  wire [63:0] input_unit_1_from_2_io_out_0_bits_flit_payload; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_2_io_out_0_bits_flit_flow_ingress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_2_io_out_0_bits_flit_flow_egress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_2_io_out_0_bits_out_virt_channel; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_2_io_debug_va_stall; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_2_io_debug_sa_stall; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_in_flit_0_valid; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_in_flit_0_bits_head; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_in_flit_0_bits_tail; // @[Router.scala 112:13]
  wire [63:0] input_unit_1_from_2_io_in_flit_0_bits_payload; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_2_io_in_flit_0_bits_flow_ingress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_2_io_in_flit_0_bits_flow_egress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_2_io_in_flit_0_bits_virt_channel_id; // @[Router.scala 112:13]
  wire [3:0] input_unit_1_from_2_io_in_credit_return; // @[Router.scala 112:13]
  wire [3:0] input_unit_1_from_2_io_in_vc_free; // @[Router.scala 112:13]
  wire  ingress_unit_2_from_3_clock; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_reset; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_router_req_valid; // @[Router.scala 116:13]
  wire [1:0] ingress_unit_2_from_3_io_router_req_bits_flow_ingress_node; // @[Router.scala 116:13]
  wire [1:0] ingress_unit_2_from_3_io_router_req_bits_flow_egress_node; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_router_resp_vc_sel_1_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_router_resp_vc_sel_1_1; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_router_resp_vc_sel_1_2; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_router_resp_vc_sel_1_3; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_router_resp_vc_sel_0_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_router_resp_vc_sel_0_1; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_router_resp_vc_sel_0_2; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_router_resp_vc_sel_0_3; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_vcalloc_req_ready; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_vcalloc_req_valid; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_vcalloc_req_bits_vc_sel_2_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_vcalloc_req_bits_vc_sel_1_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_vcalloc_req_bits_vc_sel_1_1; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_vcalloc_req_bits_vc_sel_1_2; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_vcalloc_req_bits_vc_sel_1_3; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_vcalloc_req_bits_vc_sel_0_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_vcalloc_req_bits_vc_sel_0_1; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_vcalloc_req_bits_vc_sel_0_2; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_vcalloc_req_bits_vc_sel_0_3; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_vcalloc_resp_vc_sel_2_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_vcalloc_resp_vc_sel_1_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_vcalloc_resp_vc_sel_1_1; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_vcalloc_resp_vc_sel_1_2; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_vcalloc_resp_vc_sel_1_3; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_vcalloc_resp_vc_sel_0_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_vcalloc_resp_vc_sel_0_1; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_vcalloc_resp_vc_sel_0_2; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_vcalloc_resp_vc_sel_0_3; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_out_credit_available_2_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_out_credit_available_1_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_out_credit_available_1_1; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_out_credit_available_1_2; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_out_credit_available_1_3; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_out_credit_available_0_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_out_credit_available_0_1; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_out_credit_available_0_2; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_out_credit_available_0_3; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_salloc_req_0_ready; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_salloc_req_0_valid; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_salloc_req_0_bits_vc_sel_2_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_salloc_req_0_bits_vc_sel_1_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_salloc_req_0_bits_vc_sel_1_1; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_salloc_req_0_bits_vc_sel_1_2; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_salloc_req_0_bits_vc_sel_1_3; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_salloc_req_0_bits_vc_sel_0_0; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_salloc_req_0_bits_vc_sel_0_1; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_salloc_req_0_bits_vc_sel_0_2; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_salloc_req_0_bits_vc_sel_0_3; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_salloc_req_0_bits_tail; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_out_0_valid; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_out_0_bits_flit_head; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_out_0_bits_flit_tail; // @[Router.scala 116:13]
  wire [63:0] ingress_unit_2_from_3_io_out_0_bits_flit_payload; // @[Router.scala 116:13]
  wire [1:0] ingress_unit_2_from_3_io_out_0_bits_flit_flow_ingress_node; // @[Router.scala 116:13]
  wire [1:0] ingress_unit_2_from_3_io_out_0_bits_flit_flow_egress_node; // @[Router.scala 116:13]
  wire [1:0] ingress_unit_2_from_3_io_out_0_bits_out_virt_channel; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_in_ready; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_in_valid; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_in_bits_head; // @[Router.scala 116:13]
  wire  ingress_unit_2_from_3_io_in_bits_tail; // @[Router.scala 116:13]
  wire [63:0] ingress_unit_2_from_3_io_in_bits_payload; // @[Router.scala 116:13]
  wire [1:0] ingress_unit_2_from_3_io_in_bits_egress_id; // @[Router.scala 116:13]
  wire  output_unit_0_to_0_clock; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_reset; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_in_0_valid; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_in_0_bits_head; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_in_0_bits_tail; // @[Router.scala 122:13]
  wire [63:0] output_unit_0_to_0_io_in_0_bits_payload; // @[Router.scala 122:13]
  wire [1:0] output_unit_0_to_0_io_in_0_bits_flow_ingress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_0_to_0_io_in_0_bits_flow_egress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_0_to_0_io_in_0_bits_virt_channel_id; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_credit_available_0; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_credit_available_1; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_credit_available_2; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_credit_available_3; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_channel_status_0_occupied; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_channel_status_1_occupied; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_channel_status_2_occupied; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_channel_status_3_occupied; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_allocs_0_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_allocs_1_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_allocs_2_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_allocs_3_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_credit_alloc_0_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_credit_alloc_1_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_credit_alloc_2_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_credit_alloc_3_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_out_flit_0_valid; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_out_flit_0_bits_head; // @[Router.scala 122:13]
  wire  output_unit_0_to_0_io_out_flit_0_bits_tail; // @[Router.scala 122:13]
  wire [63:0] output_unit_0_to_0_io_out_flit_0_bits_payload; // @[Router.scala 122:13]
  wire [1:0] output_unit_0_to_0_io_out_flit_0_bits_flow_ingress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_0_to_0_io_out_flit_0_bits_flow_egress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_0_to_0_io_out_flit_0_bits_virt_channel_id; // @[Router.scala 122:13]
  wire [3:0] output_unit_0_to_0_io_out_credit_return; // @[Router.scala 122:13]
  wire [3:0] output_unit_0_to_0_io_out_vc_free; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_clock; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_reset; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_in_0_valid; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_in_0_bits_head; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_in_0_bits_tail; // @[Router.scala 122:13]
  wire [63:0] output_unit_1_to_2_io_in_0_bits_payload; // @[Router.scala 122:13]
  wire [1:0] output_unit_1_to_2_io_in_0_bits_flow_ingress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_1_to_2_io_in_0_bits_flow_egress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_1_to_2_io_in_0_bits_virt_channel_id; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_credit_available_0; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_credit_available_1; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_credit_available_2; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_credit_available_3; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_channel_status_0_occupied; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_channel_status_1_occupied; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_channel_status_2_occupied; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_channel_status_3_occupied; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_allocs_0_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_allocs_1_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_allocs_2_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_allocs_3_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_credit_alloc_0_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_credit_alloc_1_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_credit_alloc_2_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_credit_alloc_3_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_out_flit_0_valid; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_out_flit_0_bits_head; // @[Router.scala 122:13]
  wire  output_unit_1_to_2_io_out_flit_0_bits_tail; // @[Router.scala 122:13]
  wire [63:0] output_unit_1_to_2_io_out_flit_0_bits_payload; // @[Router.scala 122:13]
  wire [1:0] output_unit_1_to_2_io_out_flit_0_bits_flow_ingress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_1_to_2_io_out_flit_0_bits_flow_egress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_1_to_2_io_out_flit_0_bits_virt_channel_id; // @[Router.scala 122:13]
  wire [3:0] output_unit_1_to_2_io_out_credit_return; // @[Router.scala 122:13]
  wire [3:0] output_unit_1_to_2_io_out_vc_free; // @[Router.scala 122:13]
  wire  egress_unit_2_to_3_clock; // @[Router.scala 125:13]
  wire  egress_unit_2_to_3_reset; // @[Router.scala 125:13]
  wire  egress_unit_2_to_3_io_in_0_valid; // @[Router.scala 125:13]
  wire  egress_unit_2_to_3_io_in_0_bits_head; // @[Router.scala 125:13]
  wire  egress_unit_2_to_3_io_in_0_bits_tail; // @[Router.scala 125:13]
  wire [63:0] egress_unit_2_to_3_io_in_0_bits_payload; // @[Router.scala 125:13]
  wire [1:0] egress_unit_2_to_3_io_in_0_bits_flow_ingress_node; // @[Router.scala 125:13]
  wire  egress_unit_2_to_3_io_credit_available_0; // @[Router.scala 125:13]
  wire  egress_unit_2_to_3_io_channel_status_0_occupied; // @[Router.scala 125:13]
  wire  egress_unit_2_to_3_io_allocs_0_alloc; // @[Router.scala 125:13]
  wire  egress_unit_2_to_3_io_credit_alloc_0_alloc; // @[Router.scala 125:13]
  wire  egress_unit_2_to_3_io_credit_alloc_0_tail; // @[Router.scala 125:13]
  wire  egress_unit_2_to_3_io_out_valid; // @[Router.scala 125:13]
  wire  egress_unit_2_to_3_io_out_bits_head; // @[Router.scala 125:13]
  wire  egress_unit_2_to_3_io_out_bits_tail; // @[Router.scala 125:13]
  wire [63:0] egress_unit_2_to_3_io_out_bits_payload; // @[Router.scala 125:13]
  wire [1:0] egress_unit_2_to_3_io_out_bits_ingress_id; // @[Router.scala 125:13]
  wire  switch_clock; // @[Router.scala 129:24]
  wire  switch_reset; // @[Router.scala 129:24]
  wire  switch_io_in_2_0_valid; // @[Router.scala 129:24]
  wire  switch_io_in_2_0_bits_flit_head; // @[Router.scala 129:24]
  wire  switch_io_in_2_0_bits_flit_tail; // @[Router.scala 129:24]
  wire [63:0] switch_io_in_2_0_bits_flit_payload; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_2_0_bits_flit_flow_ingress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_2_0_bits_flit_flow_egress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_2_0_bits_out_virt_channel; // @[Router.scala 129:24]
  wire  switch_io_in_1_0_valid; // @[Router.scala 129:24]
  wire  switch_io_in_1_0_bits_flit_head; // @[Router.scala 129:24]
  wire  switch_io_in_1_0_bits_flit_tail; // @[Router.scala 129:24]
  wire [63:0] switch_io_in_1_0_bits_flit_payload; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_1_0_bits_flit_flow_ingress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_1_0_bits_flit_flow_egress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_1_0_bits_out_virt_channel; // @[Router.scala 129:24]
  wire  switch_io_in_0_0_valid; // @[Router.scala 129:24]
  wire  switch_io_in_0_0_bits_flit_head; // @[Router.scala 129:24]
  wire  switch_io_in_0_0_bits_flit_tail; // @[Router.scala 129:24]
  wire [63:0] switch_io_in_0_0_bits_flit_payload; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_0_0_bits_flit_flow_ingress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_0_0_bits_flit_flow_egress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_0_0_bits_out_virt_channel; // @[Router.scala 129:24]
  wire  switch_io_out_2_0_valid; // @[Router.scala 129:24]
  wire  switch_io_out_2_0_bits_head; // @[Router.scala 129:24]
  wire  switch_io_out_2_0_bits_tail; // @[Router.scala 129:24]
  wire [63:0] switch_io_out_2_0_bits_payload; // @[Router.scala 129:24]
  wire [1:0] switch_io_out_2_0_bits_flow_ingress_node; // @[Router.scala 129:24]
  wire  switch_io_out_1_0_valid; // @[Router.scala 129:24]
  wire  switch_io_out_1_0_bits_head; // @[Router.scala 129:24]
  wire  switch_io_out_1_0_bits_tail; // @[Router.scala 129:24]
  wire [63:0] switch_io_out_1_0_bits_payload; // @[Router.scala 129:24]
  wire [1:0] switch_io_out_1_0_bits_flow_ingress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_out_1_0_bits_flow_egress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_out_1_0_bits_virt_channel_id; // @[Router.scala 129:24]
  wire  switch_io_out_0_0_valid; // @[Router.scala 129:24]
  wire  switch_io_out_0_0_bits_head; // @[Router.scala 129:24]
  wire  switch_io_out_0_0_bits_tail; // @[Router.scala 129:24]
  wire [63:0] switch_io_out_0_0_bits_payload; // @[Router.scala 129:24]
  wire [1:0] switch_io_out_0_0_bits_flow_ingress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_out_0_0_bits_flow_egress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_out_0_0_bits_virt_channel_id; // @[Router.scala 129:24]
  wire  switch_io_sel_2_0_2_0; // @[Router.scala 129:24]
  wire  switch_io_sel_2_0_1_0; // @[Router.scala 129:24]
  wire  switch_io_sel_2_0_0_0; // @[Router.scala 129:24]
  wire  switch_io_sel_1_0_2_0; // @[Router.scala 129:24]
  wire  switch_io_sel_1_0_1_0; // @[Router.scala 129:24]
  wire  switch_io_sel_1_0_0_0; // @[Router.scala 129:24]
  wire  switch_io_sel_0_0_2_0; // @[Router.scala 129:24]
  wire  switch_io_sel_0_0_1_0; // @[Router.scala 129:24]
  wire  switch_io_sel_0_0_0_0; // @[Router.scala 129:24]
  wire  switch_allocator_clock; // @[Router.scala 130:34]
  wire  switch_allocator_reset; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_ready; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_valid; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_bits_vc_sel_2_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_bits_vc_sel_1_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_bits_vc_sel_1_1; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_bits_vc_sel_1_2; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_bits_vc_sel_1_3; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_bits_vc_sel_0_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_bits_vc_sel_0_1; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_bits_vc_sel_0_2; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_bits_vc_sel_0_3; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_2_0_bits_tail; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_ready; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_valid; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_vc_sel_2_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_vc_sel_1_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_vc_sel_1_1; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_vc_sel_1_2; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_vc_sel_1_3; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_vc_sel_0_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_vc_sel_0_1; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_vc_sel_0_2; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_vc_sel_0_3; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_tail; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_ready; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_valid; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_2_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_1_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_1_1; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_1_2; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_1_3; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_0_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_0_1; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_0_2; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_0_3; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_tail; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_2_0_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_2_0_tail; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_1_0_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_1_1_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_1_2_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_1_3_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_0_0_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_0_1_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_0_2_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_0_3_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_2_0_2_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_2_0_1_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_2_0_0_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_1_0_2_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_1_0_1_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_1_0_0_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_0_0_2_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_0_0_1_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_0_0_0_0; // @[Router.scala 130:34]
  wire  vc_allocator_clock; // @[Router.scala 131:30]
  wire  vc_allocator_reset; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_ready; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_valid; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_bits_vc_sel_2_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_bits_vc_sel_1_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_bits_vc_sel_1_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_bits_vc_sel_1_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_bits_vc_sel_1_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_bits_vc_sel_0_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_bits_vc_sel_0_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_bits_vc_sel_0_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_2_bits_vc_sel_0_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_ready; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_valid; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_bits_vc_sel_2_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_bits_vc_sel_1_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_bits_vc_sel_1_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_bits_vc_sel_1_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_bits_vc_sel_1_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_bits_vc_sel_0_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_bits_vc_sel_0_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_bits_vc_sel_0_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_bits_vc_sel_0_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_ready; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_valid; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_2_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_1_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_1_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_1_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_1_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_0_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_0_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_0_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_0_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_2_vc_sel_2_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_2_vc_sel_1_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_2_vc_sel_1_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_2_vc_sel_1_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_2_vc_sel_1_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_2_vc_sel_0_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_2_vc_sel_0_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_2_vc_sel_0_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_2_vc_sel_0_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_1_vc_sel_2_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_1_vc_sel_1_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_1_vc_sel_1_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_1_vc_sel_1_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_1_vc_sel_1_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_1_vc_sel_0_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_1_vc_sel_0_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_1_vc_sel_0_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_1_vc_sel_0_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_2_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_1_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_1_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_1_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_1_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_0_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_0_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_0_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_0_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_2_0_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_1_0_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_1_1_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_1_2_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_1_3_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_0_0_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_0_1_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_0_2_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_0_3_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_2_0_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_1_0_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_1_1_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_1_2_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_1_3_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_0_0_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_0_1_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_0_2_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_0_3_alloc; // @[Router.scala 131:30]
  wire [1:0] route_computer_io_req_2_bits_flow_ingress_node; // @[Router.scala 134:32]
  wire [1:0] route_computer_io_req_2_bits_flow_egress_node; // @[Router.scala 134:32]
  wire [1:0] route_computer_io_req_1_bits_src_virt_id; // @[Router.scala 134:32]
  wire [1:0] route_computer_io_req_1_bits_flow_ingress_node; // @[Router.scala 134:32]
  wire [1:0] route_computer_io_req_1_bits_flow_egress_node; // @[Router.scala 134:32]
  wire [1:0] route_computer_io_req_0_bits_src_virt_id; // @[Router.scala 134:32]
  wire [1:0] route_computer_io_req_0_bits_flow_ingress_node; // @[Router.scala 134:32]
  wire [1:0] route_computer_io_req_0_bits_flow_egress_node; // @[Router.scala 134:32]
  wire  route_computer_io_resp_2_vc_sel_1_0; // @[Router.scala 134:32]
  wire  route_computer_io_resp_2_vc_sel_1_1; // @[Router.scala 134:32]
  wire  route_computer_io_resp_2_vc_sel_1_2; // @[Router.scala 134:32]
  wire  route_computer_io_resp_2_vc_sel_1_3; // @[Router.scala 134:32]
  wire  route_computer_io_resp_2_vc_sel_0_0; // @[Router.scala 134:32]
  wire  route_computer_io_resp_2_vc_sel_0_1; // @[Router.scala 134:32]
  wire  route_computer_io_resp_2_vc_sel_0_2; // @[Router.scala 134:32]
  wire  route_computer_io_resp_2_vc_sel_0_3; // @[Router.scala 134:32]
  wire  route_computer_io_resp_1_vc_sel_1_0; // @[Router.scala 134:32]
  wire  route_computer_io_resp_1_vc_sel_1_1; // @[Router.scala 134:32]
  wire  route_computer_io_resp_1_vc_sel_1_2; // @[Router.scala 134:32]
  wire  route_computer_io_resp_1_vc_sel_1_3; // @[Router.scala 134:32]
  wire  route_computer_io_resp_1_vc_sel_0_0; // @[Router.scala 134:32]
  wire  route_computer_io_resp_1_vc_sel_0_1; // @[Router.scala 134:32]
  wire  route_computer_io_resp_1_vc_sel_0_2; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_1_0; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_1_1; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_1_2; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_1_3; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_0_0; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_0_1; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_0_2; // @[Router.scala 134:32]
  wire [19:0] plusarg_reader_out; // @[PlusArg.scala 80:11]
  wire  _fires_count_T = vc_allocator_io_req_0_ready & vc_allocator_io_req_0_valid; // @[Decoupled.scala 51:35]
  wire  _fires_count_T_1 = vc_allocator_io_req_1_ready & vc_allocator_io_req_1_valid; // @[Decoupled.scala 51:35]
  wire  _fires_count_T_2 = vc_allocator_io_req_2_ready & vc_allocator_io_req_2_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _fires_count_T_3 = _fires_count_T_1 + _fires_count_T_2; // @[Bitwise.scala 51:90]
  wire [1:0] _GEN_5 = {{1'd0}, _fires_count_T}; // @[Bitwise.scala 51:90]
  wire [2:0] _fires_count_T_5 = _GEN_5 + _fires_count_T_3; // @[Bitwise.scala 51:90]
  reg  switch_io_sel_REG_2_0_2_0; // @[Router.scala 176:14]
  reg  switch_io_sel_REG_2_0_1_0; // @[Router.scala 176:14]
  reg  switch_io_sel_REG_2_0_0_0; // @[Router.scala 176:14]
  reg  switch_io_sel_REG_1_0_2_0; // @[Router.scala 176:14]
  reg  switch_io_sel_REG_1_0_1_0; // @[Router.scala 176:14]
  reg  switch_io_sel_REG_1_0_0_0; // @[Router.scala 176:14]
  reg  switch_io_sel_REG_0_0_2_0; // @[Router.scala 176:14]
  reg  switch_io_sel_REG_0_0_1_0; // @[Router.scala 176:14]
  reg  switch_io_sel_REG_0_0_0_0; // @[Router.scala 176:14]
  reg [63:0] debug_tsc; // @[Router.scala 193:28]
  wire [63:0] _debug_tsc_T_1 = debug_tsc + 64'h1; // @[Router.scala 194:28]
  reg [63:0] debug_sample; // @[Router.scala 195:31]
  wire [63:0] _debug_sample_T_1 = debug_sample + 64'h1; // @[Router.scala 196:34]
  wire [19:0] _T_1 = plusarg_reader_out - 20'h1; // @[Router.scala 198:40]
  wire [63:0] _GEN_6 = {{44'd0}, _T_1}; // @[Router.scala 198:24]
  wire  _T_2 = debug_sample == _GEN_6; // @[Router.scala 198:24]
  reg [63:0] util_ctr; // @[Router.scala 201:29]
  reg  fired; // @[Router.scala 202:26]
  wire [63:0] _GEN_7 = {{63'd0}, auto_dest_nodes_in_0_flit_0_valid}; // @[Router.scala 203:28]
  wire [63:0] _util_ctr_T_1 = util_ctr + _GEN_7; // @[Router.scala 203:28]
  wire  _T_8 = plusarg_reader_out != 20'h0 & _T_2 & fired; // @[Router.scala 205:71]
  reg [63:0] util_ctr_1; // @[Router.scala 201:29]
  reg  fired_1; // @[Router.scala 202:26]
  wire [63:0] _GEN_9 = {{63'd0}, auto_dest_nodes_in_1_flit_0_valid}; // @[Router.scala 203:28]
  wire [63:0] _util_ctr_T_3 = util_ctr_1 + _GEN_9; // @[Router.scala 203:28]
  wire  _T_16 = plusarg_reader_out != 20'h0 & _T_2 & fired_1; // @[Router.scala 205:71]
  wire  bundleIn_0_2_flit_ready = ingress_unit_2_from_3_io_in_ready; // @[Nodes.scala 1215:84 Router.scala 142:68]
  wire  _T_19 = bundleIn_0_2_flit_ready & auto_ingress_nodes_in_flit_valid; // @[Decoupled.scala 51:35]
  reg [63:0] util_ctr_2; // @[Router.scala 201:29]
  reg  fired_2; // @[Router.scala 202:26]
  wire [63:0] _GEN_11 = {{63'd0}, _T_19}; // @[Router.scala 203:28]
  wire [63:0] _util_ctr_T_5 = util_ctr_2 + _GEN_11; // @[Router.scala 203:28]
  wire  _T_25 = plusarg_reader_out != 20'h0 & _T_2 & fired_2; // @[Router.scala 205:71]
  wire  x1_2_flit_valid = egress_unit_2_to_3_io_out_valid; // @[Nodes.scala 1212:84 Router.scala 144:65]
  reg [63:0] util_ctr_3; // @[Router.scala 201:29]
  reg  fired_3; // @[Router.scala 202:26]
  wire [63:0] _GEN_13 = {{63'd0}, x1_2_flit_valid}; // @[Router.scala 203:28]
  wire [63:0] _util_ctr_T_7 = util_ctr_3 + _GEN_13; // @[Router.scala 203:28]
  wire  _T_34 = plusarg_reader_out != 20'h0 & _T_2 & fired_3; // @[Router.scala 205:71]
  wire [1:0] fires_count = _fires_count_T_5[1:0]; // @[Bitwise.scala 51:90]
  NoCMonitor_6 monitor ( // @[Nodes.scala 24:25]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_flit_0_valid(monitor_io_in_flit_0_valid),
    .io_in_flit_0_bits_head(monitor_io_in_flit_0_bits_head),
    .io_in_flit_0_bits_tail(monitor_io_in_flit_0_bits_tail),
    .io_in_flit_0_bits_flow_ingress_node(monitor_io_in_flit_0_bits_flow_ingress_node),
    .io_in_flit_0_bits_flow_egress_node(monitor_io_in_flit_0_bits_flow_egress_node),
    .io_in_flit_0_bits_virt_channel_id(monitor_io_in_flit_0_bits_virt_channel_id)
  );
  NoCMonitor_7 monitor_1 ( // @[Nodes.scala 24:25]
    .clock(monitor_1_clock),
    .reset(monitor_1_reset),
    .io_in_flit_0_valid(monitor_1_io_in_flit_0_valid),
    .io_in_flit_0_bits_head(monitor_1_io_in_flit_0_bits_head),
    .io_in_flit_0_bits_tail(monitor_1_io_in_flit_0_bits_tail),
    .io_in_flit_0_bits_flow_ingress_node(monitor_1_io_in_flit_0_bits_flow_ingress_node),
    .io_in_flit_0_bits_flow_egress_node(monitor_1_io_in_flit_0_bits_flow_egress_node),
    .io_in_flit_0_bits_virt_channel_id(monitor_1_io_in_flit_0_bits_virt_channel_id)
  );
  InputUnit_6 input_unit_0_from_0 ( // @[Router.scala 112:13]
    .clock(input_unit_0_from_0_clock),
    .reset(input_unit_0_from_0_reset),
    .io_router_req_valid(input_unit_0_from_0_io_router_req_valid),
    .io_router_req_bits_src_virt_id(input_unit_0_from_0_io_router_req_bits_src_virt_id),
    .io_router_req_bits_flow_ingress_node(input_unit_0_from_0_io_router_req_bits_flow_ingress_node),
    .io_router_req_bits_flow_egress_node(input_unit_0_from_0_io_router_req_bits_flow_egress_node),
    .io_router_resp_vc_sel_1_0(input_unit_0_from_0_io_router_resp_vc_sel_1_0),
    .io_router_resp_vc_sel_1_1(input_unit_0_from_0_io_router_resp_vc_sel_1_1),
    .io_router_resp_vc_sel_1_2(input_unit_0_from_0_io_router_resp_vc_sel_1_2),
    .io_router_resp_vc_sel_1_3(input_unit_0_from_0_io_router_resp_vc_sel_1_3),
    .io_router_resp_vc_sel_0_0(input_unit_0_from_0_io_router_resp_vc_sel_0_0),
    .io_router_resp_vc_sel_0_1(input_unit_0_from_0_io_router_resp_vc_sel_0_1),
    .io_router_resp_vc_sel_0_2(input_unit_0_from_0_io_router_resp_vc_sel_0_2),
    .io_vcalloc_req_ready(input_unit_0_from_0_io_vcalloc_req_ready),
    .io_vcalloc_req_valid(input_unit_0_from_0_io_vcalloc_req_valid),
    .io_vcalloc_req_bits_vc_sel_2_0(input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_2_0),
    .io_vcalloc_req_bits_vc_sel_1_0(input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_1_0),
    .io_vcalloc_req_bits_vc_sel_1_1(input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_1_1),
    .io_vcalloc_req_bits_vc_sel_1_2(input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_1_2),
    .io_vcalloc_req_bits_vc_sel_1_3(input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_1_3),
    .io_vcalloc_req_bits_vc_sel_0_0(input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_0),
    .io_vcalloc_req_bits_vc_sel_0_1(input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_1),
    .io_vcalloc_req_bits_vc_sel_0_2(input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_2),
    .io_vcalloc_resp_vc_sel_2_0(input_unit_0_from_0_io_vcalloc_resp_vc_sel_2_0),
    .io_vcalloc_resp_vc_sel_1_0(input_unit_0_from_0_io_vcalloc_resp_vc_sel_1_0),
    .io_vcalloc_resp_vc_sel_1_1(input_unit_0_from_0_io_vcalloc_resp_vc_sel_1_1),
    .io_vcalloc_resp_vc_sel_1_2(input_unit_0_from_0_io_vcalloc_resp_vc_sel_1_2),
    .io_vcalloc_resp_vc_sel_1_3(input_unit_0_from_0_io_vcalloc_resp_vc_sel_1_3),
    .io_vcalloc_resp_vc_sel_0_0(input_unit_0_from_0_io_vcalloc_resp_vc_sel_0_0),
    .io_vcalloc_resp_vc_sel_0_1(input_unit_0_from_0_io_vcalloc_resp_vc_sel_0_1),
    .io_vcalloc_resp_vc_sel_0_2(input_unit_0_from_0_io_vcalloc_resp_vc_sel_0_2),
    .io_out_credit_available_2_0(input_unit_0_from_0_io_out_credit_available_2_0),
    .io_out_credit_available_1_0(input_unit_0_from_0_io_out_credit_available_1_0),
    .io_out_credit_available_1_1(input_unit_0_from_0_io_out_credit_available_1_1),
    .io_out_credit_available_1_2(input_unit_0_from_0_io_out_credit_available_1_2),
    .io_out_credit_available_1_3(input_unit_0_from_0_io_out_credit_available_1_3),
    .io_out_credit_available_0_0(input_unit_0_from_0_io_out_credit_available_0_0),
    .io_out_credit_available_0_1(input_unit_0_from_0_io_out_credit_available_0_1),
    .io_out_credit_available_0_2(input_unit_0_from_0_io_out_credit_available_0_2),
    .io_out_credit_available_0_3(input_unit_0_from_0_io_out_credit_available_0_3),
    .io_salloc_req_0_ready(input_unit_0_from_0_io_salloc_req_0_ready),
    .io_salloc_req_0_valid(input_unit_0_from_0_io_salloc_req_0_valid),
    .io_salloc_req_0_bits_vc_sel_2_0(input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_2_0),
    .io_salloc_req_0_bits_vc_sel_1_0(input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_1_0),
    .io_salloc_req_0_bits_vc_sel_1_1(input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_1_1),
    .io_salloc_req_0_bits_vc_sel_1_2(input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_1_2),
    .io_salloc_req_0_bits_vc_sel_1_3(input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_1_3),
    .io_salloc_req_0_bits_vc_sel_0_0(input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_0),
    .io_salloc_req_0_bits_vc_sel_0_1(input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_1),
    .io_salloc_req_0_bits_vc_sel_0_2(input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_2),
    .io_salloc_req_0_bits_vc_sel_0_3(input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_3),
    .io_salloc_req_0_bits_tail(input_unit_0_from_0_io_salloc_req_0_bits_tail),
    .io_out_0_valid(input_unit_0_from_0_io_out_0_valid),
    .io_out_0_bits_flit_head(input_unit_0_from_0_io_out_0_bits_flit_head),
    .io_out_0_bits_flit_tail(input_unit_0_from_0_io_out_0_bits_flit_tail),
    .io_out_0_bits_flit_payload(input_unit_0_from_0_io_out_0_bits_flit_payload),
    .io_out_0_bits_flit_flow_ingress_node(input_unit_0_from_0_io_out_0_bits_flit_flow_ingress_node),
    .io_out_0_bits_flit_flow_egress_node(input_unit_0_from_0_io_out_0_bits_flit_flow_egress_node),
    .io_out_0_bits_out_virt_channel(input_unit_0_from_0_io_out_0_bits_out_virt_channel),
    .io_debug_va_stall(input_unit_0_from_0_io_debug_va_stall),
    .io_debug_sa_stall(input_unit_0_from_0_io_debug_sa_stall),
    .io_in_flit_0_valid(input_unit_0_from_0_io_in_flit_0_valid),
    .io_in_flit_0_bits_head(input_unit_0_from_0_io_in_flit_0_bits_head),
    .io_in_flit_0_bits_tail(input_unit_0_from_0_io_in_flit_0_bits_tail),
    .io_in_flit_0_bits_payload(input_unit_0_from_0_io_in_flit_0_bits_payload),
    .io_in_flit_0_bits_flow_ingress_node(input_unit_0_from_0_io_in_flit_0_bits_flow_ingress_node),
    .io_in_flit_0_bits_flow_egress_node(input_unit_0_from_0_io_in_flit_0_bits_flow_egress_node),
    .io_in_flit_0_bits_virt_channel_id(input_unit_0_from_0_io_in_flit_0_bits_virt_channel_id),
    .io_in_credit_return(input_unit_0_from_0_io_in_credit_return),
    .io_in_vc_free(input_unit_0_from_0_io_in_vc_free)
  );
  InputUnit_7 input_unit_1_from_2 ( // @[Router.scala 112:13]
    .clock(input_unit_1_from_2_clock),
    .reset(input_unit_1_from_2_reset),
    .io_router_req_valid(input_unit_1_from_2_io_router_req_valid),
    .io_router_req_bits_src_virt_id(input_unit_1_from_2_io_router_req_bits_src_virt_id),
    .io_router_req_bits_flow_ingress_node(input_unit_1_from_2_io_router_req_bits_flow_ingress_node),
    .io_router_req_bits_flow_egress_node(input_unit_1_from_2_io_router_req_bits_flow_egress_node),
    .io_router_resp_vc_sel_1_0(input_unit_1_from_2_io_router_resp_vc_sel_1_0),
    .io_router_resp_vc_sel_1_1(input_unit_1_from_2_io_router_resp_vc_sel_1_1),
    .io_router_resp_vc_sel_1_2(input_unit_1_from_2_io_router_resp_vc_sel_1_2),
    .io_router_resp_vc_sel_1_3(input_unit_1_from_2_io_router_resp_vc_sel_1_3),
    .io_router_resp_vc_sel_0_0(input_unit_1_from_2_io_router_resp_vc_sel_0_0),
    .io_router_resp_vc_sel_0_1(input_unit_1_from_2_io_router_resp_vc_sel_0_1),
    .io_router_resp_vc_sel_0_2(input_unit_1_from_2_io_router_resp_vc_sel_0_2),
    .io_vcalloc_req_ready(input_unit_1_from_2_io_vcalloc_req_ready),
    .io_vcalloc_req_valid(input_unit_1_from_2_io_vcalloc_req_valid),
    .io_vcalloc_req_bits_vc_sel_2_0(input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_2_0),
    .io_vcalloc_req_bits_vc_sel_1_0(input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_1_0),
    .io_vcalloc_req_bits_vc_sel_1_1(input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_1_1),
    .io_vcalloc_req_bits_vc_sel_1_2(input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_1_2),
    .io_vcalloc_req_bits_vc_sel_1_3(input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_1_3),
    .io_vcalloc_req_bits_vc_sel_0_0(input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_0_0),
    .io_vcalloc_req_bits_vc_sel_0_1(input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_0_1),
    .io_vcalloc_req_bits_vc_sel_0_2(input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_0_2),
    .io_vcalloc_resp_vc_sel_2_0(input_unit_1_from_2_io_vcalloc_resp_vc_sel_2_0),
    .io_vcalloc_resp_vc_sel_1_0(input_unit_1_from_2_io_vcalloc_resp_vc_sel_1_0),
    .io_vcalloc_resp_vc_sel_1_1(input_unit_1_from_2_io_vcalloc_resp_vc_sel_1_1),
    .io_vcalloc_resp_vc_sel_1_2(input_unit_1_from_2_io_vcalloc_resp_vc_sel_1_2),
    .io_vcalloc_resp_vc_sel_1_3(input_unit_1_from_2_io_vcalloc_resp_vc_sel_1_3),
    .io_vcalloc_resp_vc_sel_0_0(input_unit_1_from_2_io_vcalloc_resp_vc_sel_0_0),
    .io_vcalloc_resp_vc_sel_0_1(input_unit_1_from_2_io_vcalloc_resp_vc_sel_0_1),
    .io_vcalloc_resp_vc_sel_0_2(input_unit_1_from_2_io_vcalloc_resp_vc_sel_0_2),
    .io_out_credit_available_2_0(input_unit_1_from_2_io_out_credit_available_2_0),
    .io_out_credit_available_1_0(input_unit_1_from_2_io_out_credit_available_1_0),
    .io_out_credit_available_1_1(input_unit_1_from_2_io_out_credit_available_1_1),
    .io_out_credit_available_1_2(input_unit_1_from_2_io_out_credit_available_1_2),
    .io_out_credit_available_1_3(input_unit_1_from_2_io_out_credit_available_1_3),
    .io_out_credit_available_0_0(input_unit_1_from_2_io_out_credit_available_0_0),
    .io_out_credit_available_0_1(input_unit_1_from_2_io_out_credit_available_0_1),
    .io_out_credit_available_0_2(input_unit_1_from_2_io_out_credit_available_0_2),
    .io_out_credit_available_0_3(input_unit_1_from_2_io_out_credit_available_0_3),
    .io_salloc_req_0_ready(input_unit_1_from_2_io_salloc_req_0_ready),
    .io_salloc_req_0_valid(input_unit_1_from_2_io_salloc_req_0_valid),
    .io_salloc_req_0_bits_vc_sel_2_0(input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_2_0),
    .io_salloc_req_0_bits_vc_sel_1_0(input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_1_0),
    .io_salloc_req_0_bits_vc_sel_1_1(input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_1_1),
    .io_salloc_req_0_bits_vc_sel_1_2(input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_1_2),
    .io_salloc_req_0_bits_vc_sel_1_3(input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_1_3),
    .io_salloc_req_0_bits_vc_sel_0_0(input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_0_0),
    .io_salloc_req_0_bits_vc_sel_0_1(input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_0_1),
    .io_salloc_req_0_bits_vc_sel_0_2(input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_0_2),
    .io_salloc_req_0_bits_vc_sel_0_3(input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_0_3),
    .io_salloc_req_0_bits_tail(input_unit_1_from_2_io_salloc_req_0_bits_tail),
    .io_out_0_valid(input_unit_1_from_2_io_out_0_valid),
    .io_out_0_bits_flit_head(input_unit_1_from_2_io_out_0_bits_flit_head),
    .io_out_0_bits_flit_tail(input_unit_1_from_2_io_out_0_bits_flit_tail),
    .io_out_0_bits_flit_payload(input_unit_1_from_2_io_out_0_bits_flit_payload),
    .io_out_0_bits_flit_flow_ingress_node(input_unit_1_from_2_io_out_0_bits_flit_flow_ingress_node),
    .io_out_0_bits_flit_flow_egress_node(input_unit_1_from_2_io_out_0_bits_flit_flow_egress_node),
    .io_out_0_bits_out_virt_channel(input_unit_1_from_2_io_out_0_bits_out_virt_channel),
    .io_debug_va_stall(input_unit_1_from_2_io_debug_va_stall),
    .io_debug_sa_stall(input_unit_1_from_2_io_debug_sa_stall),
    .io_in_flit_0_valid(input_unit_1_from_2_io_in_flit_0_valid),
    .io_in_flit_0_bits_head(input_unit_1_from_2_io_in_flit_0_bits_head),
    .io_in_flit_0_bits_tail(input_unit_1_from_2_io_in_flit_0_bits_tail),
    .io_in_flit_0_bits_payload(input_unit_1_from_2_io_in_flit_0_bits_payload),
    .io_in_flit_0_bits_flow_ingress_node(input_unit_1_from_2_io_in_flit_0_bits_flow_ingress_node),
    .io_in_flit_0_bits_flow_egress_node(input_unit_1_from_2_io_in_flit_0_bits_flow_egress_node),
    .io_in_flit_0_bits_virt_channel_id(input_unit_1_from_2_io_in_flit_0_bits_virt_channel_id),
    .io_in_credit_return(input_unit_1_from_2_io_in_credit_return),
    .io_in_vc_free(input_unit_1_from_2_io_in_vc_free)
  );
  IngressUnit_3 ingress_unit_2_from_3 ( // @[Router.scala 116:13]
    .clock(ingress_unit_2_from_3_clock),
    .reset(ingress_unit_2_from_3_reset),
    .io_router_req_valid(ingress_unit_2_from_3_io_router_req_valid),
    .io_router_req_bits_flow_ingress_node(ingress_unit_2_from_3_io_router_req_bits_flow_ingress_node),
    .io_router_req_bits_flow_egress_node(ingress_unit_2_from_3_io_router_req_bits_flow_egress_node),
    .io_router_resp_vc_sel_1_0(ingress_unit_2_from_3_io_router_resp_vc_sel_1_0),
    .io_router_resp_vc_sel_1_1(ingress_unit_2_from_3_io_router_resp_vc_sel_1_1),
    .io_router_resp_vc_sel_1_2(ingress_unit_2_from_3_io_router_resp_vc_sel_1_2),
    .io_router_resp_vc_sel_1_3(ingress_unit_2_from_3_io_router_resp_vc_sel_1_3),
    .io_router_resp_vc_sel_0_0(ingress_unit_2_from_3_io_router_resp_vc_sel_0_0),
    .io_router_resp_vc_sel_0_1(ingress_unit_2_from_3_io_router_resp_vc_sel_0_1),
    .io_router_resp_vc_sel_0_2(ingress_unit_2_from_3_io_router_resp_vc_sel_0_2),
    .io_router_resp_vc_sel_0_3(ingress_unit_2_from_3_io_router_resp_vc_sel_0_3),
    .io_vcalloc_req_ready(ingress_unit_2_from_3_io_vcalloc_req_ready),
    .io_vcalloc_req_valid(ingress_unit_2_from_3_io_vcalloc_req_valid),
    .io_vcalloc_req_bits_vc_sel_2_0(ingress_unit_2_from_3_io_vcalloc_req_bits_vc_sel_2_0),
    .io_vcalloc_req_bits_vc_sel_1_0(ingress_unit_2_from_3_io_vcalloc_req_bits_vc_sel_1_0),
    .io_vcalloc_req_bits_vc_sel_1_1(ingress_unit_2_from_3_io_vcalloc_req_bits_vc_sel_1_1),
    .io_vcalloc_req_bits_vc_sel_1_2(ingress_unit_2_from_3_io_vcalloc_req_bits_vc_sel_1_2),
    .io_vcalloc_req_bits_vc_sel_1_3(ingress_unit_2_from_3_io_vcalloc_req_bits_vc_sel_1_3),
    .io_vcalloc_req_bits_vc_sel_0_0(ingress_unit_2_from_3_io_vcalloc_req_bits_vc_sel_0_0),
    .io_vcalloc_req_bits_vc_sel_0_1(ingress_unit_2_from_3_io_vcalloc_req_bits_vc_sel_0_1),
    .io_vcalloc_req_bits_vc_sel_0_2(ingress_unit_2_from_3_io_vcalloc_req_bits_vc_sel_0_2),
    .io_vcalloc_req_bits_vc_sel_0_3(ingress_unit_2_from_3_io_vcalloc_req_bits_vc_sel_0_3),
    .io_vcalloc_resp_vc_sel_2_0(ingress_unit_2_from_3_io_vcalloc_resp_vc_sel_2_0),
    .io_vcalloc_resp_vc_sel_1_0(ingress_unit_2_from_3_io_vcalloc_resp_vc_sel_1_0),
    .io_vcalloc_resp_vc_sel_1_1(ingress_unit_2_from_3_io_vcalloc_resp_vc_sel_1_1),
    .io_vcalloc_resp_vc_sel_1_2(ingress_unit_2_from_3_io_vcalloc_resp_vc_sel_1_2),
    .io_vcalloc_resp_vc_sel_1_3(ingress_unit_2_from_3_io_vcalloc_resp_vc_sel_1_3),
    .io_vcalloc_resp_vc_sel_0_0(ingress_unit_2_from_3_io_vcalloc_resp_vc_sel_0_0),
    .io_vcalloc_resp_vc_sel_0_1(ingress_unit_2_from_3_io_vcalloc_resp_vc_sel_0_1),
    .io_vcalloc_resp_vc_sel_0_2(ingress_unit_2_from_3_io_vcalloc_resp_vc_sel_0_2),
    .io_vcalloc_resp_vc_sel_0_3(ingress_unit_2_from_3_io_vcalloc_resp_vc_sel_0_3),
    .io_out_credit_available_2_0(ingress_unit_2_from_3_io_out_credit_available_2_0),
    .io_out_credit_available_1_0(ingress_unit_2_from_3_io_out_credit_available_1_0),
    .io_out_credit_available_1_1(ingress_unit_2_from_3_io_out_credit_available_1_1),
    .io_out_credit_available_1_2(ingress_unit_2_from_3_io_out_credit_available_1_2),
    .io_out_credit_available_1_3(ingress_unit_2_from_3_io_out_credit_available_1_3),
    .io_out_credit_available_0_0(ingress_unit_2_from_3_io_out_credit_available_0_0),
    .io_out_credit_available_0_1(ingress_unit_2_from_3_io_out_credit_available_0_1),
    .io_out_credit_available_0_2(ingress_unit_2_from_3_io_out_credit_available_0_2),
    .io_out_credit_available_0_3(ingress_unit_2_from_3_io_out_credit_available_0_3),
    .io_salloc_req_0_ready(ingress_unit_2_from_3_io_salloc_req_0_ready),
    .io_salloc_req_0_valid(ingress_unit_2_from_3_io_salloc_req_0_valid),
    .io_salloc_req_0_bits_vc_sel_2_0(ingress_unit_2_from_3_io_salloc_req_0_bits_vc_sel_2_0),
    .io_salloc_req_0_bits_vc_sel_1_0(ingress_unit_2_from_3_io_salloc_req_0_bits_vc_sel_1_0),
    .io_salloc_req_0_bits_vc_sel_1_1(ingress_unit_2_from_3_io_salloc_req_0_bits_vc_sel_1_1),
    .io_salloc_req_0_bits_vc_sel_1_2(ingress_unit_2_from_3_io_salloc_req_0_bits_vc_sel_1_2),
    .io_salloc_req_0_bits_vc_sel_1_3(ingress_unit_2_from_3_io_salloc_req_0_bits_vc_sel_1_3),
    .io_salloc_req_0_bits_vc_sel_0_0(ingress_unit_2_from_3_io_salloc_req_0_bits_vc_sel_0_0),
    .io_salloc_req_0_bits_vc_sel_0_1(ingress_unit_2_from_3_io_salloc_req_0_bits_vc_sel_0_1),
    .io_salloc_req_0_bits_vc_sel_0_2(ingress_unit_2_from_3_io_salloc_req_0_bits_vc_sel_0_2),
    .io_salloc_req_0_bits_vc_sel_0_3(ingress_unit_2_from_3_io_salloc_req_0_bits_vc_sel_0_3),
    .io_salloc_req_0_bits_tail(ingress_unit_2_from_3_io_salloc_req_0_bits_tail),
    .io_out_0_valid(ingress_unit_2_from_3_io_out_0_valid),
    .io_out_0_bits_flit_head(ingress_unit_2_from_3_io_out_0_bits_flit_head),
    .io_out_0_bits_flit_tail(ingress_unit_2_from_3_io_out_0_bits_flit_tail),
    .io_out_0_bits_flit_payload(ingress_unit_2_from_3_io_out_0_bits_flit_payload),
    .io_out_0_bits_flit_flow_ingress_node(ingress_unit_2_from_3_io_out_0_bits_flit_flow_ingress_node),
    .io_out_0_bits_flit_flow_egress_node(ingress_unit_2_from_3_io_out_0_bits_flit_flow_egress_node),
    .io_out_0_bits_out_virt_channel(ingress_unit_2_from_3_io_out_0_bits_out_virt_channel),
    .io_in_ready(ingress_unit_2_from_3_io_in_ready),
    .io_in_valid(ingress_unit_2_from_3_io_in_valid),
    .io_in_bits_head(ingress_unit_2_from_3_io_in_bits_head),
    .io_in_bits_tail(ingress_unit_2_from_3_io_in_bits_tail),
    .io_in_bits_payload(ingress_unit_2_from_3_io_in_bits_payload),
    .io_in_bits_egress_id(ingress_unit_2_from_3_io_in_bits_egress_id)
  );
  OutputUnit output_unit_0_to_0 ( // @[Router.scala 122:13]
    .clock(output_unit_0_to_0_clock),
    .reset(output_unit_0_to_0_reset),
    .io_in_0_valid(output_unit_0_to_0_io_in_0_valid),
    .io_in_0_bits_head(output_unit_0_to_0_io_in_0_bits_head),
    .io_in_0_bits_tail(output_unit_0_to_0_io_in_0_bits_tail),
    .io_in_0_bits_payload(output_unit_0_to_0_io_in_0_bits_payload),
    .io_in_0_bits_flow_ingress_node(output_unit_0_to_0_io_in_0_bits_flow_ingress_node),
    .io_in_0_bits_flow_egress_node(output_unit_0_to_0_io_in_0_bits_flow_egress_node),
    .io_in_0_bits_virt_channel_id(output_unit_0_to_0_io_in_0_bits_virt_channel_id),
    .io_credit_available_0(output_unit_0_to_0_io_credit_available_0),
    .io_credit_available_1(output_unit_0_to_0_io_credit_available_1),
    .io_credit_available_2(output_unit_0_to_0_io_credit_available_2),
    .io_credit_available_3(output_unit_0_to_0_io_credit_available_3),
    .io_channel_status_0_occupied(output_unit_0_to_0_io_channel_status_0_occupied),
    .io_channel_status_1_occupied(output_unit_0_to_0_io_channel_status_1_occupied),
    .io_channel_status_2_occupied(output_unit_0_to_0_io_channel_status_2_occupied),
    .io_channel_status_3_occupied(output_unit_0_to_0_io_channel_status_3_occupied),
    .io_allocs_0_alloc(output_unit_0_to_0_io_allocs_0_alloc),
    .io_allocs_1_alloc(output_unit_0_to_0_io_allocs_1_alloc),
    .io_allocs_2_alloc(output_unit_0_to_0_io_allocs_2_alloc),
    .io_allocs_3_alloc(output_unit_0_to_0_io_allocs_3_alloc),
    .io_credit_alloc_0_alloc(output_unit_0_to_0_io_credit_alloc_0_alloc),
    .io_credit_alloc_1_alloc(output_unit_0_to_0_io_credit_alloc_1_alloc),
    .io_credit_alloc_2_alloc(output_unit_0_to_0_io_credit_alloc_2_alloc),
    .io_credit_alloc_3_alloc(output_unit_0_to_0_io_credit_alloc_3_alloc),
    .io_out_flit_0_valid(output_unit_0_to_0_io_out_flit_0_valid),
    .io_out_flit_0_bits_head(output_unit_0_to_0_io_out_flit_0_bits_head),
    .io_out_flit_0_bits_tail(output_unit_0_to_0_io_out_flit_0_bits_tail),
    .io_out_flit_0_bits_payload(output_unit_0_to_0_io_out_flit_0_bits_payload),
    .io_out_flit_0_bits_flow_ingress_node(output_unit_0_to_0_io_out_flit_0_bits_flow_ingress_node),
    .io_out_flit_0_bits_flow_egress_node(output_unit_0_to_0_io_out_flit_0_bits_flow_egress_node),
    .io_out_flit_0_bits_virt_channel_id(output_unit_0_to_0_io_out_flit_0_bits_virt_channel_id),
    .io_out_credit_return(output_unit_0_to_0_io_out_credit_return),
    .io_out_vc_free(output_unit_0_to_0_io_out_vc_free)
  );
  OutputUnit output_unit_1_to_2 ( // @[Router.scala 122:13]
    .clock(output_unit_1_to_2_clock),
    .reset(output_unit_1_to_2_reset),
    .io_in_0_valid(output_unit_1_to_2_io_in_0_valid),
    .io_in_0_bits_head(output_unit_1_to_2_io_in_0_bits_head),
    .io_in_0_bits_tail(output_unit_1_to_2_io_in_0_bits_tail),
    .io_in_0_bits_payload(output_unit_1_to_2_io_in_0_bits_payload),
    .io_in_0_bits_flow_ingress_node(output_unit_1_to_2_io_in_0_bits_flow_ingress_node),
    .io_in_0_bits_flow_egress_node(output_unit_1_to_2_io_in_0_bits_flow_egress_node),
    .io_in_0_bits_virt_channel_id(output_unit_1_to_2_io_in_0_bits_virt_channel_id),
    .io_credit_available_0(output_unit_1_to_2_io_credit_available_0),
    .io_credit_available_1(output_unit_1_to_2_io_credit_available_1),
    .io_credit_available_2(output_unit_1_to_2_io_credit_available_2),
    .io_credit_available_3(output_unit_1_to_2_io_credit_available_3),
    .io_channel_status_0_occupied(output_unit_1_to_2_io_channel_status_0_occupied),
    .io_channel_status_1_occupied(output_unit_1_to_2_io_channel_status_1_occupied),
    .io_channel_status_2_occupied(output_unit_1_to_2_io_channel_status_2_occupied),
    .io_channel_status_3_occupied(output_unit_1_to_2_io_channel_status_3_occupied),
    .io_allocs_0_alloc(output_unit_1_to_2_io_allocs_0_alloc),
    .io_allocs_1_alloc(output_unit_1_to_2_io_allocs_1_alloc),
    .io_allocs_2_alloc(output_unit_1_to_2_io_allocs_2_alloc),
    .io_allocs_3_alloc(output_unit_1_to_2_io_allocs_3_alloc),
    .io_credit_alloc_0_alloc(output_unit_1_to_2_io_credit_alloc_0_alloc),
    .io_credit_alloc_1_alloc(output_unit_1_to_2_io_credit_alloc_1_alloc),
    .io_credit_alloc_2_alloc(output_unit_1_to_2_io_credit_alloc_2_alloc),
    .io_credit_alloc_3_alloc(output_unit_1_to_2_io_credit_alloc_3_alloc),
    .io_out_flit_0_valid(output_unit_1_to_2_io_out_flit_0_valid),
    .io_out_flit_0_bits_head(output_unit_1_to_2_io_out_flit_0_bits_head),
    .io_out_flit_0_bits_tail(output_unit_1_to_2_io_out_flit_0_bits_tail),
    .io_out_flit_0_bits_payload(output_unit_1_to_2_io_out_flit_0_bits_payload),
    .io_out_flit_0_bits_flow_ingress_node(output_unit_1_to_2_io_out_flit_0_bits_flow_ingress_node),
    .io_out_flit_0_bits_flow_egress_node(output_unit_1_to_2_io_out_flit_0_bits_flow_egress_node),
    .io_out_flit_0_bits_virt_channel_id(output_unit_1_to_2_io_out_flit_0_bits_virt_channel_id),
    .io_out_credit_return(output_unit_1_to_2_io_out_credit_return),
    .io_out_vc_free(output_unit_1_to_2_io_out_vc_free)
  );
  EgressUnit egress_unit_2_to_3 ( // @[Router.scala 125:13]
    .clock(egress_unit_2_to_3_clock),
    .reset(egress_unit_2_to_3_reset),
    .io_in_0_valid(egress_unit_2_to_3_io_in_0_valid),
    .io_in_0_bits_head(egress_unit_2_to_3_io_in_0_bits_head),
    .io_in_0_bits_tail(egress_unit_2_to_3_io_in_0_bits_tail),
    .io_in_0_bits_payload(egress_unit_2_to_3_io_in_0_bits_payload),
    .io_in_0_bits_flow_ingress_node(egress_unit_2_to_3_io_in_0_bits_flow_ingress_node),
    .io_credit_available_0(egress_unit_2_to_3_io_credit_available_0),
    .io_channel_status_0_occupied(egress_unit_2_to_3_io_channel_status_0_occupied),
    .io_allocs_0_alloc(egress_unit_2_to_3_io_allocs_0_alloc),
    .io_credit_alloc_0_alloc(egress_unit_2_to_3_io_credit_alloc_0_alloc),
    .io_credit_alloc_0_tail(egress_unit_2_to_3_io_credit_alloc_0_tail),
    .io_out_valid(egress_unit_2_to_3_io_out_valid),
    .io_out_bits_head(egress_unit_2_to_3_io_out_bits_head),
    .io_out_bits_tail(egress_unit_2_to_3_io_out_bits_tail),
    .io_out_bits_payload(egress_unit_2_to_3_io_out_bits_payload),
    .io_out_bits_ingress_id(egress_unit_2_to_3_io_out_bits_ingress_id)
  );
  Switch switch ( // @[Router.scala 129:24]
    .clock(switch_clock),
    .reset(switch_reset),
    .io_in_2_0_valid(switch_io_in_2_0_valid),
    .io_in_2_0_bits_flit_head(switch_io_in_2_0_bits_flit_head),
    .io_in_2_0_bits_flit_tail(switch_io_in_2_0_bits_flit_tail),
    .io_in_2_0_bits_flit_payload(switch_io_in_2_0_bits_flit_payload),
    .io_in_2_0_bits_flit_flow_ingress_node(switch_io_in_2_0_bits_flit_flow_ingress_node),
    .io_in_2_0_bits_flit_flow_egress_node(switch_io_in_2_0_bits_flit_flow_egress_node),
    .io_in_2_0_bits_out_virt_channel(switch_io_in_2_0_bits_out_virt_channel),
    .io_in_1_0_valid(switch_io_in_1_0_valid),
    .io_in_1_0_bits_flit_head(switch_io_in_1_0_bits_flit_head),
    .io_in_1_0_bits_flit_tail(switch_io_in_1_0_bits_flit_tail),
    .io_in_1_0_bits_flit_payload(switch_io_in_1_0_bits_flit_payload),
    .io_in_1_0_bits_flit_flow_ingress_node(switch_io_in_1_0_bits_flit_flow_ingress_node),
    .io_in_1_0_bits_flit_flow_egress_node(switch_io_in_1_0_bits_flit_flow_egress_node),
    .io_in_1_0_bits_out_virt_channel(switch_io_in_1_0_bits_out_virt_channel),
    .io_in_0_0_valid(switch_io_in_0_0_valid),
    .io_in_0_0_bits_flit_head(switch_io_in_0_0_bits_flit_head),
    .io_in_0_0_bits_flit_tail(switch_io_in_0_0_bits_flit_tail),
    .io_in_0_0_bits_flit_payload(switch_io_in_0_0_bits_flit_payload),
    .io_in_0_0_bits_flit_flow_ingress_node(switch_io_in_0_0_bits_flit_flow_ingress_node),
    .io_in_0_0_bits_flit_flow_egress_node(switch_io_in_0_0_bits_flit_flow_egress_node),
    .io_in_0_0_bits_out_virt_channel(switch_io_in_0_0_bits_out_virt_channel),
    .io_out_2_0_valid(switch_io_out_2_0_valid),
    .io_out_2_0_bits_head(switch_io_out_2_0_bits_head),
    .io_out_2_0_bits_tail(switch_io_out_2_0_bits_tail),
    .io_out_2_0_bits_payload(switch_io_out_2_0_bits_payload),
    .io_out_2_0_bits_flow_ingress_node(switch_io_out_2_0_bits_flow_ingress_node),
    .io_out_1_0_valid(switch_io_out_1_0_valid),
    .io_out_1_0_bits_head(switch_io_out_1_0_bits_head),
    .io_out_1_0_bits_tail(switch_io_out_1_0_bits_tail),
    .io_out_1_0_bits_payload(switch_io_out_1_0_bits_payload),
    .io_out_1_0_bits_flow_ingress_node(switch_io_out_1_0_bits_flow_ingress_node),
    .io_out_1_0_bits_flow_egress_node(switch_io_out_1_0_bits_flow_egress_node),
    .io_out_1_0_bits_virt_channel_id(switch_io_out_1_0_bits_virt_channel_id),
    .io_out_0_0_valid(switch_io_out_0_0_valid),
    .io_out_0_0_bits_head(switch_io_out_0_0_bits_head),
    .io_out_0_0_bits_tail(switch_io_out_0_0_bits_tail),
    .io_out_0_0_bits_payload(switch_io_out_0_0_bits_payload),
    .io_out_0_0_bits_flow_ingress_node(switch_io_out_0_0_bits_flow_ingress_node),
    .io_out_0_0_bits_flow_egress_node(switch_io_out_0_0_bits_flow_egress_node),
    .io_out_0_0_bits_virt_channel_id(switch_io_out_0_0_bits_virt_channel_id),
    .io_sel_2_0_2_0(switch_io_sel_2_0_2_0),
    .io_sel_2_0_1_0(switch_io_sel_2_0_1_0),
    .io_sel_2_0_0_0(switch_io_sel_2_0_0_0),
    .io_sel_1_0_2_0(switch_io_sel_1_0_2_0),
    .io_sel_1_0_1_0(switch_io_sel_1_0_1_0),
    .io_sel_1_0_0_0(switch_io_sel_1_0_0_0),
    .io_sel_0_0_2_0(switch_io_sel_0_0_2_0),
    .io_sel_0_0_1_0(switch_io_sel_0_0_1_0),
    .io_sel_0_0_0_0(switch_io_sel_0_0_0_0)
  );
  SwitchAllocator switch_allocator ( // @[Router.scala 130:34]
    .clock(switch_allocator_clock),
    .reset(switch_allocator_reset),
    .io_req_2_0_ready(switch_allocator_io_req_2_0_ready),
    .io_req_2_0_valid(switch_allocator_io_req_2_0_valid),
    .io_req_2_0_bits_vc_sel_2_0(switch_allocator_io_req_2_0_bits_vc_sel_2_0),
    .io_req_2_0_bits_vc_sel_1_0(switch_allocator_io_req_2_0_bits_vc_sel_1_0),
    .io_req_2_0_bits_vc_sel_1_1(switch_allocator_io_req_2_0_bits_vc_sel_1_1),
    .io_req_2_0_bits_vc_sel_1_2(switch_allocator_io_req_2_0_bits_vc_sel_1_2),
    .io_req_2_0_bits_vc_sel_1_3(switch_allocator_io_req_2_0_bits_vc_sel_1_3),
    .io_req_2_0_bits_vc_sel_0_0(switch_allocator_io_req_2_0_bits_vc_sel_0_0),
    .io_req_2_0_bits_vc_sel_0_1(switch_allocator_io_req_2_0_bits_vc_sel_0_1),
    .io_req_2_0_bits_vc_sel_0_2(switch_allocator_io_req_2_0_bits_vc_sel_0_2),
    .io_req_2_0_bits_vc_sel_0_3(switch_allocator_io_req_2_0_bits_vc_sel_0_3),
    .io_req_2_0_bits_tail(switch_allocator_io_req_2_0_bits_tail),
    .io_req_1_0_ready(switch_allocator_io_req_1_0_ready),
    .io_req_1_0_valid(switch_allocator_io_req_1_0_valid),
    .io_req_1_0_bits_vc_sel_2_0(switch_allocator_io_req_1_0_bits_vc_sel_2_0),
    .io_req_1_0_bits_vc_sel_1_0(switch_allocator_io_req_1_0_bits_vc_sel_1_0),
    .io_req_1_0_bits_vc_sel_1_1(switch_allocator_io_req_1_0_bits_vc_sel_1_1),
    .io_req_1_0_bits_vc_sel_1_2(switch_allocator_io_req_1_0_bits_vc_sel_1_2),
    .io_req_1_0_bits_vc_sel_1_3(switch_allocator_io_req_1_0_bits_vc_sel_1_3),
    .io_req_1_0_bits_vc_sel_0_0(switch_allocator_io_req_1_0_bits_vc_sel_0_0),
    .io_req_1_0_bits_vc_sel_0_1(switch_allocator_io_req_1_0_bits_vc_sel_0_1),
    .io_req_1_0_bits_vc_sel_0_2(switch_allocator_io_req_1_0_bits_vc_sel_0_2),
    .io_req_1_0_bits_vc_sel_0_3(switch_allocator_io_req_1_0_bits_vc_sel_0_3),
    .io_req_1_0_bits_tail(switch_allocator_io_req_1_0_bits_tail),
    .io_req_0_0_ready(switch_allocator_io_req_0_0_ready),
    .io_req_0_0_valid(switch_allocator_io_req_0_0_valid),
    .io_req_0_0_bits_vc_sel_2_0(switch_allocator_io_req_0_0_bits_vc_sel_2_0),
    .io_req_0_0_bits_vc_sel_1_0(switch_allocator_io_req_0_0_bits_vc_sel_1_0),
    .io_req_0_0_bits_vc_sel_1_1(switch_allocator_io_req_0_0_bits_vc_sel_1_1),
    .io_req_0_0_bits_vc_sel_1_2(switch_allocator_io_req_0_0_bits_vc_sel_1_2),
    .io_req_0_0_bits_vc_sel_1_3(switch_allocator_io_req_0_0_bits_vc_sel_1_3),
    .io_req_0_0_bits_vc_sel_0_0(switch_allocator_io_req_0_0_bits_vc_sel_0_0),
    .io_req_0_0_bits_vc_sel_0_1(switch_allocator_io_req_0_0_bits_vc_sel_0_1),
    .io_req_0_0_bits_vc_sel_0_2(switch_allocator_io_req_0_0_bits_vc_sel_0_2),
    .io_req_0_0_bits_vc_sel_0_3(switch_allocator_io_req_0_0_bits_vc_sel_0_3),
    .io_req_0_0_bits_tail(switch_allocator_io_req_0_0_bits_tail),
    .io_credit_alloc_2_0_alloc(switch_allocator_io_credit_alloc_2_0_alloc),
    .io_credit_alloc_2_0_tail(switch_allocator_io_credit_alloc_2_0_tail),
    .io_credit_alloc_1_0_alloc(switch_allocator_io_credit_alloc_1_0_alloc),
    .io_credit_alloc_1_1_alloc(switch_allocator_io_credit_alloc_1_1_alloc),
    .io_credit_alloc_1_2_alloc(switch_allocator_io_credit_alloc_1_2_alloc),
    .io_credit_alloc_1_3_alloc(switch_allocator_io_credit_alloc_1_3_alloc),
    .io_credit_alloc_0_0_alloc(switch_allocator_io_credit_alloc_0_0_alloc),
    .io_credit_alloc_0_1_alloc(switch_allocator_io_credit_alloc_0_1_alloc),
    .io_credit_alloc_0_2_alloc(switch_allocator_io_credit_alloc_0_2_alloc),
    .io_credit_alloc_0_3_alloc(switch_allocator_io_credit_alloc_0_3_alloc),
    .io_switch_sel_2_0_2_0(switch_allocator_io_switch_sel_2_0_2_0),
    .io_switch_sel_2_0_1_0(switch_allocator_io_switch_sel_2_0_1_0),
    .io_switch_sel_2_0_0_0(switch_allocator_io_switch_sel_2_0_0_0),
    .io_switch_sel_1_0_2_0(switch_allocator_io_switch_sel_1_0_2_0),
    .io_switch_sel_1_0_1_0(switch_allocator_io_switch_sel_1_0_1_0),
    .io_switch_sel_1_0_0_0(switch_allocator_io_switch_sel_1_0_0_0),
    .io_switch_sel_0_0_2_0(switch_allocator_io_switch_sel_0_0_2_0),
    .io_switch_sel_0_0_1_0(switch_allocator_io_switch_sel_0_0_1_0),
    .io_switch_sel_0_0_0_0(switch_allocator_io_switch_sel_0_0_0_0)
  );
  RotatingSingleVCAllocator vc_allocator ( // @[Router.scala 131:30]
    .clock(vc_allocator_clock),
    .reset(vc_allocator_reset),
    .io_req_2_ready(vc_allocator_io_req_2_ready),
    .io_req_2_valid(vc_allocator_io_req_2_valid),
    .io_req_2_bits_vc_sel_2_0(vc_allocator_io_req_2_bits_vc_sel_2_0),
    .io_req_2_bits_vc_sel_1_0(vc_allocator_io_req_2_bits_vc_sel_1_0),
    .io_req_2_bits_vc_sel_1_1(vc_allocator_io_req_2_bits_vc_sel_1_1),
    .io_req_2_bits_vc_sel_1_2(vc_allocator_io_req_2_bits_vc_sel_1_2),
    .io_req_2_bits_vc_sel_1_3(vc_allocator_io_req_2_bits_vc_sel_1_3),
    .io_req_2_bits_vc_sel_0_0(vc_allocator_io_req_2_bits_vc_sel_0_0),
    .io_req_2_bits_vc_sel_0_1(vc_allocator_io_req_2_bits_vc_sel_0_1),
    .io_req_2_bits_vc_sel_0_2(vc_allocator_io_req_2_bits_vc_sel_0_2),
    .io_req_2_bits_vc_sel_0_3(vc_allocator_io_req_2_bits_vc_sel_0_3),
    .io_req_1_ready(vc_allocator_io_req_1_ready),
    .io_req_1_valid(vc_allocator_io_req_1_valid),
    .io_req_1_bits_vc_sel_2_0(vc_allocator_io_req_1_bits_vc_sel_2_0),
    .io_req_1_bits_vc_sel_1_0(vc_allocator_io_req_1_bits_vc_sel_1_0),
    .io_req_1_bits_vc_sel_1_1(vc_allocator_io_req_1_bits_vc_sel_1_1),
    .io_req_1_bits_vc_sel_1_2(vc_allocator_io_req_1_bits_vc_sel_1_2),
    .io_req_1_bits_vc_sel_1_3(vc_allocator_io_req_1_bits_vc_sel_1_3),
    .io_req_1_bits_vc_sel_0_0(vc_allocator_io_req_1_bits_vc_sel_0_0),
    .io_req_1_bits_vc_sel_0_1(vc_allocator_io_req_1_bits_vc_sel_0_1),
    .io_req_1_bits_vc_sel_0_2(vc_allocator_io_req_1_bits_vc_sel_0_2),
    .io_req_1_bits_vc_sel_0_3(vc_allocator_io_req_1_bits_vc_sel_0_3),
    .io_req_0_ready(vc_allocator_io_req_0_ready),
    .io_req_0_valid(vc_allocator_io_req_0_valid),
    .io_req_0_bits_vc_sel_2_0(vc_allocator_io_req_0_bits_vc_sel_2_0),
    .io_req_0_bits_vc_sel_1_0(vc_allocator_io_req_0_bits_vc_sel_1_0),
    .io_req_0_bits_vc_sel_1_1(vc_allocator_io_req_0_bits_vc_sel_1_1),
    .io_req_0_bits_vc_sel_1_2(vc_allocator_io_req_0_bits_vc_sel_1_2),
    .io_req_0_bits_vc_sel_1_3(vc_allocator_io_req_0_bits_vc_sel_1_3),
    .io_req_0_bits_vc_sel_0_0(vc_allocator_io_req_0_bits_vc_sel_0_0),
    .io_req_0_bits_vc_sel_0_1(vc_allocator_io_req_0_bits_vc_sel_0_1),
    .io_req_0_bits_vc_sel_0_2(vc_allocator_io_req_0_bits_vc_sel_0_2),
    .io_req_0_bits_vc_sel_0_3(vc_allocator_io_req_0_bits_vc_sel_0_3),
    .io_resp_2_vc_sel_2_0(vc_allocator_io_resp_2_vc_sel_2_0),
    .io_resp_2_vc_sel_1_0(vc_allocator_io_resp_2_vc_sel_1_0),
    .io_resp_2_vc_sel_1_1(vc_allocator_io_resp_2_vc_sel_1_1),
    .io_resp_2_vc_sel_1_2(vc_allocator_io_resp_2_vc_sel_1_2),
    .io_resp_2_vc_sel_1_3(vc_allocator_io_resp_2_vc_sel_1_3),
    .io_resp_2_vc_sel_0_0(vc_allocator_io_resp_2_vc_sel_0_0),
    .io_resp_2_vc_sel_0_1(vc_allocator_io_resp_2_vc_sel_0_1),
    .io_resp_2_vc_sel_0_2(vc_allocator_io_resp_2_vc_sel_0_2),
    .io_resp_2_vc_sel_0_3(vc_allocator_io_resp_2_vc_sel_0_3),
    .io_resp_1_vc_sel_2_0(vc_allocator_io_resp_1_vc_sel_2_0),
    .io_resp_1_vc_sel_1_0(vc_allocator_io_resp_1_vc_sel_1_0),
    .io_resp_1_vc_sel_1_1(vc_allocator_io_resp_1_vc_sel_1_1),
    .io_resp_1_vc_sel_1_2(vc_allocator_io_resp_1_vc_sel_1_2),
    .io_resp_1_vc_sel_1_3(vc_allocator_io_resp_1_vc_sel_1_3),
    .io_resp_1_vc_sel_0_0(vc_allocator_io_resp_1_vc_sel_0_0),
    .io_resp_1_vc_sel_0_1(vc_allocator_io_resp_1_vc_sel_0_1),
    .io_resp_1_vc_sel_0_2(vc_allocator_io_resp_1_vc_sel_0_2),
    .io_resp_1_vc_sel_0_3(vc_allocator_io_resp_1_vc_sel_0_3),
    .io_resp_0_vc_sel_2_0(vc_allocator_io_resp_0_vc_sel_2_0),
    .io_resp_0_vc_sel_1_0(vc_allocator_io_resp_0_vc_sel_1_0),
    .io_resp_0_vc_sel_1_1(vc_allocator_io_resp_0_vc_sel_1_1),
    .io_resp_0_vc_sel_1_2(vc_allocator_io_resp_0_vc_sel_1_2),
    .io_resp_0_vc_sel_1_3(vc_allocator_io_resp_0_vc_sel_1_3),
    .io_resp_0_vc_sel_0_0(vc_allocator_io_resp_0_vc_sel_0_0),
    .io_resp_0_vc_sel_0_1(vc_allocator_io_resp_0_vc_sel_0_1),
    .io_resp_0_vc_sel_0_2(vc_allocator_io_resp_0_vc_sel_0_2),
    .io_resp_0_vc_sel_0_3(vc_allocator_io_resp_0_vc_sel_0_3),
    .io_channel_status_2_0_occupied(vc_allocator_io_channel_status_2_0_occupied),
    .io_channel_status_1_0_occupied(vc_allocator_io_channel_status_1_0_occupied),
    .io_channel_status_1_1_occupied(vc_allocator_io_channel_status_1_1_occupied),
    .io_channel_status_1_2_occupied(vc_allocator_io_channel_status_1_2_occupied),
    .io_channel_status_1_3_occupied(vc_allocator_io_channel_status_1_3_occupied),
    .io_channel_status_0_0_occupied(vc_allocator_io_channel_status_0_0_occupied),
    .io_channel_status_0_1_occupied(vc_allocator_io_channel_status_0_1_occupied),
    .io_channel_status_0_2_occupied(vc_allocator_io_channel_status_0_2_occupied),
    .io_channel_status_0_3_occupied(vc_allocator_io_channel_status_0_3_occupied),
    .io_out_allocs_2_0_alloc(vc_allocator_io_out_allocs_2_0_alloc),
    .io_out_allocs_1_0_alloc(vc_allocator_io_out_allocs_1_0_alloc),
    .io_out_allocs_1_1_alloc(vc_allocator_io_out_allocs_1_1_alloc),
    .io_out_allocs_1_2_alloc(vc_allocator_io_out_allocs_1_2_alloc),
    .io_out_allocs_1_3_alloc(vc_allocator_io_out_allocs_1_3_alloc),
    .io_out_allocs_0_0_alloc(vc_allocator_io_out_allocs_0_0_alloc),
    .io_out_allocs_0_1_alloc(vc_allocator_io_out_allocs_0_1_alloc),
    .io_out_allocs_0_2_alloc(vc_allocator_io_out_allocs_0_2_alloc),
    .io_out_allocs_0_3_alloc(vc_allocator_io_out_allocs_0_3_alloc)
  );
  RouteComputer_3 route_computer ( // @[Router.scala 134:32]
    .io_req_2_bits_flow_ingress_node(route_computer_io_req_2_bits_flow_ingress_node),
    .io_req_2_bits_flow_egress_node(route_computer_io_req_2_bits_flow_egress_node),
    .io_req_1_bits_src_virt_id(route_computer_io_req_1_bits_src_virt_id),
    .io_req_1_bits_flow_ingress_node(route_computer_io_req_1_bits_flow_ingress_node),
    .io_req_1_bits_flow_egress_node(route_computer_io_req_1_bits_flow_egress_node),
    .io_req_0_bits_src_virt_id(route_computer_io_req_0_bits_src_virt_id),
    .io_req_0_bits_flow_ingress_node(route_computer_io_req_0_bits_flow_ingress_node),
    .io_req_0_bits_flow_egress_node(route_computer_io_req_0_bits_flow_egress_node),
    .io_resp_2_vc_sel_1_0(route_computer_io_resp_2_vc_sel_1_0),
    .io_resp_2_vc_sel_1_1(route_computer_io_resp_2_vc_sel_1_1),
    .io_resp_2_vc_sel_1_2(route_computer_io_resp_2_vc_sel_1_2),
    .io_resp_2_vc_sel_1_3(route_computer_io_resp_2_vc_sel_1_3),
    .io_resp_2_vc_sel_0_0(route_computer_io_resp_2_vc_sel_0_0),
    .io_resp_2_vc_sel_0_1(route_computer_io_resp_2_vc_sel_0_1),
    .io_resp_2_vc_sel_0_2(route_computer_io_resp_2_vc_sel_0_2),
    .io_resp_2_vc_sel_0_3(route_computer_io_resp_2_vc_sel_0_3),
    .io_resp_1_vc_sel_1_0(route_computer_io_resp_1_vc_sel_1_0),
    .io_resp_1_vc_sel_1_1(route_computer_io_resp_1_vc_sel_1_1),
    .io_resp_1_vc_sel_1_2(route_computer_io_resp_1_vc_sel_1_2),
    .io_resp_1_vc_sel_1_3(route_computer_io_resp_1_vc_sel_1_3),
    .io_resp_1_vc_sel_0_0(route_computer_io_resp_1_vc_sel_0_0),
    .io_resp_1_vc_sel_0_1(route_computer_io_resp_1_vc_sel_0_1),
    .io_resp_1_vc_sel_0_2(route_computer_io_resp_1_vc_sel_0_2),
    .io_resp_0_vc_sel_1_0(route_computer_io_resp_0_vc_sel_1_0),
    .io_resp_0_vc_sel_1_1(route_computer_io_resp_0_vc_sel_1_1),
    .io_resp_0_vc_sel_1_2(route_computer_io_resp_0_vc_sel_1_2),
    .io_resp_0_vc_sel_1_3(route_computer_io_resp_0_vc_sel_1_3),
    .io_resp_0_vc_sel_0_0(route_computer_io_resp_0_vc_sel_0_0),
    .io_resp_0_vc_sel_0_1(route_computer_io_resp_0_vc_sel_0_1),
    .io_resp_0_vc_sel_0_2(route_computer_io_resp_0_vc_sel_0_2)
  );
  plusarg_reader #(.FORMAT("noc_util_sample_rate=%d"), .DEFAULT(0), .WIDTH(20)) plusarg_reader ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_out)
  );
  assign auto_debug_out_va_stall_0 = input_unit_0_from_0_io_debug_va_stall; // @[Nodes.scala 1212:84 Router.scala 190:92]
  assign auto_debug_out_va_stall_1 = input_unit_1_from_2_io_debug_va_stall; // @[Nodes.scala 1212:84 Router.scala 190:92]
  assign auto_debug_out_sa_stall_0 = input_unit_0_from_0_io_debug_sa_stall; // @[Nodes.scala 1212:84 Router.scala 191:92]
  assign auto_debug_out_sa_stall_1 = input_unit_1_from_2_io_debug_sa_stall; // @[Nodes.scala 1212:84 Router.scala 191:92]
  assign auto_egress_nodes_out_flit_valid = egress_unit_2_to_3_io_out_valid; // @[Nodes.scala 1212:84 Router.scala 144:65]
  assign auto_egress_nodes_out_flit_bits_head = egress_unit_2_to_3_io_out_bits_head; // @[Nodes.scala 1212:84 Router.scala 144:65]
  assign auto_egress_nodes_out_flit_bits_tail = egress_unit_2_to_3_io_out_bits_tail; // @[Nodes.scala 1212:84 Router.scala 144:65]
  assign auto_egress_nodes_out_flit_bits_payload = egress_unit_2_to_3_io_out_bits_payload; // @[Nodes.scala 1212:84 Router.scala 144:65]
  assign auto_egress_nodes_out_flit_bits_ingress_id = egress_unit_2_to_3_io_out_bits_ingress_id; // @[Nodes.scala 1212:84 Router.scala 144:65]
  assign auto_ingress_nodes_in_flit_ready = ingress_unit_2_from_3_io_in_ready; // @[Nodes.scala 1215:84 Router.scala 142:68]
  assign auto_source_nodes_out_1_flit_0_valid = output_unit_1_to_2_io_out_flit_0_valid; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_1_flit_0_bits_head = output_unit_1_to_2_io_out_flit_0_bits_head; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_1_flit_0_bits_tail = output_unit_1_to_2_io_out_flit_0_bits_tail; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_1_flit_0_bits_payload = output_unit_1_to_2_io_out_flit_0_bits_payload; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_1_flit_0_bits_flow_ingress_node = output_unit_1_to_2_io_out_flit_0_bits_flow_ingress_node
    ; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_1_flit_0_bits_flow_egress_node = output_unit_1_to_2_io_out_flit_0_bits_flow_egress_node; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_1_flit_0_bits_virt_channel_id = output_unit_1_to_2_io_out_flit_0_bits_virt_channel_id; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_0_flit_0_valid = output_unit_0_to_0_io_out_flit_0_valid; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_0_flit_0_bits_head = output_unit_0_to_0_io_out_flit_0_bits_head; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_0_flit_0_bits_tail = output_unit_0_to_0_io_out_flit_0_bits_tail; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_0_flit_0_bits_payload = output_unit_0_to_0_io_out_flit_0_bits_payload; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_0_flit_0_bits_flow_ingress_node = output_unit_0_to_0_io_out_flit_0_bits_flow_ingress_node
    ; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_0_flit_0_bits_flow_egress_node = output_unit_0_to_0_io_out_flit_0_bits_flow_egress_node; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_0_flit_0_bits_virt_channel_id = output_unit_0_to_0_io_out_flit_0_bits_virt_channel_id; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_dest_nodes_in_1_credit_return = input_unit_1_from_2_io_in_credit_return; // @[Nodes.scala 1215:84 Router.scala 141:68]
  assign auto_dest_nodes_in_1_vc_free = input_unit_1_from_2_io_in_vc_free; // @[Nodes.scala 1215:84 Router.scala 141:68]
  assign auto_dest_nodes_in_0_credit_return = input_unit_0_from_0_io_in_credit_return; // @[Nodes.scala 1215:84 Router.scala 141:68]
  assign auto_dest_nodes_in_0_vc_free = input_unit_0_from_0_io_in_vc_free; // @[Nodes.scala 1215:84 Router.scala 141:68]
  assign monitor_clock = clock;
  assign monitor_reset = reset;
  assign monitor_io_in_flit_0_valid = auto_dest_nodes_in_0_flit_0_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_io_in_flit_0_bits_head = auto_dest_nodes_in_0_flit_0_bits_head; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_io_in_flit_0_bits_tail = auto_dest_nodes_in_0_flit_0_bits_tail; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_io_in_flit_0_bits_flow_ingress_node = auto_dest_nodes_in_0_flit_0_bits_flow_ingress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_io_in_flit_0_bits_flow_egress_node = auto_dest_nodes_in_0_flit_0_bits_flow_egress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_io_in_flit_0_bits_virt_channel_id = auto_dest_nodes_in_0_flit_0_bits_virt_channel_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_1_clock = clock;
  assign monitor_1_reset = reset;
  assign monitor_1_io_in_flit_0_valid = auto_dest_nodes_in_1_flit_0_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_1_io_in_flit_0_bits_head = auto_dest_nodes_in_1_flit_0_bits_head; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_1_io_in_flit_0_bits_tail = auto_dest_nodes_in_1_flit_0_bits_tail; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_1_io_in_flit_0_bits_flow_ingress_node = auto_dest_nodes_in_1_flit_0_bits_flow_ingress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_1_io_in_flit_0_bits_flow_egress_node = auto_dest_nodes_in_1_flit_0_bits_flow_egress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_1_io_in_flit_0_bits_virt_channel_id = auto_dest_nodes_in_1_flit_0_bits_virt_channel_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_0_clock = clock;
  assign input_unit_0_from_0_reset = reset;
  assign input_unit_0_from_0_io_router_resp_vc_sel_1_0 = route_computer_io_resp_0_vc_sel_1_0; // @[Router.scala 148:38]
  assign input_unit_0_from_0_io_router_resp_vc_sel_1_1 = route_computer_io_resp_0_vc_sel_1_1; // @[Router.scala 148:38]
  assign input_unit_0_from_0_io_router_resp_vc_sel_1_2 = route_computer_io_resp_0_vc_sel_1_2; // @[Router.scala 148:38]
  assign input_unit_0_from_0_io_router_resp_vc_sel_1_3 = route_computer_io_resp_0_vc_sel_1_3; // @[Router.scala 148:38]
  assign input_unit_0_from_0_io_router_resp_vc_sel_0_0 = route_computer_io_resp_0_vc_sel_0_0; // @[Router.scala 148:38]
  assign input_unit_0_from_0_io_router_resp_vc_sel_0_1 = route_computer_io_resp_0_vc_sel_0_1; // @[Router.scala 148:38]
  assign input_unit_0_from_0_io_router_resp_vc_sel_0_2 = route_computer_io_resp_0_vc_sel_0_2; // @[Router.scala 148:38]
  assign input_unit_0_from_0_io_vcalloc_req_ready = vc_allocator_io_req_0_ready; // @[Router.scala 151:23]
  assign input_unit_0_from_0_io_vcalloc_resp_vc_sel_2_0 = vc_allocator_io_resp_0_vc_sel_2_0; // @[Router.scala 153:39]
  assign input_unit_0_from_0_io_vcalloc_resp_vc_sel_1_0 = vc_allocator_io_resp_0_vc_sel_1_0; // @[Router.scala 153:39]
  assign input_unit_0_from_0_io_vcalloc_resp_vc_sel_1_1 = vc_allocator_io_resp_0_vc_sel_1_1; // @[Router.scala 153:39]
  assign input_unit_0_from_0_io_vcalloc_resp_vc_sel_1_2 = vc_allocator_io_resp_0_vc_sel_1_2; // @[Router.scala 153:39]
  assign input_unit_0_from_0_io_vcalloc_resp_vc_sel_1_3 = vc_allocator_io_resp_0_vc_sel_1_3; // @[Router.scala 153:39]
  assign input_unit_0_from_0_io_vcalloc_resp_vc_sel_0_0 = vc_allocator_io_resp_0_vc_sel_0_0; // @[Router.scala 153:39]
  assign input_unit_0_from_0_io_vcalloc_resp_vc_sel_0_1 = vc_allocator_io_resp_0_vc_sel_0_1; // @[Router.scala 153:39]
  assign input_unit_0_from_0_io_vcalloc_resp_vc_sel_0_2 = vc_allocator_io_resp_0_vc_sel_0_2; // @[Router.scala 153:39]
  assign input_unit_0_from_0_io_out_credit_available_2_0 = egress_unit_2_to_3_io_credit_available_0; // @[Router.scala 162:42]
  assign input_unit_0_from_0_io_out_credit_available_1_0 = output_unit_1_to_2_io_credit_available_0; // @[Router.scala 162:42]
  assign input_unit_0_from_0_io_out_credit_available_1_1 = output_unit_1_to_2_io_credit_available_1; // @[Router.scala 162:42]
  assign input_unit_0_from_0_io_out_credit_available_1_2 = output_unit_1_to_2_io_credit_available_2; // @[Router.scala 162:42]
  assign input_unit_0_from_0_io_out_credit_available_1_3 = output_unit_1_to_2_io_credit_available_3; // @[Router.scala 162:42]
  assign input_unit_0_from_0_io_out_credit_available_0_0 = output_unit_0_to_0_io_credit_available_0; // @[Router.scala 162:42]
  assign input_unit_0_from_0_io_out_credit_available_0_1 = output_unit_0_to_0_io_credit_available_1; // @[Router.scala 162:42]
  assign input_unit_0_from_0_io_out_credit_available_0_2 = output_unit_0_to_0_io_credit_available_2; // @[Router.scala 162:42]
  assign input_unit_0_from_0_io_out_credit_available_0_3 = output_unit_0_to_0_io_credit_available_3; // @[Router.scala 162:42]
  assign input_unit_0_from_0_io_salloc_req_0_ready = switch_allocator_io_req_0_0_ready; // @[Router.scala 165:23]
  assign input_unit_0_from_0_io_in_flit_0_valid = auto_dest_nodes_in_0_flit_0_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_0_io_in_flit_0_bits_head = auto_dest_nodes_in_0_flit_0_bits_head; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_0_io_in_flit_0_bits_tail = auto_dest_nodes_in_0_flit_0_bits_tail; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_0_io_in_flit_0_bits_payload = auto_dest_nodes_in_0_flit_0_bits_payload; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_0_io_in_flit_0_bits_flow_ingress_node = auto_dest_nodes_in_0_flit_0_bits_flow_ingress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_0_io_in_flit_0_bits_flow_egress_node = auto_dest_nodes_in_0_flit_0_bits_flow_egress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_0_io_in_flit_0_bits_virt_channel_id = auto_dest_nodes_in_0_flit_0_bits_virt_channel_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_1_from_2_clock = clock;
  assign input_unit_1_from_2_reset = reset;
  assign input_unit_1_from_2_io_router_resp_vc_sel_1_0 = route_computer_io_resp_1_vc_sel_1_0; // @[Router.scala 148:38]
  assign input_unit_1_from_2_io_router_resp_vc_sel_1_1 = route_computer_io_resp_1_vc_sel_1_1; // @[Router.scala 148:38]
  assign input_unit_1_from_2_io_router_resp_vc_sel_1_2 = route_computer_io_resp_1_vc_sel_1_2; // @[Router.scala 148:38]
  assign input_unit_1_from_2_io_router_resp_vc_sel_1_3 = route_computer_io_resp_1_vc_sel_1_3; // @[Router.scala 148:38]
  assign input_unit_1_from_2_io_router_resp_vc_sel_0_0 = route_computer_io_resp_1_vc_sel_0_0; // @[Router.scala 148:38]
  assign input_unit_1_from_2_io_router_resp_vc_sel_0_1 = route_computer_io_resp_1_vc_sel_0_1; // @[Router.scala 148:38]
  assign input_unit_1_from_2_io_router_resp_vc_sel_0_2 = route_computer_io_resp_1_vc_sel_0_2; // @[Router.scala 148:38]
  assign input_unit_1_from_2_io_vcalloc_req_ready = vc_allocator_io_req_1_ready; // @[Router.scala 151:23]
  assign input_unit_1_from_2_io_vcalloc_resp_vc_sel_2_0 = vc_allocator_io_resp_1_vc_sel_2_0; // @[Router.scala 153:39]
  assign input_unit_1_from_2_io_vcalloc_resp_vc_sel_1_0 = vc_allocator_io_resp_1_vc_sel_1_0; // @[Router.scala 153:39]
  assign input_unit_1_from_2_io_vcalloc_resp_vc_sel_1_1 = vc_allocator_io_resp_1_vc_sel_1_1; // @[Router.scala 153:39]
  assign input_unit_1_from_2_io_vcalloc_resp_vc_sel_1_2 = vc_allocator_io_resp_1_vc_sel_1_2; // @[Router.scala 153:39]
  assign input_unit_1_from_2_io_vcalloc_resp_vc_sel_1_3 = vc_allocator_io_resp_1_vc_sel_1_3; // @[Router.scala 153:39]
  assign input_unit_1_from_2_io_vcalloc_resp_vc_sel_0_0 = vc_allocator_io_resp_1_vc_sel_0_0; // @[Router.scala 153:39]
  assign input_unit_1_from_2_io_vcalloc_resp_vc_sel_0_1 = vc_allocator_io_resp_1_vc_sel_0_1; // @[Router.scala 153:39]
  assign input_unit_1_from_2_io_vcalloc_resp_vc_sel_0_2 = vc_allocator_io_resp_1_vc_sel_0_2; // @[Router.scala 153:39]
  assign input_unit_1_from_2_io_out_credit_available_2_0 = egress_unit_2_to_3_io_credit_available_0; // @[Router.scala 162:42]
  assign input_unit_1_from_2_io_out_credit_available_1_0 = output_unit_1_to_2_io_credit_available_0; // @[Router.scala 162:42]
  assign input_unit_1_from_2_io_out_credit_available_1_1 = output_unit_1_to_2_io_credit_available_1; // @[Router.scala 162:42]
  assign input_unit_1_from_2_io_out_credit_available_1_2 = output_unit_1_to_2_io_credit_available_2; // @[Router.scala 162:42]
  assign input_unit_1_from_2_io_out_credit_available_1_3 = output_unit_1_to_2_io_credit_available_3; // @[Router.scala 162:42]
  assign input_unit_1_from_2_io_out_credit_available_0_0 = output_unit_0_to_0_io_credit_available_0; // @[Router.scala 162:42]
  assign input_unit_1_from_2_io_out_credit_available_0_1 = output_unit_0_to_0_io_credit_available_1; // @[Router.scala 162:42]
  assign input_unit_1_from_2_io_out_credit_available_0_2 = output_unit_0_to_0_io_credit_available_2; // @[Router.scala 162:42]
  assign input_unit_1_from_2_io_out_credit_available_0_3 = output_unit_0_to_0_io_credit_available_3; // @[Router.scala 162:42]
  assign input_unit_1_from_2_io_salloc_req_0_ready = switch_allocator_io_req_1_0_ready; // @[Router.scala 165:23]
  assign input_unit_1_from_2_io_in_flit_0_valid = auto_dest_nodes_in_1_flit_0_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_1_from_2_io_in_flit_0_bits_head = auto_dest_nodes_in_1_flit_0_bits_head; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_1_from_2_io_in_flit_0_bits_tail = auto_dest_nodes_in_1_flit_0_bits_tail; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_1_from_2_io_in_flit_0_bits_payload = auto_dest_nodes_in_1_flit_0_bits_payload; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_1_from_2_io_in_flit_0_bits_flow_ingress_node = auto_dest_nodes_in_1_flit_0_bits_flow_ingress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_1_from_2_io_in_flit_0_bits_flow_egress_node = auto_dest_nodes_in_1_flit_0_bits_flow_egress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_1_from_2_io_in_flit_0_bits_virt_channel_id = auto_dest_nodes_in_1_flit_0_bits_virt_channel_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign ingress_unit_2_from_3_clock = clock;
  assign ingress_unit_2_from_3_reset = reset;
  assign ingress_unit_2_from_3_io_router_resp_vc_sel_1_0 = route_computer_io_resp_2_vc_sel_1_0; // @[Router.scala 148:38]
  assign ingress_unit_2_from_3_io_router_resp_vc_sel_1_1 = route_computer_io_resp_2_vc_sel_1_1; // @[Router.scala 148:38]
  assign ingress_unit_2_from_3_io_router_resp_vc_sel_1_2 = route_computer_io_resp_2_vc_sel_1_2; // @[Router.scala 148:38]
  assign ingress_unit_2_from_3_io_router_resp_vc_sel_1_3 = route_computer_io_resp_2_vc_sel_1_3; // @[Router.scala 148:38]
  assign ingress_unit_2_from_3_io_router_resp_vc_sel_0_0 = route_computer_io_resp_2_vc_sel_0_0; // @[Router.scala 148:38]
  assign ingress_unit_2_from_3_io_router_resp_vc_sel_0_1 = route_computer_io_resp_2_vc_sel_0_1; // @[Router.scala 148:38]
  assign ingress_unit_2_from_3_io_router_resp_vc_sel_0_2 = route_computer_io_resp_2_vc_sel_0_2; // @[Router.scala 148:38]
  assign ingress_unit_2_from_3_io_router_resp_vc_sel_0_3 = route_computer_io_resp_2_vc_sel_0_3; // @[Router.scala 148:38]
  assign ingress_unit_2_from_3_io_vcalloc_req_ready = vc_allocator_io_req_2_ready; // @[Router.scala 151:23]
  assign ingress_unit_2_from_3_io_vcalloc_resp_vc_sel_2_0 = vc_allocator_io_resp_2_vc_sel_2_0; // @[Router.scala 153:39]
  assign ingress_unit_2_from_3_io_vcalloc_resp_vc_sel_1_0 = vc_allocator_io_resp_2_vc_sel_1_0; // @[Router.scala 153:39]
  assign ingress_unit_2_from_3_io_vcalloc_resp_vc_sel_1_1 = vc_allocator_io_resp_2_vc_sel_1_1; // @[Router.scala 153:39]
  assign ingress_unit_2_from_3_io_vcalloc_resp_vc_sel_1_2 = vc_allocator_io_resp_2_vc_sel_1_2; // @[Router.scala 153:39]
  assign ingress_unit_2_from_3_io_vcalloc_resp_vc_sel_1_3 = vc_allocator_io_resp_2_vc_sel_1_3; // @[Router.scala 153:39]
  assign ingress_unit_2_from_3_io_vcalloc_resp_vc_sel_0_0 = vc_allocator_io_resp_2_vc_sel_0_0; // @[Router.scala 153:39]
  assign ingress_unit_2_from_3_io_vcalloc_resp_vc_sel_0_1 = vc_allocator_io_resp_2_vc_sel_0_1; // @[Router.scala 153:39]
  assign ingress_unit_2_from_3_io_vcalloc_resp_vc_sel_0_2 = vc_allocator_io_resp_2_vc_sel_0_2; // @[Router.scala 153:39]
  assign ingress_unit_2_from_3_io_vcalloc_resp_vc_sel_0_3 = vc_allocator_io_resp_2_vc_sel_0_3; // @[Router.scala 153:39]
  assign ingress_unit_2_from_3_io_out_credit_available_2_0 = egress_unit_2_to_3_io_credit_available_0; // @[Router.scala 162:42]
  assign ingress_unit_2_from_3_io_out_credit_available_1_0 = output_unit_1_to_2_io_credit_available_0; // @[Router.scala 162:42]
  assign ingress_unit_2_from_3_io_out_credit_available_1_1 = output_unit_1_to_2_io_credit_available_1; // @[Router.scala 162:42]
  assign ingress_unit_2_from_3_io_out_credit_available_1_2 = output_unit_1_to_2_io_credit_available_2; // @[Router.scala 162:42]
  assign ingress_unit_2_from_3_io_out_credit_available_1_3 = output_unit_1_to_2_io_credit_available_3; // @[Router.scala 162:42]
  assign ingress_unit_2_from_3_io_out_credit_available_0_0 = output_unit_0_to_0_io_credit_available_0; // @[Router.scala 162:42]
  assign ingress_unit_2_from_3_io_out_credit_available_0_1 = output_unit_0_to_0_io_credit_available_1; // @[Router.scala 162:42]
  assign ingress_unit_2_from_3_io_out_credit_available_0_2 = output_unit_0_to_0_io_credit_available_2; // @[Router.scala 162:42]
  assign ingress_unit_2_from_3_io_out_credit_available_0_3 = output_unit_0_to_0_io_credit_available_3; // @[Router.scala 162:42]
  assign ingress_unit_2_from_3_io_salloc_req_0_ready = switch_allocator_io_req_2_0_ready; // @[Router.scala 165:23]
  assign ingress_unit_2_from_3_io_in_valid = auto_ingress_nodes_in_flit_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign ingress_unit_2_from_3_io_in_bits_head = auto_ingress_nodes_in_flit_bits_head; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign ingress_unit_2_from_3_io_in_bits_tail = auto_ingress_nodes_in_flit_bits_tail; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign ingress_unit_2_from_3_io_in_bits_payload = auto_ingress_nodes_in_flit_bits_payload; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign ingress_unit_2_from_3_io_in_bits_egress_id = auto_ingress_nodes_in_flit_bits_egress_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign output_unit_0_to_0_clock = clock;
  assign output_unit_0_to_0_reset = reset;
  assign output_unit_0_to_0_io_in_0_valid = switch_io_out_0_0_valid; // @[Router.scala 172:29]
  assign output_unit_0_to_0_io_in_0_bits_head = switch_io_out_0_0_bits_head; // @[Router.scala 172:29]
  assign output_unit_0_to_0_io_in_0_bits_tail = switch_io_out_0_0_bits_tail; // @[Router.scala 172:29]
  assign output_unit_0_to_0_io_in_0_bits_payload = switch_io_out_0_0_bits_payload; // @[Router.scala 172:29]
  assign output_unit_0_to_0_io_in_0_bits_flow_ingress_node = switch_io_out_0_0_bits_flow_ingress_node; // @[Router.scala 172:29]
  assign output_unit_0_to_0_io_in_0_bits_flow_egress_node = switch_io_out_0_0_bits_flow_egress_node; // @[Router.scala 172:29]
  assign output_unit_0_to_0_io_in_0_bits_virt_channel_id = switch_io_out_0_0_bits_virt_channel_id; // @[Router.scala 172:29]
  assign output_unit_0_to_0_io_allocs_0_alloc = vc_allocator_io_out_allocs_0_0_alloc; // @[Router.scala 157:33]
  assign output_unit_0_to_0_io_allocs_1_alloc = vc_allocator_io_out_allocs_0_1_alloc; // @[Router.scala 157:33]
  assign output_unit_0_to_0_io_allocs_2_alloc = vc_allocator_io_out_allocs_0_2_alloc; // @[Router.scala 157:33]
  assign output_unit_0_to_0_io_allocs_3_alloc = vc_allocator_io_out_allocs_0_3_alloc; // @[Router.scala 157:33]
  assign output_unit_0_to_0_io_credit_alloc_0_alloc = switch_allocator_io_credit_alloc_0_0_alloc; // @[Router.scala 167:39]
  assign output_unit_0_to_0_io_credit_alloc_1_alloc = switch_allocator_io_credit_alloc_0_1_alloc; // @[Router.scala 167:39]
  assign output_unit_0_to_0_io_credit_alloc_2_alloc = switch_allocator_io_credit_alloc_0_2_alloc; // @[Router.scala 167:39]
  assign output_unit_0_to_0_io_credit_alloc_3_alloc = switch_allocator_io_credit_alloc_0_3_alloc; // @[Router.scala 167:39]
  assign output_unit_0_to_0_io_out_credit_return = auto_source_nodes_out_0_credit_return; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign output_unit_0_to_0_io_out_vc_free = auto_source_nodes_out_0_vc_free; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign output_unit_1_to_2_clock = clock;
  assign output_unit_1_to_2_reset = reset;
  assign output_unit_1_to_2_io_in_0_valid = switch_io_out_1_0_valid; // @[Router.scala 172:29]
  assign output_unit_1_to_2_io_in_0_bits_head = switch_io_out_1_0_bits_head; // @[Router.scala 172:29]
  assign output_unit_1_to_2_io_in_0_bits_tail = switch_io_out_1_0_bits_tail; // @[Router.scala 172:29]
  assign output_unit_1_to_2_io_in_0_bits_payload = switch_io_out_1_0_bits_payload; // @[Router.scala 172:29]
  assign output_unit_1_to_2_io_in_0_bits_flow_ingress_node = switch_io_out_1_0_bits_flow_ingress_node; // @[Router.scala 172:29]
  assign output_unit_1_to_2_io_in_0_bits_flow_egress_node = switch_io_out_1_0_bits_flow_egress_node; // @[Router.scala 172:29]
  assign output_unit_1_to_2_io_in_0_bits_virt_channel_id = switch_io_out_1_0_bits_virt_channel_id; // @[Router.scala 172:29]
  assign output_unit_1_to_2_io_allocs_0_alloc = vc_allocator_io_out_allocs_1_0_alloc; // @[Router.scala 157:33]
  assign output_unit_1_to_2_io_allocs_1_alloc = vc_allocator_io_out_allocs_1_1_alloc; // @[Router.scala 157:33]
  assign output_unit_1_to_2_io_allocs_2_alloc = vc_allocator_io_out_allocs_1_2_alloc; // @[Router.scala 157:33]
  assign output_unit_1_to_2_io_allocs_3_alloc = vc_allocator_io_out_allocs_1_3_alloc; // @[Router.scala 157:33]
  assign output_unit_1_to_2_io_credit_alloc_0_alloc = switch_allocator_io_credit_alloc_1_0_alloc; // @[Router.scala 167:39]
  assign output_unit_1_to_2_io_credit_alloc_1_alloc = switch_allocator_io_credit_alloc_1_1_alloc; // @[Router.scala 167:39]
  assign output_unit_1_to_2_io_credit_alloc_2_alloc = switch_allocator_io_credit_alloc_1_2_alloc; // @[Router.scala 167:39]
  assign output_unit_1_to_2_io_credit_alloc_3_alloc = switch_allocator_io_credit_alloc_1_3_alloc; // @[Router.scala 167:39]
  assign output_unit_1_to_2_io_out_credit_return = auto_source_nodes_out_1_credit_return; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign output_unit_1_to_2_io_out_vc_free = auto_source_nodes_out_1_vc_free; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign egress_unit_2_to_3_clock = clock;
  assign egress_unit_2_to_3_reset = reset;
  assign egress_unit_2_to_3_io_in_0_valid = switch_io_out_2_0_valid; // @[Router.scala 172:29]
  assign egress_unit_2_to_3_io_in_0_bits_head = switch_io_out_2_0_bits_head; // @[Router.scala 172:29]
  assign egress_unit_2_to_3_io_in_0_bits_tail = switch_io_out_2_0_bits_tail; // @[Router.scala 172:29]
  assign egress_unit_2_to_3_io_in_0_bits_payload = switch_io_out_2_0_bits_payload; // @[Router.scala 172:29]
  assign egress_unit_2_to_3_io_in_0_bits_flow_ingress_node = switch_io_out_2_0_bits_flow_ingress_node; // @[Router.scala 172:29]
  assign egress_unit_2_to_3_io_allocs_0_alloc = vc_allocator_io_out_allocs_2_0_alloc; // @[Router.scala 157:33]
  assign egress_unit_2_to_3_io_credit_alloc_0_alloc = switch_allocator_io_credit_alloc_2_0_alloc; // @[Router.scala 167:39]
  assign egress_unit_2_to_3_io_credit_alloc_0_tail = switch_allocator_io_credit_alloc_2_0_tail; // @[Router.scala 167:39]
  assign switch_clock = clock;
  assign switch_reset = reset;
  assign switch_io_in_2_0_valid = ingress_unit_2_from_3_io_out_0_valid; // @[Router.scala 170:23]
  assign switch_io_in_2_0_bits_flit_head = ingress_unit_2_from_3_io_out_0_bits_flit_head; // @[Router.scala 170:23]
  assign switch_io_in_2_0_bits_flit_tail = ingress_unit_2_from_3_io_out_0_bits_flit_tail; // @[Router.scala 170:23]
  assign switch_io_in_2_0_bits_flit_payload = ingress_unit_2_from_3_io_out_0_bits_flit_payload; // @[Router.scala 170:23]
  assign switch_io_in_2_0_bits_flit_flow_ingress_node = ingress_unit_2_from_3_io_out_0_bits_flit_flow_ingress_node; // @[Router.scala 170:23]
  assign switch_io_in_2_0_bits_flit_flow_egress_node = ingress_unit_2_from_3_io_out_0_bits_flit_flow_egress_node; // @[Router.scala 170:23]
  assign switch_io_in_2_0_bits_out_virt_channel = ingress_unit_2_from_3_io_out_0_bits_out_virt_channel; // @[Router.scala 170:23]
  assign switch_io_in_1_0_valid = input_unit_1_from_2_io_out_0_valid; // @[Router.scala 170:23]
  assign switch_io_in_1_0_bits_flit_head = input_unit_1_from_2_io_out_0_bits_flit_head; // @[Router.scala 170:23]
  assign switch_io_in_1_0_bits_flit_tail = input_unit_1_from_2_io_out_0_bits_flit_tail; // @[Router.scala 170:23]
  assign switch_io_in_1_0_bits_flit_payload = input_unit_1_from_2_io_out_0_bits_flit_payload; // @[Router.scala 170:23]
  assign switch_io_in_1_0_bits_flit_flow_ingress_node = input_unit_1_from_2_io_out_0_bits_flit_flow_ingress_node; // @[Router.scala 170:23]
  assign switch_io_in_1_0_bits_flit_flow_egress_node = input_unit_1_from_2_io_out_0_bits_flit_flow_egress_node; // @[Router.scala 170:23]
  assign switch_io_in_1_0_bits_out_virt_channel = input_unit_1_from_2_io_out_0_bits_out_virt_channel; // @[Router.scala 170:23]
  assign switch_io_in_0_0_valid = input_unit_0_from_0_io_out_0_valid; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_head = input_unit_0_from_0_io_out_0_bits_flit_head; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_tail = input_unit_0_from_0_io_out_0_bits_flit_tail; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_payload = input_unit_0_from_0_io_out_0_bits_flit_payload; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_flow_ingress_node = input_unit_0_from_0_io_out_0_bits_flit_flow_ingress_node; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_flow_egress_node = input_unit_0_from_0_io_out_0_bits_flit_flow_egress_node; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_out_virt_channel = input_unit_0_from_0_io_out_0_bits_out_virt_channel; // @[Router.scala 170:23]
  assign switch_io_sel_2_0_2_0 = switch_io_sel_REG_2_0_2_0; // @[Router.scala 173:19]
  assign switch_io_sel_2_0_1_0 = switch_io_sel_REG_2_0_1_0; // @[Router.scala 173:19]
  assign switch_io_sel_2_0_0_0 = switch_io_sel_REG_2_0_0_0; // @[Router.scala 173:19]
  assign switch_io_sel_1_0_2_0 = switch_io_sel_REG_1_0_2_0; // @[Router.scala 173:19]
  assign switch_io_sel_1_0_1_0 = switch_io_sel_REG_1_0_1_0; // @[Router.scala 173:19]
  assign switch_io_sel_1_0_0_0 = switch_io_sel_REG_1_0_0_0; // @[Router.scala 173:19]
  assign switch_io_sel_0_0_2_0 = switch_io_sel_REG_0_0_2_0; // @[Router.scala 173:19]
  assign switch_io_sel_0_0_1_0 = switch_io_sel_REG_0_0_1_0; // @[Router.scala 173:19]
  assign switch_io_sel_0_0_0_0 = switch_io_sel_REG_0_0_0_0; // @[Router.scala 173:19]
  assign switch_allocator_clock = clock;
  assign switch_allocator_reset = reset;
  assign switch_allocator_io_req_2_0_valid = ingress_unit_2_from_3_io_salloc_req_0_valid; // @[Router.scala 165:23]
  assign switch_allocator_io_req_2_0_bits_vc_sel_2_0 = ingress_unit_2_from_3_io_salloc_req_0_bits_vc_sel_2_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_2_0_bits_vc_sel_1_0 = ingress_unit_2_from_3_io_salloc_req_0_bits_vc_sel_1_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_2_0_bits_vc_sel_1_1 = ingress_unit_2_from_3_io_salloc_req_0_bits_vc_sel_1_1; // @[Router.scala 165:23]
  assign switch_allocator_io_req_2_0_bits_vc_sel_1_2 = ingress_unit_2_from_3_io_salloc_req_0_bits_vc_sel_1_2; // @[Router.scala 165:23]
  assign switch_allocator_io_req_2_0_bits_vc_sel_1_3 = ingress_unit_2_from_3_io_salloc_req_0_bits_vc_sel_1_3; // @[Router.scala 165:23]
  assign switch_allocator_io_req_2_0_bits_vc_sel_0_0 = ingress_unit_2_from_3_io_salloc_req_0_bits_vc_sel_0_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_2_0_bits_vc_sel_0_1 = ingress_unit_2_from_3_io_salloc_req_0_bits_vc_sel_0_1; // @[Router.scala 165:23]
  assign switch_allocator_io_req_2_0_bits_vc_sel_0_2 = ingress_unit_2_from_3_io_salloc_req_0_bits_vc_sel_0_2; // @[Router.scala 165:23]
  assign switch_allocator_io_req_2_0_bits_vc_sel_0_3 = ingress_unit_2_from_3_io_salloc_req_0_bits_vc_sel_0_3; // @[Router.scala 165:23]
  assign switch_allocator_io_req_2_0_bits_tail = ingress_unit_2_from_3_io_salloc_req_0_bits_tail; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_valid = input_unit_1_from_2_io_salloc_req_0_valid; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_vc_sel_2_0 = input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_2_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_vc_sel_1_0 = input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_1_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_vc_sel_1_1 = input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_1_1; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_vc_sel_1_2 = input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_1_2; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_vc_sel_1_3 = input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_1_3; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_vc_sel_0_0 = input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_0_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_vc_sel_0_1 = input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_0_1; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_vc_sel_0_2 = input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_0_2; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_vc_sel_0_3 = input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_0_3; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_tail = input_unit_1_from_2_io_salloc_req_0_bits_tail; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_valid = input_unit_0_from_0_io_salloc_req_0_valid; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_2_0 = input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_2_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_1_0 = input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_1_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_1_1 = input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_1_1; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_1_2 = input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_1_2; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_1_3 = input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_1_3; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_0_0 = input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_0_1 = input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_1; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_0_2 = input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_2; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_0_3 = input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_3; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_tail = input_unit_0_from_0_io_salloc_req_0_bits_tail; // @[Router.scala 165:23]
  assign vc_allocator_clock = clock;
  assign vc_allocator_reset = reset;
  assign vc_allocator_io_req_2_valid = ingress_unit_2_from_3_io_vcalloc_req_valid; // @[Router.scala 151:23]
  assign vc_allocator_io_req_2_bits_vc_sel_2_0 = ingress_unit_2_from_3_io_vcalloc_req_bits_vc_sel_2_0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_2_bits_vc_sel_1_0 = ingress_unit_2_from_3_io_vcalloc_req_bits_vc_sel_1_0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_2_bits_vc_sel_1_1 = ingress_unit_2_from_3_io_vcalloc_req_bits_vc_sel_1_1; // @[Router.scala 151:23]
  assign vc_allocator_io_req_2_bits_vc_sel_1_2 = ingress_unit_2_from_3_io_vcalloc_req_bits_vc_sel_1_2; // @[Router.scala 151:23]
  assign vc_allocator_io_req_2_bits_vc_sel_1_3 = ingress_unit_2_from_3_io_vcalloc_req_bits_vc_sel_1_3; // @[Router.scala 151:23]
  assign vc_allocator_io_req_2_bits_vc_sel_0_0 = ingress_unit_2_from_3_io_vcalloc_req_bits_vc_sel_0_0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_2_bits_vc_sel_0_1 = ingress_unit_2_from_3_io_vcalloc_req_bits_vc_sel_0_1; // @[Router.scala 151:23]
  assign vc_allocator_io_req_2_bits_vc_sel_0_2 = ingress_unit_2_from_3_io_vcalloc_req_bits_vc_sel_0_2; // @[Router.scala 151:23]
  assign vc_allocator_io_req_2_bits_vc_sel_0_3 = ingress_unit_2_from_3_io_vcalloc_req_bits_vc_sel_0_3; // @[Router.scala 151:23]
  assign vc_allocator_io_req_1_valid = input_unit_1_from_2_io_vcalloc_req_valid; // @[Router.scala 151:23]
  assign vc_allocator_io_req_1_bits_vc_sel_2_0 = input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_2_0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_1_bits_vc_sel_1_0 = input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_1_0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_1_bits_vc_sel_1_1 = input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_1_1; // @[Router.scala 151:23]
  assign vc_allocator_io_req_1_bits_vc_sel_1_2 = input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_1_2; // @[Router.scala 151:23]
  assign vc_allocator_io_req_1_bits_vc_sel_1_3 = input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_1_3; // @[Router.scala 151:23]
  assign vc_allocator_io_req_1_bits_vc_sel_0_0 = input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_0_0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_1_bits_vc_sel_0_1 = input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_0_1; // @[Router.scala 151:23]
  assign vc_allocator_io_req_1_bits_vc_sel_0_2 = input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_0_2; // @[Router.scala 151:23]
  assign vc_allocator_io_req_1_bits_vc_sel_0_3 = 1'h0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_valid = input_unit_0_from_0_io_vcalloc_req_valid; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_2_0 = input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_2_0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_1_0 = input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_1_0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_1_1 = input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_1_1; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_1_2 = input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_1_2; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_1_3 = input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_1_3; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_0_0 = input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_0_1 = input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_1; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_0_2 = input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_2; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_0_3 = 1'h0; // @[Router.scala 151:23]
  assign vc_allocator_io_channel_status_2_0_occupied = egress_unit_2_to_3_io_channel_status_0_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_1_0_occupied = output_unit_1_to_2_io_channel_status_0_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_1_1_occupied = output_unit_1_to_2_io_channel_status_1_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_1_2_occupied = output_unit_1_to_2_io_channel_status_2_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_1_3_occupied = output_unit_1_to_2_io_channel_status_3_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_0_0_occupied = output_unit_0_to_0_io_channel_status_0_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_0_1_occupied = output_unit_0_to_0_io_channel_status_1_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_0_2_occupied = output_unit_0_to_0_io_channel_status_2_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_0_3_occupied = output_unit_0_to_0_io_channel_status_3_occupied; // @[Router.scala 159:23]
  assign route_computer_io_req_2_bits_flow_ingress_node = ingress_unit_2_from_3_io_router_req_bits_flow_ingress_node; // @[Router.scala 146:23]
  assign route_computer_io_req_2_bits_flow_egress_node = ingress_unit_2_from_3_io_router_req_bits_flow_egress_node; // @[Router.scala 146:23]
  assign route_computer_io_req_1_bits_src_virt_id = input_unit_1_from_2_io_router_req_bits_src_virt_id; // @[Router.scala 146:23]
  assign route_computer_io_req_1_bits_flow_ingress_node = input_unit_1_from_2_io_router_req_bits_flow_ingress_node; // @[Router.scala 146:23]
  assign route_computer_io_req_1_bits_flow_egress_node = input_unit_1_from_2_io_router_req_bits_flow_egress_node; // @[Router.scala 146:23]
  assign route_computer_io_req_0_bits_src_virt_id = input_unit_0_from_0_io_router_req_bits_src_virt_id; // @[Router.scala 146:23]
  assign route_computer_io_req_0_bits_flow_ingress_node = input_unit_0_from_0_io_router_req_bits_flow_ingress_node; // @[Router.scala 146:23]
  assign route_computer_io_req_0_bits_flow_egress_node = input_unit_0_from_0_io_router_req_bits_flow_egress_node; // @[Router.scala 146:23]
  always @(posedge clock) begin
    switch_io_sel_REG_2_0_2_0 <= switch_allocator_io_switch_sel_2_0_2_0; // @[Router.scala 176:14]
    switch_io_sel_REG_2_0_1_0 <= switch_allocator_io_switch_sel_2_0_1_0; // @[Router.scala 176:14]
    switch_io_sel_REG_2_0_0_0 <= switch_allocator_io_switch_sel_2_0_0_0; // @[Router.scala 176:14]
    switch_io_sel_REG_1_0_2_0 <= switch_allocator_io_switch_sel_1_0_2_0; // @[Router.scala 176:14]
    switch_io_sel_REG_1_0_1_0 <= switch_allocator_io_switch_sel_1_0_1_0; // @[Router.scala 176:14]
    switch_io_sel_REG_1_0_0_0 <= switch_allocator_io_switch_sel_1_0_0_0; // @[Router.scala 176:14]
    switch_io_sel_REG_0_0_2_0 <= switch_allocator_io_switch_sel_0_0_2_0; // @[Router.scala 176:14]
    switch_io_sel_REG_0_0_1_0 <= switch_allocator_io_switch_sel_0_0_1_0; // @[Router.scala 176:14]
    switch_io_sel_REG_0_0_0_0 <= switch_allocator_io_switch_sel_0_0_0_0; // @[Router.scala 176:14]
    if (reset) begin // @[Router.scala 193:28]
      debug_tsc <= 64'h0; // @[Router.scala 193:28]
    end else begin
      debug_tsc <= _debug_tsc_T_1; // @[Router.scala 194:15]
    end
    if (reset) begin // @[Router.scala 195:31]
      debug_sample <= 64'h0; // @[Router.scala 195:31]
    end else if (debug_sample == _GEN_6) begin // @[Router.scala 198:47]
      debug_sample <= 64'h0; // @[Router.scala 198:62]
    end else begin
      debug_sample <= _debug_sample_T_1; // @[Router.scala 196:18]
    end
    if (reset) begin // @[Router.scala 201:29]
      util_ctr <= 64'h0; // @[Router.scala 201:29]
    end else begin
      util_ctr <= _util_ctr_T_1; // @[Router.scala 203:16]
    end
    if (reset) begin // @[Router.scala 202:26]
      fired <= 1'h0; // @[Router.scala 202:26]
    end else if (plusarg_reader_out != 20'h0 & _T_2 & fired) begin // @[Router.scala 205:81]
      fired <= auto_dest_nodes_in_0_flit_0_valid; // @[Router.scala 208:15]
    end else begin
      fired <= fired | auto_dest_nodes_in_0_flit_0_valid; // @[Router.scala 204:13]
    end
    if (reset) begin // @[Router.scala 201:29]
      util_ctr_1 <= 64'h0; // @[Router.scala 201:29]
    end else begin
      util_ctr_1 <= _util_ctr_T_3; // @[Router.scala 203:16]
    end
    if (reset) begin // @[Router.scala 202:26]
      fired_1 <= 1'h0; // @[Router.scala 202:26]
    end else if (plusarg_reader_out != 20'h0 & _T_2 & fired_1) begin // @[Router.scala 205:81]
      fired_1 <= auto_dest_nodes_in_1_flit_0_valid; // @[Router.scala 208:15]
    end else begin
      fired_1 <= fired_1 | auto_dest_nodes_in_1_flit_0_valid; // @[Router.scala 204:13]
    end
    if (reset) begin // @[Router.scala 201:29]
      util_ctr_2 <= 64'h0; // @[Router.scala 201:29]
    end else begin
      util_ctr_2 <= _util_ctr_T_5; // @[Router.scala 203:16]
    end
    if (reset) begin // @[Router.scala 202:26]
      fired_2 <= 1'h0; // @[Router.scala 202:26]
    end else if (plusarg_reader_out != 20'h0 & _T_2 & fired_2) begin // @[Router.scala 205:81]
      fired_2 <= _T_19; // @[Router.scala 208:15]
    end else begin
      fired_2 <= fired_2 | _T_19; // @[Router.scala 204:13]
    end
    if (reset) begin // @[Router.scala 201:29]
      util_ctr_3 <= 64'h0; // @[Router.scala 201:29]
    end else begin
      util_ctr_3 <= _util_ctr_T_7; // @[Router.scala 203:16]
    end
    if (reset) begin // @[Router.scala 202:26]
      fired_3 <= 1'h0; // @[Router.scala 202:26]
    end else if (plusarg_reader_out != 20'h0 & _T_2 & fired_3) begin // @[Router.scala 205:81]
      fired_3 <= x1_2_flit_valid; // @[Router.scala 208:15]
    end else begin
      fired_3 <= fired_3 | x1_2_flit_valid; // @[Router.scala 204:13]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8 & ~reset) begin
          $fwrite(32'h80000002,"nocsample %d 0 3 %d\n",debug_tsc,util_ctr); // @[Router.scala 207:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_16 & ~reset) begin
          $fwrite(32'h80000002,"nocsample %d 2 3 %d\n",debug_tsc,util_ctr_1); // @[Router.scala 207:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_25 & ~reset) begin
          $fwrite(32'h80000002,"nocsample %d i3 3 %d\n",debug_tsc,util_ctr_2); // @[Router.scala 207:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_34 & ~reset) begin
          $fwrite(32'h80000002,"nocsample %d 3 e3 %d\n",debug_tsc,util_ctr_3); // @[Router.scala 207:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  switch_io_sel_REG_2_0_2_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  switch_io_sel_REG_2_0_1_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  switch_io_sel_REG_2_0_0_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  switch_io_sel_REG_1_0_2_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  switch_io_sel_REG_1_0_1_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  switch_io_sel_REG_1_0_0_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  switch_io_sel_REG_0_0_2_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  switch_io_sel_REG_0_0_1_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  switch_io_sel_REG_0_0_0_0 = _RAND_8[0:0];
  _RAND_9 = {2{`RANDOM}};
  debug_tsc = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  debug_sample = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  util_ctr = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  fired = _RAND_12[0:0];
  _RAND_13 = {2{`RANDOM}};
  util_ctr_1 = _RAND_13[63:0];
  _RAND_14 = {1{`RANDOM}};
  fired_1 = _RAND_14[0:0];
  _RAND_15 = {2{`RANDOM}};
  util_ctr_2 = _RAND_15[63:0];
  _RAND_16 = {1{`RANDOM}};
  fired_2 = _RAND_16[0:0];
  _RAND_17 = {2{`RANDOM}};
  util_ctr_3 = _RAND_17[63:0];
  _RAND_18 = {1{`RANDOM}};
  fired_3 = _RAND_18[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ClockSinkDomain_3(
  output [1:0]  auto_routers_debug_out_va_stall_0,
  output [1:0]  auto_routers_debug_out_va_stall_1,
  output [1:0]  auto_routers_debug_out_sa_stall_0,
  output [1:0]  auto_routers_debug_out_sa_stall_1,
  output        auto_routers_egress_nodes_out_flit_valid,
  output        auto_routers_egress_nodes_out_flit_bits_head,
  output        auto_routers_egress_nodes_out_flit_bits_tail,
  output [63:0] auto_routers_egress_nodes_out_flit_bits_payload,
  output [1:0]  auto_routers_egress_nodes_out_flit_bits_ingress_id,
  output        auto_routers_ingress_nodes_in_flit_ready,
  input         auto_routers_ingress_nodes_in_flit_valid,
  input         auto_routers_ingress_nodes_in_flit_bits_head,
  input         auto_routers_ingress_nodes_in_flit_bits_tail,
  input  [63:0] auto_routers_ingress_nodes_in_flit_bits_payload,
  input  [1:0]  auto_routers_ingress_nodes_in_flit_bits_egress_id,
  output        auto_routers_source_nodes_out_1_flit_0_valid,
  output        auto_routers_source_nodes_out_1_flit_0_bits_head,
  output        auto_routers_source_nodes_out_1_flit_0_bits_tail,
  output [63:0] auto_routers_source_nodes_out_1_flit_0_bits_payload,
  output [1:0]  auto_routers_source_nodes_out_1_flit_0_bits_flow_ingress_node,
  output [1:0]  auto_routers_source_nodes_out_1_flit_0_bits_flow_egress_node,
  output [1:0]  auto_routers_source_nodes_out_1_flit_0_bits_virt_channel_id,
  input  [3:0]  auto_routers_source_nodes_out_1_credit_return,
  input  [3:0]  auto_routers_source_nodes_out_1_vc_free,
  output        auto_routers_source_nodes_out_0_flit_0_valid,
  output        auto_routers_source_nodes_out_0_flit_0_bits_head,
  output        auto_routers_source_nodes_out_0_flit_0_bits_tail,
  output [63:0] auto_routers_source_nodes_out_0_flit_0_bits_payload,
  output [1:0]  auto_routers_source_nodes_out_0_flit_0_bits_flow_ingress_node,
  output [1:0]  auto_routers_source_nodes_out_0_flit_0_bits_flow_egress_node,
  output [1:0]  auto_routers_source_nodes_out_0_flit_0_bits_virt_channel_id,
  input  [3:0]  auto_routers_source_nodes_out_0_credit_return,
  input  [3:0]  auto_routers_source_nodes_out_0_vc_free,
  input         auto_routers_dest_nodes_in_1_flit_0_valid,
  input         auto_routers_dest_nodes_in_1_flit_0_bits_head,
  input         auto_routers_dest_nodes_in_1_flit_0_bits_tail,
  input  [63:0] auto_routers_dest_nodes_in_1_flit_0_bits_payload,
  input  [1:0]  auto_routers_dest_nodes_in_1_flit_0_bits_flow_ingress_node,
  input  [1:0]  auto_routers_dest_nodes_in_1_flit_0_bits_flow_egress_node,
  input  [1:0]  auto_routers_dest_nodes_in_1_flit_0_bits_virt_channel_id,
  output [3:0]  auto_routers_dest_nodes_in_1_credit_return,
  output [3:0]  auto_routers_dest_nodes_in_1_vc_free,
  input         auto_routers_dest_nodes_in_0_flit_0_valid,
  input         auto_routers_dest_nodes_in_0_flit_0_bits_head,
  input         auto_routers_dest_nodes_in_0_flit_0_bits_tail,
  input  [63:0] auto_routers_dest_nodes_in_0_flit_0_bits_payload,
  input  [1:0]  auto_routers_dest_nodes_in_0_flit_0_bits_flow_ingress_node,
  input  [1:0]  auto_routers_dest_nodes_in_0_flit_0_bits_flow_egress_node,
  input  [1:0]  auto_routers_dest_nodes_in_0_flit_0_bits_virt_channel_id,
  output [3:0]  auto_routers_dest_nodes_in_0_credit_return,
  output [3:0]  auto_routers_dest_nodes_in_0_vc_free,
  input         auto_clock_in_clock,
  input         auto_clock_in_reset
);
  wire  routers_clock; // @[NoC.scala 64:22]
  wire  routers_reset; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_debug_out_va_stall_0; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_debug_out_va_stall_1; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_debug_out_sa_stall_0; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_debug_out_sa_stall_1; // @[NoC.scala 64:22]
  wire  routers_auto_egress_nodes_out_flit_valid; // @[NoC.scala 64:22]
  wire  routers_auto_egress_nodes_out_flit_bits_head; // @[NoC.scala 64:22]
  wire  routers_auto_egress_nodes_out_flit_bits_tail; // @[NoC.scala 64:22]
  wire [63:0] routers_auto_egress_nodes_out_flit_bits_payload; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_egress_nodes_out_flit_bits_ingress_id; // @[NoC.scala 64:22]
  wire  routers_auto_ingress_nodes_in_flit_ready; // @[NoC.scala 64:22]
  wire  routers_auto_ingress_nodes_in_flit_valid; // @[NoC.scala 64:22]
  wire  routers_auto_ingress_nodes_in_flit_bits_head; // @[NoC.scala 64:22]
  wire  routers_auto_ingress_nodes_in_flit_bits_tail; // @[NoC.scala 64:22]
  wire [63:0] routers_auto_ingress_nodes_in_flit_bits_payload; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_ingress_nodes_in_flit_bits_egress_id; // @[NoC.scala 64:22]
  wire  routers_auto_source_nodes_out_1_flit_0_valid; // @[NoC.scala 64:22]
  wire  routers_auto_source_nodes_out_1_flit_0_bits_head; // @[NoC.scala 64:22]
  wire  routers_auto_source_nodes_out_1_flit_0_bits_tail; // @[NoC.scala 64:22]
  wire [63:0] routers_auto_source_nodes_out_1_flit_0_bits_payload; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_source_nodes_out_1_flit_0_bits_flow_ingress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_source_nodes_out_1_flit_0_bits_flow_egress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_source_nodes_out_1_flit_0_bits_virt_channel_id; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_source_nodes_out_1_credit_return; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_source_nodes_out_1_vc_free; // @[NoC.scala 64:22]
  wire  routers_auto_source_nodes_out_0_flit_0_valid; // @[NoC.scala 64:22]
  wire  routers_auto_source_nodes_out_0_flit_0_bits_head; // @[NoC.scala 64:22]
  wire  routers_auto_source_nodes_out_0_flit_0_bits_tail; // @[NoC.scala 64:22]
  wire [63:0] routers_auto_source_nodes_out_0_flit_0_bits_payload; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_source_nodes_out_0_flit_0_bits_flow_ingress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_source_nodes_out_0_flit_0_bits_flow_egress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_source_nodes_out_0_flit_0_bits_virt_channel_id; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_source_nodes_out_0_credit_return; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_source_nodes_out_0_vc_free; // @[NoC.scala 64:22]
  wire  routers_auto_dest_nodes_in_1_flit_0_valid; // @[NoC.scala 64:22]
  wire  routers_auto_dest_nodes_in_1_flit_0_bits_head; // @[NoC.scala 64:22]
  wire  routers_auto_dest_nodes_in_1_flit_0_bits_tail; // @[NoC.scala 64:22]
  wire [63:0] routers_auto_dest_nodes_in_1_flit_0_bits_payload; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_dest_nodes_in_1_flit_0_bits_flow_ingress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_dest_nodes_in_1_flit_0_bits_flow_egress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_dest_nodes_in_1_flit_0_bits_virt_channel_id; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_dest_nodes_in_1_credit_return; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_dest_nodes_in_1_vc_free; // @[NoC.scala 64:22]
  wire  routers_auto_dest_nodes_in_0_flit_0_valid; // @[NoC.scala 64:22]
  wire  routers_auto_dest_nodes_in_0_flit_0_bits_head; // @[NoC.scala 64:22]
  wire  routers_auto_dest_nodes_in_0_flit_0_bits_tail; // @[NoC.scala 64:22]
  wire [63:0] routers_auto_dest_nodes_in_0_flit_0_bits_payload; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_dest_nodes_in_0_flit_0_bits_flow_ingress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_dest_nodes_in_0_flit_0_bits_flow_egress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_dest_nodes_in_0_flit_0_bits_virt_channel_id; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_dest_nodes_in_0_credit_return; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_dest_nodes_in_0_vc_free; // @[NoC.scala 64:22]
  Router_3 routers ( // @[NoC.scala 64:22]
    .clock(routers_clock),
    .reset(routers_reset),
    .auto_debug_out_va_stall_0(routers_auto_debug_out_va_stall_0),
    .auto_debug_out_va_stall_1(routers_auto_debug_out_va_stall_1),
    .auto_debug_out_sa_stall_0(routers_auto_debug_out_sa_stall_0),
    .auto_debug_out_sa_stall_1(routers_auto_debug_out_sa_stall_1),
    .auto_egress_nodes_out_flit_valid(routers_auto_egress_nodes_out_flit_valid),
    .auto_egress_nodes_out_flit_bits_head(routers_auto_egress_nodes_out_flit_bits_head),
    .auto_egress_nodes_out_flit_bits_tail(routers_auto_egress_nodes_out_flit_bits_tail),
    .auto_egress_nodes_out_flit_bits_payload(routers_auto_egress_nodes_out_flit_bits_payload),
    .auto_egress_nodes_out_flit_bits_ingress_id(routers_auto_egress_nodes_out_flit_bits_ingress_id),
    .auto_ingress_nodes_in_flit_ready(routers_auto_ingress_nodes_in_flit_ready),
    .auto_ingress_nodes_in_flit_valid(routers_auto_ingress_nodes_in_flit_valid),
    .auto_ingress_nodes_in_flit_bits_head(routers_auto_ingress_nodes_in_flit_bits_head),
    .auto_ingress_nodes_in_flit_bits_tail(routers_auto_ingress_nodes_in_flit_bits_tail),
    .auto_ingress_nodes_in_flit_bits_payload(routers_auto_ingress_nodes_in_flit_bits_payload),
    .auto_ingress_nodes_in_flit_bits_egress_id(routers_auto_ingress_nodes_in_flit_bits_egress_id),
    .auto_source_nodes_out_1_flit_0_valid(routers_auto_source_nodes_out_1_flit_0_valid),
    .auto_source_nodes_out_1_flit_0_bits_head(routers_auto_source_nodes_out_1_flit_0_bits_head),
    .auto_source_nodes_out_1_flit_0_bits_tail(routers_auto_source_nodes_out_1_flit_0_bits_tail),
    .auto_source_nodes_out_1_flit_0_bits_payload(routers_auto_source_nodes_out_1_flit_0_bits_payload),
    .auto_source_nodes_out_1_flit_0_bits_flow_ingress_node(routers_auto_source_nodes_out_1_flit_0_bits_flow_ingress_node
      ),
    .auto_source_nodes_out_1_flit_0_bits_flow_egress_node(routers_auto_source_nodes_out_1_flit_0_bits_flow_egress_node),
    .auto_source_nodes_out_1_flit_0_bits_virt_channel_id(routers_auto_source_nodes_out_1_flit_0_bits_virt_channel_id),
    .auto_source_nodes_out_1_credit_return(routers_auto_source_nodes_out_1_credit_return),
    .auto_source_nodes_out_1_vc_free(routers_auto_source_nodes_out_1_vc_free),
    .auto_source_nodes_out_0_flit_0_valid(routers_auto_source_nodes_out_0_flit_0_valid),
    .auto_source_nodes_out_0_flit_0_bits_head(routers_auto_source_nodes_out_0_flit_0_bits_head),
    .auto_source_nodes_out_0_flit_0_bits_tail(routers_auto_source_nodes_out_0_flit_0_bits_tail),
    .auto_source_nodes_out_0_flit_0_bits_payload(routers_auto_source_nodes_out_0_flit_0_bits_payload),
    .auto_source_nodes_out_0_flit_0_bits_flow_ingress_node(routers_auto_source_nodes_out_0_flit_0_bits_flow_ingress_node
      ),
    .auto_source_nodes_out_0_flit_0_bits_flow_egress_node(routers_auto_source_nodes_out_0_flit_0_bits_flow_egress_node),
    .auto_source_nodes_out_0_flit_0_bits_virt_channel_id(routers_auto_source_nodes_out_0_flit_0_bits_virt_channel_id),
    .auto_source_nodes_out_0_credit_return(routers_auto_source_nodes_out_0_credit_return),
    .auto_source_nodes_out_0_vc_free(routers_auto_source_nodes_out_0_vc_free),
    .auto_dest_nodes_in_1_flit_0_valid(routers_auto_dest_nodes_in_1_flit_0_valid),
    .auto_dest_nodes_in_1_flit_0_bits_head(routers_auto_dest_nodes_in_1_flit_0_bits_head),
    .auto_dest_nodes_in_1_flit_0_bits_tail(routers_auto_dest_nodes_in_1_flit_0_bits_tail),
    .auto_dest_nodes_in_1_flit_0_bits_payload(routers_auto_dest_nodes_in_1_flit_0_bits_payload),
    .auto_dest_nodes_in_1_flit_0_bits_flow_ingress_node(routers_auto_dest_nodes_in_1_flit_0_bits_flow_ingress_node),
    .auto_dest_nodes_in_1_flit_0_bits_flow_egress_node(routers_auto_dest_nodes_in_1_flit_0_bits_flow_egress_node),
    .auto_dest_nodes_in_1_flit_0_bits_virt_channel_id(routers_auto_dest_nodes_in_1_flit_0_bits_virt_channel_id),
    .auto_dest_nodes_in_1_credit_return(routers_auto_dest_nodes_in_1_credit_return),
    .auto_dest_nodes_in_1_vc_free(routers_auto_dest_nodes_in_1_vc_free),
    .auto_dest_nodes_in_0_flit_0_valid(routers_auto_dest_nodes_in_0_flit_0_valid),
    .auto_dest_nodes_in_0_flit_0_bits_head(routers_auto_dest_nodes_in_0_flit_0_bits_head),
    .auto_dest_nodes_in_0_flit_0_bits_tail(routers_auto_dest_nodes_in_0_flit_0_bits_tail),
    .auto_dest_nodes_in_0_flit_0_bits_payload(routers_auto_dest_nodes_in_0_flit_0_bits_payload),
    .auto_dest_nodes_in_0_flit_0_bits_flow_ingress_node(routers_auto_dest_nodes_in_0_flit_0_bits_flow_ingress_node),
    .auto_dest_nodes_in_0_flit_0_bits_flow_egress_node(routers_auto_dest_nodes_in_0_flit_0_bits_flow_egress_node),
    .auto_dest_nodes_in_0_flit_0_bits_virt_channel_id(routers_auto_dest_nodes_in_0_flit_0_bits_virt_channel_id),
    .auto_dest_nodes_in_0_credit_return(routers_auto_dest_nodes_in_0_credit_return),
    .auto_dest_nodes_in_0_vc_free(routers_auto_dest_nodes_in_0_vc_free)
  );
  assign auto_routers_debug_out_va_stall_0 = routers_auto_debug_out_va_stall_0; // @[LazyModule.scala 368:12]
  assign auto_routers_debug_out_va_stall_1 = routers_auto_debug_out_va_stall_1; // @[LazyModule.scala 368:12]
  assign auto_routers_debug_out_sa_stall_0 = routers_auto_debug_out_sa_stall_0; // @[LazyModule.scala 368:12]
  assign auto_routers_debug_out_sa_stall_1 = routers_auto_debug_out_sa_stall_1; // @[LazyModule.scala 368:12]
  assign auto_routers_egress_nodes_out_flit_valid = routers_auto_egress_nodes_out_flit_valid; // @[LazyModule.scala 368:12]
  assign auto_routers_egress_nodes_out_flit_bits_head = routers_auto_egress_nodes_out_flit_bits_head; // @[LazyModule.scala 368:12]
  assign auto_routers_egress_nodes_out_flit_bits_tail = routers_auto_egress_nodes_out_flit_bits_tail; // @[LazyModule.scala 368:12]
  assign auto_routers_egress_nodes_out_flit_bits_payload = routers_auto_egress_nodes_out_flit_bits_payload; // @[LazyModule.scala 368:12]
  assign auto_routers_egress_nodes_out_flit_bits_ingress_id = routers_auto_egress_nodes_out_flit_bits_ingress_id; // @[LazyModule.scala 368:12]
  assign auto_routers_ingress_nodes_in_flit_ready = routers_auto_ingress_nodes_in_flit_ready; // @[LazyModule.scala 366:16]
  assign auto_routers_source_nodes_out_1_flit_0_valid = routers_auto_source_nodes_out_1_flit_0_valid; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_1_flit_0_bits_head = routers_auto_source_nodes_out_1_flit_0_bits_head; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_1_flit_0_bits_tail = routers_auto_source_nodes_out_1_flit_0_bits_tail; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_1_flit_0_bits_payload = routers_auto_source_nodes_out_1_flit_0_bits_payload; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_1_flit_0_bits_flow_ingress_node =
    routers_auto_source_nodes_out_1_flit_0_bits_flow_ingress_node; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_1_flit_0_bits_flow_egress_node =
    routers_auto_source_nodes_out_1_flit_0_bits_flow_egress_node; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_1_flit_0_bits_virt_channel_id =
    routers_auto_source_nodes_out_1_flit_0_bits_virt_channel_id; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_0_flit_0_valid = routers_auto_source_nodes_out_0_flit_0_valid; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_0_flit_0_bits_head = routers_auto_source_nodes_out_0_flit_0_bits_head; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_0_flit_0_bits_tail = routers_auto_source_nodes_out_0_flit_0_bits_tail; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_0_flit_0_bits_payload = routers_auto_source_nodes_out_0_flit_0_bits_payload; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_0_flit_0_bits_flow_ingress_node =
    routers_auto_source_nodes_out_0_flit_0_bits_flow_ingress_node; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_0_flit_0_bits_flow_egress_node =
    routers_auto_source_nodes_out_0_flit_0_bits_flow_egress_node; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_0_flit_0_bits_virt_channel_id =
    routers_auto_source_nodes_out_0_flit_0_bits_virt_channel_id; // @[LazyModule.scala 368:12]
  assign auto_routers_dest_nodes_in_1_credit_return = routers_auto_dest_nodes_in_1_credit_return; // @[LazyModule.scala 366:16]
  assign auto_routers_dest_nodes_in_1_vc_free = routers_auto_dest_nodes_in_1_vc_free; // @[LazyModule.scala 366:16]
  assign auto_routers_dest_nodes_in_0_credit_return = routers_auto_dest_nodes_in_0_credit_return; // @[LazyModule.scala 366:16]
  assign auto_routers_dest_nodes_in_0_vc_free = routers_auto_dest_nodes_in_0_vc_free; // @[LazyModule.scala 366:16]
  assign routers_clock = auto_clock_in_clock; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign routers_reset = auto_clock_in_reset; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign routers_auto_ingress_nodes_in_flit_valid = auto_routers_ingress_nodes_in_flit_valid; // @[LazyModule.scala 366:16]
  assign routers_auto_ingress_nodes_in_flit_bits_head = auto_routers_ingress_nodes_in_flit_bits_head; // @[LazyModule.scala 366:16]
  assign routers_auto_ingress_nodes_in_flit_bits_tail = auto_routers_ingress_nodes_in_flit_bits_tail; // @[LazyModule.scala 366:16]
  assign routers_auto_ingress_nodes_in_flit_bits_payload = auto_routers_ingress_nodes_in_flit_bits_payload; // @[LazyModule.scala 366:16]
  assign routers_auto_ingress_nodes_in_flit_bits_egress_id = auto_routers_ingress_nodes_in_flit_bits_egress_id; // @[LazyModule.scala 366:16]
  assign routers_auto_source_nodes_out_1_credit_return = auto_routers_source_nodes_out_1_credit_return; // @[LazyModule.scala 368:12]
  assign routers_auto_source_nodes_out_1_vc_free = auto_routers_source_nodes_out_1_vc_free; // @[LazyModule.scala 368:12]
  assign routers_auto_source_nodes_out_0_credit_return = auto_routers_source_nodes_out_0_credit_return; // @[LazyModule.scala 368:12]
  assign routers_auto_source_nodes_out_0_vc_free = auto_routers_source_nodes_out_0_vc_free; // @[LazyModule.scala 368:12]
  assign routers_auto_dest_nodes_in_1_flit_0_valid = auto_routers_dest_nodes_in_1_flit_0_valid; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_1_flit_0_bits_head = auto_routers_dest_nodes_in_1_flit_0_bits_head; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_1_flit_0_bits_tail = auto_routers_dest_nodes_in_1_flit_0_bits_tail; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_1_flit_0_bits_payload = auto_routers_dest_nodes_in_1_flit_0_bits_payload; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_1_flit_0_bits_flow_ingress_node =
    auto_routers_dest_nodes_in_1_flit_0_bits_flow_ingress_node; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_1_flit_0_bits_flow_egress_node =
    auto_routers_dest_nodes_in_1_flit_0_bits_flow_egress_node; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_1_flit_0_bits_virt_channel_id =
    auto_routers_dest_nodes_in_1_flit_0_bits_virt_channel_id; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_0_flit_0_valid = auto_routers_dest_nodes_in_0_flit_0_valid; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_0_flit_0_bits_head = auto_routers_dest_nodes_in_0_flit_0_bits_head; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_0_flit_0_bits_tail = auto_routers_dest_nodes_in_0_flit_0_bits_tail; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_0_flit_0_bits_payload = auto_routers_dest_nodes_in_0_flit_0_bits_payload; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_0_flit_0_bits_flow_ingress_node =
    auto_routers_dest_nodes_in_0_flit_0_bits_flow_ingress_node; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_0_flit_0_bits_flow_egress_node =
    auto_routers_dest_nodes_in_0_flit_0_bits_flow_egress_node; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_0_flit_0_bits_virt_channel_id =
    auto_routers_dest_nodes_in_0_flit_0_bits_virt_channel_id; // @[LazyModule.scala 366:16]
endmodule
module NoC(
  input         clock,
  input         reset,
  output        io_ingress_3_flit_ready,
  input         io_ingress_3_flit_valid,
  input         io_ingress_3_flit_bits_head,
  input         io_ingress_3_flit_bits_tail,
  input  [63:0] io_ingress_3_flit_bits_payload,
  input  [1:0]  io_ingress_3_flit_bits_egress_id,
  output        io_ingress_2_flit_ready,
  input         io_ingress_2_flit_valid,
  input         io_ingress_2_flit_bits_head,
  input         io_ingress_2_flit_bits_tail,
  input  [63:0] io_ingress_2_flit_bits_payload,
  input  [1:0]  io_ingress_2_flit_bits_egress_id,
  output        io_ingress_1_flit_ready,
  input         io_ingress_1_flit_valid,
  input         io_ingress_1_flit_bits_head,
  input         io_ingress_1_flit_bits_tail,
  input  [63:0] io_ingress_1_flit_bits_payload,
  input  [1:0]  io_ingress_1_flit_bits_egress_id,
  output        io_ingress_0_flit_ready,
  input         io_ingress_0_flit_valid,
  input         io_ingress_0_flit_bits_head,
  input         io_ingress_0_flit_bits_tail,
  input  [63:0] io_ingress_0_flit_bits_payload,
  input  [1:0]  io_ingress_0_flit_bits_egress_id,
  output        io_egress_3_flit_valid,
  output        io_egress_3_flit_bits_head,
  output        io_egress_3_flit_bits_tail,
  output [63:0] io_egress_3_flit_bits_payload,
  output [1:0]  io_egress_3_flit_bits_ingress_id,
  output        io_egress_2_flit_valid,
  output        io_egress_2_flit_bits_head,
  output        io_egress_2_flit_bits_tail,
  output [63:0] io_egress_2_flit_bits_payload,
  output [1:0]  io_egress_2_flit_bits_ingress_id,
  output        io_egress_1_flit_valid,
  output        io_egress_1_flit_bits_head,
  output        io_egress_1_flit_bits_tail,
  output [63:0] io_egress_1_flit_bits_payload,
  output [1:0]  io_egress_1_flit_bits_ingress_id,
  output        io_egress_0_flit_valid,
  output        io_egress_0_flit_bits_head,
  output        io_egress_0_flit_bits_tail,
  output [63:0] io_egress_0_flit_bits_payload,
  output [1:0]  io_egress_0_flit_bits_ingress_id,
  input         io_router_clocks_0_clock,
  input         io_router_clocks_0_reset,
  input         io_router_clocks_1_clock,
  input         io_router_clocks_1_reset,
  input         io_router_clocks_2_clock,
  input         io_router_clocks_2_reset,
  input         io_router_clocks_3_clock,
  input         io_router_clocks_3_reset
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire [1:0] router_sink_domain_auto_routers_debug_out_va_stall_0; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_auto_routers_debug_out_va_stall_1; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_auto_routers_debug_out_sa_stall_0; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_auto_routers_debug_out_sa_stall_1; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_routers_egress_nodes_out_flit_valid; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_routers_egress_nodes_out_flit_bits_head; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_routers_egress_nodes_out_flit_bits_tail; // @[NoC.scala 38:40]
  wire [63:0] router_sink_domain_auto_routers_egress_nodes_out_flit_bits_payload; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_auto_routers_egress_nodes_out_flit_bits_ingress_id; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_routers_ingress_nodes_in_flit_ready; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_routers_ingress_nodes_in_flit_valid; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_routers_ingress_nodes_in_flit_bits_head; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_routers_ingress_nodes_in_flit_bits_tail; // @[NoC.scala 38:40]
  wire [63:0] router_sink_domain_auto_routers_ingress_nodes_in_flit_bits_payload; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_auto_routers_ingress_nodes_in_flit_bits_egress_id; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_routers_source_nodes_out_1_flit_0_valid; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_routers_source_nodes_out_1_flit_0_bits_head; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_routers_source_nodes_out_1_flit_0_bits_tail; // @[NoC.scala 38:40]
  wire [63:0] router_sink_domain_auto_routers_source_nodes_out_1_flit_0_bits_payload; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_auto_routers_source_nodes_out_1_flit_0_bits_flow_ingress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_auto_routers_source_nodes_out_1_flit_0_bits_flow_egress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_auto_routers_source_nodes_out_1_flit_0_bits_virt_channel_id; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_auto_routers_source_nodes_out_1_credit_return; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_auto_routers_source_nodes_out_1_vc_free; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_routers_source_nodes_out_0_flit_0_valid; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_routers_source_nodes_out_0_flit_0_bits_head; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_routers_source_nodes_out_0_flit_0_bits_tail; // @[NoC.scala 38:40]
  wire [63:0] router_sink_domain_auto_routers_source_nodes_out_0_flit_0_bits_payload; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_auto_routers_source_nodes_out_0_flit_0_bits_flow_ingress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_auto_routers_source_nodes_out_0_flit_0_bits_flow_egress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_auto_routers_source_nodes_out_0_flit_0_bits_virt_channel_id; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_auto_routers_source_nodes_out_0_credit_return; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_auto_routers_source_nodes_out_0_vc_free; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_routers_dest_nodes_in_1_flit_0_valid; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_routers_dest_nodes_in_1_flit_0_bits_head; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_routers_dest_nodes_in_1_flit_0_bits_tail; // @[NoC.scala 38:40]
  wire [63:0] router_sink_domain_auto_routers_dest_nodes_in_1_flit_0_bits_payload; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_auto_routers_dest_nodes_in_1_flit_0_bits_flow_ingress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_auto_routers_dest_nodes_in_1_flit_0_bits_flow_egress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_auto_routers_dest_nodes_in_1_flit_0_bits_virt_channel_id; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_auto_routers_dest_nodes_in_1_credit_return; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_auto_routers_dest_nodes_in_1_vc_free; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_routers_dest_nodes_in_0_flit_0_valid; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_routers_dest_nodes_in_0_flit_0_bits_head; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_routers_dest_nodes_in_0_flit_0_bits_tail; // @[NoC.scala 38:40]
  wire [63:0] router_sink_domain_auto_routers_dest_nodes_in_0_flit_0_bits_payload; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_auto_routers_dest_nodes_in_0_flit_0_bits_flow_ingress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_auto_routers_dest_nodes_in_0_flit_0_bits_flow_egress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_auto_routers_dest_nodes_in_0_flit_0_bits_virt_channel_id; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_auto_routers_dest_nodes_in_0_credit_return; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_auto_routers_dest_nodes_in_0_vc_free; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_clock_in_clock; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_clock_in_reset; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_1_auto_routers_debug_out_va_stall_0; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_1_auto_routers_debug_out_va_stall_1; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_1_auto_routers_debug_out_sa_stall_0; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_1_auto_routers_debug_out_sa_stall_1; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_routers_egress_nodes_out_flit_valid; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_routers_egress_nodes_out_flit_bits_head; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_routers_egress_nodes_out_flit_bits_tail; // @[NoC.scala 38:40]
  wire [63:0] router_sink_domain_1_auto_routers_egress_nodes_out_flit_bits_payload; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_1_auto_routers_egress_nodes_out_flit_bits_ingress_id; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_routers_ingress_nodes_in_flit_ready; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_routers_ingress_nodes_in_flit_valid; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_routers_ingress_nodes_in_flit_bits_head; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_routers_ingress_nodes_in_flit_bits_tail; // @[NoC.scala 38:40]
  wire [63:0] router_sink_domain_1_auto_routers_ingress_nodes_in_flit_bits_payload; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_1_auto_routers_ingress_nodes_in_flit_bits_egress_id; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_routers_source_nodes_out_1_flit_0_valid; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_routers_source_nodes_out_1_flit_0_bits_head; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_routers_source_nodes_out_1_flit_0_bits_tail; // @[NoC.scala 38:40]
  wire [63:0] router_sink_domain_1_auto_routers_source_nodes_out_1_flit_0_bits_payload; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_1_auto_routers_source_nodes_out_1_flit_0_bits_flow_ingress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_1_auto_routers_source_nodes_out_1_flit_0_bits_flow_egress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_1_auto_routers_source_nodes_out_1_flit_0_bits_virt_channel_id; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_1_auto_routers_source_nodes_out_1_credit_return; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_1_auto_routers_source_nodes_out_1_vc_free; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_routers_source_nodes_out_0_flit_0_valid; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_routers_source_nodes_out_0_flit_0_bits_head; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_routers_source_nodes_out_0_flit_0_bits_tail; // @[NoC.scala 38:40]
  wire [63:0] router_sink_domain_1_auto_routers_source_nodes_out_0_flit_0_bits_payload; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_1_auto_routers_source_nodes_out_0_flit_0_bits_flow_ingress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_1_auto_routers_source_nodes_out_0_flit_0_bits_flow_egress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_1_auto_routers_source_nodes_out_0_flit_0_bits_virt_channel_id; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_1_auto_routers_source_nodes_out_0_credit_return; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_1_auto_routers_source_nodes_out_0_vc_free; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_routers_dest_nodes_in_1_flit_0_valid; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_routers_dest_nodes_in_1_flit_0_bits_head; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_routers_dest_nodes_in_1_flit_0_bits_tail; // @[NoC.scala 38:40]
  wire [63:0] router_sink_domain_1_auto_routers_dest_nodes_in_1_flit_0_bits_payload; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_1_auto_routers_dest_nodes_in_1_flit_0_bits_flow_ingress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_1_auto_routers_dest_nodes_in_1_flit_0_bits_flow_egress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_1_auto_routers_dest_nodes_in_1_flit_0_bits_virt_channel_id; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_1_auto_routers_dest_nodes_in_1_credit_return; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_1_auto_routers_dest_nodes_in_1_vc_free; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_routers_dest_nodes_in_0_flit_0_valid; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_routers_dest_nodes_in_0_flit_0_bits_head; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_routers_dest_nodes_in_0_flit_0_bits_tail; // @[NoC.scala 38:40]
  wire [63:0] router_sink_domain_1_auto_routers_dest_nodes_in_0_flit_0_bits_payload; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_1_auto_routers_dest_nodes_in_0_flit_0_bits_flow_ingress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_1_auto_routers_dest_nodes_in_0_flit_0_bits_flow_egress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_1_auto_routers_dest_nodes_in_0_flit_0_bits_virt_channel_id; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_1_auto_routers_dest_nodes_in_0_credit_return; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_1_auto_routers_dest_nodes_in_0_vc_free; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_clock_in_clock; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_clock_in_reset; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_2_auto_routers_debug_out_va_stall_0; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_2_auto_routers_debug_out_va_stall_1; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_2_auto_routers_debug_out_sa_stall_0; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_2_auto_routers_debug_out_sa_stall_1; // @[NoC.scala 38:40]
  wire  router_sink_domain_2_auto_routers_egress_nodes_out_flit_valid; // @[NoC.scala 38:40]
  wire  router_sink_domain_2_auto_routers_egress_nodes_out_flit_bits_head; // @[NoC.scala 38:40]
  wire  router_sink_domain_2_auto_routers_egress_nodes_out_flit_bits_tail; // @[NoC.scala 38:40]
  wire [63:0] router_sink_domain_2_auto_routers_egress_nodes_out_flit_bits_payload; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_2_auto_routers_egress_nodes_out_flit_bits_ingress_id; // @[NoC.scala 38:40]
  wire  router_sink_domain_2_auto_routers_ingress_nodes_in_flit_ready; // @[NoC.scala 38:40]
  wire  router_sink_domain_2_auto_routers_ingress_nodes_in_flit_valid; // @[NoC.scala 38:40]
  wire  router_sink_domain_2_auto_routers_ingress_nodes_in_flit_bits_head; // @[NoC.scala 38:40]
  wire  router_sink_domain_2_auto_routers_ingress_nodes_in_flit_bits_tail; // @[NoC.scala 38:40]
  wire [63:0] router_sink_domain_2_auto_routers_ingress_nodes_in_flit_bits_payload; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_2_auto_routers_ingress_nodes_in_flit_bits_egress_id; // @[NoC.scala 38:40]
  wire  router_sink_domain_2_auto_routers_source_nodes_out_1_flit_0_valid; // @[NoC.scala 38:40]
  wire  router_sink_domain_2_auto_routers_source_nodes_out_1_flit_0_bits_head; // @[NoC.scala 38:40]
  wire  router_sink_domain_2_auto_routers_source_nodes_out_1_flit_0_bits_tail; // @[NoC.scala 38:40]
  wire [63:0] router_sink_domain_2_auto_routers_source_nodes_out_1_flit_0_bits_payload; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_2_auto_routers_source_nodes_out_1_flit_0_bits_flow_ingress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_2_auto_routers_source_nodes_out_1_flit_0_bits_flow_egress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_2_auto_routers_source_nodes_out_1_flit_0_bits_virt_channel_id; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_2_auto_routers_source_nodes_out_1_credit_return; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_2_auto_routers_source_nodes_out_1_vc_free; // @[NoC.scala 38:40]
  wire  router_sink_domain_2_auto_routers_source_nodes_out_0_flit_0_valid; // @[NoC.scala 38:40]
  wire  router_sink_domain_2_auto_routers_source_nodes_out_0_flit_0_bits_head; // @[NoC.scala 38:40]
  wire  router_sink_domain_2_auto_routers_source_nodes_out_0_flit_0_bits_tail; // @[NoC.scala 38:40]
  wire [63:0] router_sink_domain_2_auto_routers_source_nodes_out_0_flit_0_bits_payload; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_2_auto_routers_source_nodes_out_0_flit_0_bits_flow_ingress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_2_auto_routers_source_nodes_out_0_flit_0_bits_flow_egress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_2_auto_routers_source_nodes_out_0_flit_0_bits_virt_channel_id; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_2_auto_routers_source_nodes_out_0_credit_return; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_2_auto_routers_source_nodes_out_0_vc_free; // @[NoC.scala 38:40]
  wire  router_sink_domain_2_auto_routers_dest_nodes_in_1_flit_0_valid; // @[NoC.scala 38:40]
  wire  router_sink_domain_2_auto_routers_dest_nodes_in_1_flit_0_bits_head; // @[NoC.scala 38:40]
  wire  router_sink_domain_2_auto_routers_dest_nodes_in_1_flit_0_bits_tail; // @[NoC.scala 38:40]
  wire [63:0] router_sink_domain_2_auto_routers_dest_nodes_in_1_flit_0_bits_payload; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_2_auto_routers_dest_nodes_in_1_flit_0_bits_flow_ingress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_2_auto_routers_dest_nodes_in_1_flit_0_bits_flow_egress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_2_auto_routers_dest_nodes_in_1_flit_0_bits_virt_channel_id; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_2_auto_routers_dest_nodes_in_1_credit_return; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_2_auto_routers_dest_nodes_in_1_vc_free; // @[NoC.scala 38:40]
  wire  router_sink_domain_2_auto_routers_dest_nodes_in_0_flit_0_valid; // @[NoC.scala 38:40]
  wire  router_sink_domain_2_auto_routers_dest_nodes_in_0_flit_0_bits_head; // @[NoC.scala 38:40]
  wire  router_sink_domain_2_auto_routers_dest_nodes_in_0_flit_0_bits_tail; // @[NoC.scala 38:40]
  wire [63:0] router_sink_domain_2_auto_routers_dest_nodes_in_0_flit_0_bits_payload; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_2_auto_routers_dest_nodes_in_0_flit_0_bits_flow_ingress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_2_auto_routers_dest_nodes_in_0_flit_0_bits_flow_egress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_2_auto_routers_dest_nodes_in_0_flit_0_bits_virt_channel_id; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_2_auto_routers_dest_nodes_in_0_credit_return; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_2_auto_routers_dest_nodes_in_0_vc_free; // @[NoC.scala 38:40]
  wire  router_sink_domain_2_auto_clock_in_clock; // @[NoC.scala 38:40]
  wire  router_sink_domain_2_auto_clock_in_reset; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_3_auto_routers_debug_out_va_stall_0; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_3_auto_routers_debug_out_va_stall_1; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_3_auto_routers_debug_out_sa_stall_0; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_3_auto_routers_debug_out_sa_stall_1; // @[NoC.scala 38:40]
  wire  router_sink_domain_3_auto_routers_egress_nodes_out_flit_valid; // @[NoC.scala 38:40]
  wire  router_sink_domain_3_auto_routers_egress_nodes_out_flit_bits_head; // @[NoC.scala 38:40]
  wire  router_sink_domain_3_auto_routers_egress_nodes_out_flit_bits_tail; // @[NoC.scala 38:40]
  wire [63:0] router_sink_domain_3_auto_routers_egress_nodes_out_flit_bits_payload; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_3_auto_routers_egress_nodes_out_flit_bits_ingress_id; // @[NoC.scala 38:40]
  wire  router_sink_domain_3_auto_routers_ingress_nodes_in_flit_ready; // @[NoC.scala 38:40]
  wire  router_sink_domain_3_auto_routers_ingress_nodes_in_flit_valid; // @[NoC.scala 38:40]
  wire  router_sink_domain_3_auto_routers_ingress_nodes_in_flit_bits_head; // @[NoC.scala 38:40]
  wire  router_sink_domain_3_auto_routers_ingress_nodes_in_flit_bits_tail; // @[NoC.scala 38:40]
  wire [63:0] router_sink_domain_3_auto_routers_ingress_nodes_in_flit_bits_payload; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_3_auto_routers_ingress_nodes_in_flit_bits_egress_id; // @[NoC.scala 38:40]
  wire  router_sink_domain_3_auto_routers_source_nodes_out_1_flit_0_valid; // @[NoC.scala 38:40]
  wire  router_sink_domain_3_auto_routers_source_nodes_out_1_flit_0_bits_head; // @[NoC.scala 38:40]
  wire  router_sink_domain_3_auto_routers_source_nodes_out_1_flit_0_bits_tail; // @[NoC.scala 38:40]
  wire [63:0] router_sink_domain_3_auto_routers_source_nodes_out_1_flit_0_bits_payload; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_3_auto_routers_source_nodes_out_1_flit_0_bits_flow_ingress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_3_auto_routers_source_nodes_out_1_flit_0_bits_flow_egress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_3_auto_routers_source_nodes_out_1_flit_0_bits_virt_channel_id; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_3_auto_routers_source_nodes_out_1_credit_return; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_3_auto_routers_source_nodes_out_1_vc_free; // @[NoC.scala 38:40]
  wire  router_sink_domain_3_auto_routers_source_nodes_out_0_flit_0_valid; // @[NoC.scala 38:40]
  wire  router_sink_domain_3_auto_routers_source_nodes_out_0_flit_0_bits_head; // @[NoC.scala 38:40]
  wire  router_sink_domain_3_auto_routers_source_nodes_out_0_flit_0_bits_tail; // @[NoC.scala 38:40]
  wire [63:0] router_sink_domain_3_auto_routers_source_nodes_out_0_flit_0_bits_payload; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_3_auto_routers_source_nodes_out_0_flit_0_bits_flow_ingress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_3_auto_routers_source_nodes_out_0_flit_0_bits_flow_egress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_3_auto_routers_source_nodes_out_0_flit_0_bits_virt_channel_id; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_3_auto_routers_source_nodes_out_0_credit_return; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_3_auto_routers_source_nodes_out_0_vc_free; // @[NoC.scala 38:40]
  wire  router_sink_domain_3_auto_routers_dest_nodes_in_1_flit_0_valid; // @[NoC.scala 38:40]
  wire  router_sink_domain_3_auto_routers_dest_nodes_in_1_flit_0_bits_head; // @[NoC.scala 38:40]
  wire  router_sink_domain_3_auto_routers_dest_nodes_in_1_flit_0_bits_tail; // @[NoC.scala 38:40]
  wire [63:0] router_sink_domain_3_auto_routers_dest_nodes_in_1_flit_0_bits_payload; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_3_auto_routers_dest_nodes_in_1_flit_0_bits_flow_ingress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_3_auto_routers_dest_nodes_in_1_flit_0_bits_flow_egress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_3_auto_routers_dest_nodes_in_1_flit_0_bits_virt_channel_id; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_3_auto_routers_dest_nodes_in_1_credit_return; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_3_auto_routers_dest_nodes_in_1_vc_free; // @[NoC.scala 38:40]
  wire  router_sink_domain_3_auto_routers_dest_nodes_in_0_flit_0_valid; // @[NoC.scala 38:40]
  wire  router_sink_domain_3_auto_routers_dest_nodes_in_0_flit_0_bits_head; // @[NoC.scala 38:40]
  wire  router_sink_domain_3_auto_routers_dest_nodes_in_0_flit_0_bits_tail; // @[NoC.scala 38:40]
  wire [63:0] router_sink_domain_3_auto_routers_dest_nodes_in_0_flit_0_bits_payload; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_3_auto_routers_dest_nodes_in_0_flit_0_bits_flow_ingress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_3_auto_routers_dest_nodes_in_0_flit_0_bits_flow_egress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_3_auto_routers_dest_nodes_in_0_flit_0_bits_virt_channel_id; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_3_auto_routers_dest_nodes_in_0_credit_return; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_3_auto_routers_dest_nodes_in_0_vc_free; // @[NoC.scala 38:40]
  wire  router_sink_domain_3_auto_clock_in_clock; // @[NoC.scala 38:40]
  wire  router_sink_domain_3_auto_clock_in_reset; // @[NoC.scala 38:40]
  reg [63:0] debug_va_stall_ctr; // @[NoC.scala 160:37]
  reg [63:0] debug_sa_stall_ctr; // @[NoC.scala 161:37]
  wire [63:0] debug_any_stall_ctr = debug_va_stall_ctr + debug_sa_stall_ctr; // @[NoC.scala 162:50]
  wire [1:0] bundleIn_0_4_va_stall_0 = router_sink_domain_auto_routers_debug_out_va_stall_0; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  wire [1:0] bundleIn_0_4_va_stall_1 = router_sink_domain_auto_routers_debug_out_va_stall_1; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  wire [1:0] _debug_va_stall_ctr_T_1 = bundleIn_0_4_va_stall_0 + bundleIn_0_4_va_stall_1; // @[NoC.scala 163:91]
  wire [2:0] _debug_va_stall_ctr_T_2 = {{1'd0}, _debug_va_stall_ctr_T_1}; // @[NoC.scala 163:91]
  wire [1:0] bundleIn_0_5_va_stall_0 = router_sink_domain_1_auto_routers_debug_out_va_stall_0; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  wire [1:0] bundleIn_0_5_va_stall_1 = router_sink_domain_1_auto_routers_debug_out_va_stall_1; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  wire [1:0] _debug_va_stall_ctr_T_5 = bundleIn_0_5_va_stall_0 + bundleIn_0_5_va_stall_1; // @[NoC.scala 163:91]
  wire [2:0] _debug_va_stall_ctr_T_6 = {{1'd0}, _debug_va_stall_ctr_T_5}; // @[NoC.scala 163:91]
  wire [1:0] bundleIn_0_6_va_stall_0 = router_sink_domain_2_auto_routers_debug_out_va_stall_0; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  wire [1:0] bundleIn_0_6_va_stall_1 = router_sink_domain_2_auto_routers_debug_out_va_stall_1; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  wire [1:0] _debug_va_stall_ctr_T_9 = bundleIn_0_6_va_stall_0 + bundleIn_0_6_va_stall_1; // @[NoC.scala 163:91]
  wire [2:0] _debug_va_stall_ctr_T_10 = {{1'd0}, _debug_va_stall_ctr_T_9}; // @[NoC.scala 163:91]
  wire [1:0] bundleIn_0_7_va_stall_0 = router_sink_domain_3_auto_routers_debug_out_va_stall_0; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  wire [1:0] bundleIn_0_7_va_stall_1 = router_sink_domain_3_auto_routers_debug_out_va_stall_1; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  wire [1:0] _debug_va_stall_ctr_T_13 = bundleIn_0_7_va_stall_0 + bundleIn_0_7_va_stall_1; // @[NoC.scala 163:91]
  wire [2:0] _debug_va_stall_ctr_T_14 = {{1'd0}, _debug_va_stall_ctr_T_13}; // @[NoC.scala 163:91]
  wire [1:0] _debug_va_stall_ctr_T_17 = _debug_va_stall_ctr_T_2[1:0] + _debug_va_stall_ctr_T_6[1:0]; // @[NoC.scala 163:104]
  wire [1:0] _debug_va_stall_ctr_T_19 = _debug_va_stall_ctr_T_17 + _debug_va_stall_ctr_T_10[1:0]; // @[NoC.scala 163:104]
  wire [1:0] _debug_va_stall_ctr_T_21 = _debug_va_stall_ctr_T_19 + _debug_va_stall_ctr_T_14[1:0]; // @[NoC.scala 163:104]
  wire [63:0] _GEN_0 = {{62'd0}, _debug_va_stall_ctr_T_21}; // @[NoC.scala 163:46]
  wire [63:0] _debug_va_stall_ctr_T_23 = debug_va_stall_ctr + _GEN_0; // @[NoC.scala 163:46]
  wire [1:0] bundleIn_0_4_sa_stall_0 = router_sink_domain_auto_routers_debug_out_sa_stall_0; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  wire [1:0] bundleIn_0_4_sa_stall_1 = router_sink_domain_auto_routers_debug_out_sa_stall_1; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  wire [1:0] _debug_sa_stall_ctr_T_1 = bundleIn_0_4_sa_stall_0 + bundleIn_0_4_sa_stall_1; // @[NoC.scala 164:91]
  wire [2:0] _debug_sa_stall_ctr_T_2 = {{1'd0}, _debug_sa_stall_ctr_T_1}; // @[NoC.scala 164:91]
  wire [1:0] bundleIn_0_5_sa_stall_0 = router_sink_domain_1_auto_routers_debug_out_sa_stall_0; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  wire [1:0] bundleIn_0_5_sa_stall_1 = router_sink_domain_1_auto_routers_debug_out_sa_stall_1; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  wire [1:0] _debug_sa_stall_ctr_T_5 = bundleIn_0_5_sa_stall_0 + bundleIn_0_5_sa_stall_1; // @[NoC.scala 164:91]
  wire [2:0] _debug_sa_stall_ctr_T_6 = {{1'd0}, _debug_sa_stall_ctr_T_5}; // @[NoC.scala 164:91]
  wire [1:0] bundleIn_0_6_sa_stall_0 = router_sink_domain_2_auto_routers_debug_out_sa_stall_0; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  wire [1:0] bundleIn_0_6_sa_stall_1 = router_sink_domain_2_auto_routers_debug_out_sa_stall_1; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  wire [1:0] _debug_sa_stall_ctr_T_9 = bundleIn_0_6_sa_stall_0 + bundleIn_0_6_sa_stall_1; // @[NoC.scala 164:91]
  wire [2:0] _debug_sa_stall_ctr_T_10 = {{1'd0}, _debug_sa_stall_ctr_T_9}; // @[NoC.scala 164:91]
  wire [1:0] bundleIn_0_7_sa_stall_0 = router_sink_domain_3_auto_routers_debug_out_sa_stall_0; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  wire [1:0] bundleIn_0_7_sa_stall_1 = router_sink_domain_3_auto_routers_debug_out_sa_stall_1; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  wire [1:0] _debug_sa_stall_ctr_T_13 = bundleIn_0_7_sa_stall_0 + bundleIn_0_7_sa_stall_1; // @[NoC.scala 164:91]
  wire [2:0] _debug_sa_stall_ctr_T_14 = {{1'd0}, _debug_sa_stall_ctr_T_13}; // @[NoC.scala 164:91]
  wire [1:0] _debug_sa_stall_ctr_T_17 = _debug_sa_stall_ctr_T_2[1:0] + _debug_sa_stall_ctr_T_6[1:0]; // @[NoC.scala 164:104]
  wire [1:0] _debug_sa_stall_ctr_T_19 = _debug_sa_stall_ctr_T_17 + _debug_sa_stall_ctr_T_10[1:0]; // @[NoC.scala 164:104]
  wire [1:0] _debug_sa_stall_ctr_T_21 = _debug_sa_stall_ctr_T_19 + _debug_sa_stall_ctr_T_14[1:0]; // @[NoC.scala 164:104]
  wire [63:0] _GEN_1 = {{62'd0}, _debug_sa_stall_ctr_T_21}; // @[NoC.scala 164:46]
  wire [63:0] _debug_sa_stall_ctr_T_23 = debug_sa_stall_ctr + _GEN_1; // @[NoC.scala 164:46]
  ClockSinkDomain router_sink_domain ( // @[NoC.scala 38:40]
    .auto_routers_debug_out_va_stall_0(router_sink_domain_auto_routers_debug_out_va_stall_0),
    .auto_routers_debug_out_va_stall_1(router_sink_domain_auto_routers_debug_out_va_stall_1),
    .auto_routers_debug_out_sa_stall_0(router_sink_domain_auto_routers_debug_out_sa_stall_0),
    .auto_routers_debug_out_sa_stall_1(router_sink_domain_auto_routers_debug_out_sa_stall_1),
    .auto_routers_egress_nodes_out_flit_valid(router_sink_domain_auto_routers_egress_nodes_out_flit_valid),
    .auto_routers_egress_nodes_out_flit_bits_head(router_sink_domain_auto_routers_egress_nodes_out_flit_bits_head),
    .auto_routers_egress_nodes_out_flit_bits_tail(router_sink_domain_auto_routers_egress_nodes_out_flit_bits_tail),
    .auto_routers_egress_nodes_out_flit_bits_payload(router_sink_domain_auto_routers_egress_nodes_out_flit_bits_payload)
      ,
    .auto_routers_egress_nodes_out_flit_bits_ingress_id(
      router_sink_domain_auto_routers_egress_nodes_out_flit_bits_ingress_id),
    .auto_routers_ingress_nodes_in_flit_ready(router_sink_domain_auto_routers_ingress_nodes_in_flit_ready),
    .auto_routers_ingress_nodes_in_flit_valid(router_sink_domain_auto_routers_ingress_nodes_in_flit_valid),
    .auto_routers_ingress_nodes_in_flit_bits_head(router_sink_domain_auto_routers_ingress_nodes_in_flit_bits_head),
    .auto_routers_ingress_nodes_in_flit_bits_tail(router_sink_domain_auto_routers_ingress_nodes_in_flit_bits_tail),
    .auto_routers_ingress_nodes_in_flit_bits_payload(router_sink_domain_auto_routers_ingress_nodes_in_flit_bits_payload)
      ,
    .auto_routers_ingress_nodes_in_flit_bits_egress_id(
      router_sink_domain_auto_routers_ingress_nodes_in_flit_bits_egress_id),
    .auto_routers_source_nodes_out_1_flit_0_valid(router_sink_domain_auto_routers_source_nodes_out_1_flit_0_valid),
    .auto_routers_source_nodes_out_1_flit_0_bits_head(
      router_sink_domain_auto_routers_source_nodes_out_1_flit_0_bits_head),
    .auto_routers_source_nodes_out_1_flit_0_bits_tail(
      router_sink_domain_auto_routers_source_nodes_out_1_flit_0_bits_tail),
    .auto_routers_source_nodes_out_1_flit_0_bits_payload(
      router_sink_domain_auto_routers_source_nodes_out_1_flit_0_bits_payload),
    .auto_routers_source_nodes_out_1_flit_0_bits_flow_ingress_node(
      router_sink_domain_auto_routers_source_nodes_out_1_flit_0_bits_flow_ingress_node),
    .auto_routers_source_nodes_out_1_flit_0_bits_flow_egress_node(
      router_sink_domain_auto_routers_source_nodes_out_1_flit_0_bits_flow_egress_node),
    .auto_routers_source_nodes_out_1_flit_0_bits_virt_channel_id(
      router_sink_domain_auto_routers_source_nodes_out_1_flit_0_bits_virt_channel_id),
    .auto_routers_source_nodes_out_1_credit_return(router_sink_domain_auto_routers_source_nodes_out_1_credit_return),
    .auto_routers_source_nodes_out_1_vc_free(router_sink_domain_auto_routers_source_nodes_out_1_vc_free),
    .auto_routers_source_nodes_out_0_flit_0_valid(router_sink_domain_auto_routers_source_nodes_out_0_flit_0_valid),
    .auto_routers_source_nodes_out_0_flit_0_bits_head(
      router_sink_domain_auto_routers_source_nodes_out_0_flit_0_bits_head),
    .auto_routers_source_nodes_out_0_flit_0_bits_tail(
      router_sink_domain_auto_routers_source_nodes_out_0_flit_0_bits_tail),
    .auto_routers_source_nodes_out_0_flit_0_bits_payload(
      router_sink_domain_auto_routers_source_nodes_out_0_flit_0_bits_payload),
    .auto_routers_source_nodes_out_0_flit_0_bits_flow_ingress_node(
      router_sink_domain_auto_routers_source_nodes_out_0_flit_0_bits_flow_ingress_node),
    .auto_routers_source_nodes_out_0_flit_0_bits_flow_egress_node(
      router_sink_domain_auto_routers_source_nodes_out_0_flit_0_bits_flow_egress_node),
    .auto_routers_source_nodes_out_0_flit_0_bits_virt_channel_id(
      router_sink_domain_auto_routers_source_nodes_out_0_flit_0_bits_virt_channel_id),
    .auto_routers_source_nodes_out_0_credit_return(router_sink_domain_auto_routers_source_nodes_out_0_credit_return),
    .auto_routers_source_nodes_out_0_vc_free(router_sink_domain_auto_routers_source_nodes_out_0_vc_free),
    .auto_routers_dest_nodes_in_1_flit_0_valid(router_sink_domain_auto_routers_dest_nodes_in_1_flit_0_valid),
    .auto_routers_dest_nodes_in_1_flit_0_bits_head(router_sink_domain_auto_routers_dest_nodes_in_1_flit_0_bits_head),
    .auto_routers_dest_nodes_in_1_flit_0_bits_tail(router_sink_domain_auto_routers_dest_nodes_in_1_flit_0_bits_tail),
    .auto_routers_dest_nodes_in_1_flit_0_bits_payload(
      router_sink_domain_auto_routers_dest_nodes_in_1_flit_0_bits_payload),
    .auto_routers_dest_nodes_in_1_flit_0_bits_flow_ingress_node(
      router_sink_domain_auto_routers_dest_nodes_in_1_flit_0_bits_flow_ingress_node),
    .auto_routers_dest_nodes_in_1_flit_0_bits_flow_egress_node(
      router_sink_domain_auto_routers_dest_nodes_in_1_flit_0_bits_flow_egress_node),
    .auto_routers_dest_nodes_in_1_flit_0_bits_virt_channel_id(
      router_sink_domain_auto_routers_dest_nodes_in_1_flit_0_bits_virt_channel_id),
    .auto_routers_dest_nodes_in_1_credit_return(router_sink_domain_auto_routers_dest_nodes_in_1_credit_return),
    .auto_routers_dest_nodes_in_1_vc_free(router_sink_domain_auto_routers_dest_nodes_in_1_vc_free),
    .auto_routers_dest_nodes_in_0_flit_0_valid(router_sink_domain_auto_routers_dest_nodes_in_0_flit_0_valid),
    .auto_routers_dest_nodes_in_0_flit_0_bits_head(router_sink_domain_auto_routers_dest_nodes_in_0_flit_0_bits_head),
    .auto_routers_dest_nodes_in_0_flit_0_bits_tail(router_sink_domain_auto_routers_dest_nodes_in_0_flit_0_bits_tail),
    .auto_routers_dest_nodes_in_0_flit_0_bits_payload(
      router_sink_domain_auto_routers_dest_nodes_in_0_flit_0_bits_payload),
    .auto_routers_dest_nodes_in_0_flit_0_bits_flow_ingress_node(
      router_sink_domain_auto_routers_dest_nodes_in_0_flit_0_bits_flow_ingress_node),
    .auto_routers_dest_nodes_in_0_flit_0_bits_flow_egress_node(
      router_sink_domain_auto_routers_dest_nodes_in_0_flit_0_bits_flow_egress_node),
    .auto_routers_dest_nodes_in_0_flit_0_bits_virt_channel_id(
      router_sink_domain_auto_routers_dest_nodes_in_0_flit_0_bits_virt_channel_id),
    .auto_routers_dest_nodes_in_0_credit_return(router_sink_domain_auto_routers_dest_nodes_in_0_credit_return),
    .auto_routers_dest_nodes_in_0_vc_free(router_sink_domain_auto_routers_dest_nodes_in_0_vc_free),
    .auto_clock_in_clock(router_sink_domain_auto_clock_in_clock),
    .auto_clock_in_reset(router_sink_domain_auto_clock_in_reset)
  );
  ClockSinkDomain_1 router_sink_domain_1 ( // @[NoC.scala 38:40]
    .auto_routers_debug_out_va_stall_0(router_sink_domain_1_auto_routers_debug_out_va_stall_0),
    .auto_routers_debug_out_va_stall_1(router_sink_domain_1_auto_routers_debug_out_va_stall_1),
    .auto_routers_debug_out_sa_stall_0(router_sink_domain_1_auto_routers_debug_out_sa_stall_0),
    .auto_routers_debug_out_sa_stall_1(router_sink_domain_1_auto_routers_debug_out_sa_stall_1),
    .auto_routers_egress_nodes_out_flit_valid(router_sink_domain_1_auto_routers_egress_nodes_out_flit_valid),
    .auto_routers_egress_nodes_out_flit_bits_head(router_sink_domain_1_auto_routers_egress_nodes_out_flit_bits_head),
    .auto_routers_egress_nodes_out_flit_bits_tail(router_sink_domain_1_auto_routers_egress_nodes_out_flit_bits_tail),
    .auto_routers_egress_nodes_out_flit_bits_payload(
      router_sink_domain_1_auto_routers_egress_nodes_out_flit_bits_payload),
    .auto_routers_egress_nodes_out_flit_bits_ingress_id(
      router_sink_domain_1_auto_routers_egress_nodes_out_flit_bits_ingress_id),
    .auto_routers_ingress_nodes_in_flit_ready(router_sink_domain_1_auto_routers_ingress_nodes_in_flit_ready),
    .auto_routers_ingress_nodes_in_flit_valid(router_sink_domain_1_auto_routers_ingress_nodes_in_flit_valid),
    .auto_routers_ingress_nodes_in_flit_bits_head(router_sink_domain_1_auto_routers_ingress_nodes_in_flit_bits_head),
    .auto_routers_ingress_nodes_in_flit_bits_tail(router_sink_domain_1_auto_routers_ingress_nodes_in_flit_bits_tail),
    .auto_routers_ingress_nodes_in_flit_bits_payload(
      router_sink_domain_1_auto_routers_ingress_nodes_in_flit_bits_payload),
    .auto_routers_ingress_nodes_in_flit_bits_egress_id(
      router_sink_domain_1_auto_routers_ingress_nodes_in_flit_bits_egress_id),
    .auto_routers_source_nodes_out_1_flit_0_valid(router_sink_domain_1_auto_routers_source_nodes_out_1_flit_0_valid),
    .auto_routers_source_nodes_out_1_flit_0_bits_head(
      router_sink_domain_1_auto_routers_source_nodes_out_1_flit_0_bits_head),
    .auto_routers_source_nodes_out_1_flit_0_bits_tail(
      router_sink_domain_1_auto_routers_source_nodes_out_1_flit_0_bits_tail),
    .auto_routers_source_nodes_out_1_flit_0_bits_payload(
      router_sink_domain_1_auto_routers_source_nodes_out_1_flit_0_bits_payload),
    .auto_routers_source_nodes_out_1_flit_0_bits_flow_ingress_node(
      router_sink_domain_1_auto_routers_source_nodes_out_1_flit_0_bits_flow_ingress_node),
    .auto_routers_source_nodes_out_1_flit_0_bits_flow_egress_node(
      router_sink_domain_1_auto_routers_source_nodes_out_1_flit_0_bits_flow_egress_node),
    .auto_routers_source_nodes_out_1_flit_0_bits_virt_channel_id(
      router_sink_domain_1_auto_routers_source_nodes_out_1_flit_0_bits_virt_channel_id),
    .auto_routers_source_nodes_out_1_credit_return(router_sink_domain_1_auto_routers_source_nodes_out_1_credit_return),
    .auto_routers_source_nodes_out_1_vc_free(router_sink_domain_1_auto_routers_source_nodes_out_1_vc_free),
    .auto_routers_source_nodes_out_0_flit_0_valid(router_sink_domain_1_auto_routers_source_nodes_out_0_flit_0_valid),
    .auto_routers_source_nodes_out_0_flit_0_bits_head(
      router_sink_domain_1_auto_routers_source_nodes_out_0_flit_0_bits_head),
    .auto_routers_source_nodes_out_0_flit_0_bits_tail(
      router_sink_domain_1_auto_routers_source_nodes_out_0_flit_0_bits_tail),
    .auto_routers_source_nodes_out_0_flit_0_bits_payload(
      router_sink_domain_1_auto_routers_source_nodes_out_0_flit_0_bits_payload),
    .auto_routers_source_nodes_out_0_flit_0_bits_flow_ingress_node(
      router_sink_domain_1_auto_routers_source_nodes_out_0_flit_0_bits_flow_ingress_node),
    .auto_routers_source_nodes_out_0_flit_0_bits_flow_egress_node(
      router_sink_domain_1_auto_routers_source_nodes_out_0_flit_0_bits_flow_egress_node),
    .auto_routers_source_nodes_out_0_flit_0_bits_virt_channel_id(
      router_sink_domain_1_auto_routers_source_nodes_out_0_flit_0_bits_virt_channel_id),
    .auto_routers_source_nodes_out_0_credit_return(router_sink_domain_1_auto_routers_source_nodes_out_0_credit_return),
    .auto_routers_source_nodes_out_0_vc_free(router_sink_domain_1_auto_routers_source_nodes_out_0_vc_free),
    .auto_routers_dest_nodes_in_1_flit_0_valid(router_sink_domain_1_auto_routers_dest_nodes_in_1_flit_0_valid),
    .auto_routers_dest_nodes_in_1_flit_0_bits_head(router_sink_domain_1_auto_routers_dest_nodes_in_1_flit_0_bits_head),
    .auto_routers_dest_nodes_in_1_flit_0_bits_tail(router_sink_domain_1_auto_routers_dest_nodes_in_1_flit_0_bits_tail),
    .auto_routers_dest_nodes_in_1_flit_0_bits_payload(
      router_sink_domain_1_auto_routers_dest_nodes_in_1_flit_0_bits_payload),
    .auto_routers_dest_nodes_in_1_flit_0_bits_flow_ingress_node(
      router_sink_domain_1_auto_routers_dest_nodes_in_1_flit_0_bits_flow_ingress_node),
    .auto_routers_dest_nodes_in_1_flit_0_bits_flow_egress_node(
      router_sink_domain_1_auto_routers_dest_nodes_in_1_flit_0_bits_flow_egress_node),
    .auto_routers_dest_nodes_in_1_flit_0_bits_virt_channel_id(
      router_sink_domain_1_auto_routers_dest_nodes_in_1_flit_0_bits_virt_channel_id),
    .auto_routers_dest_nodes_in_1_credit_return(router_sink_domain_1_auto_routers_dest_nodes_in_1_credit_return),
    .auto_routers_dest_nodes_in_1_vc_free(router_sink_domain_1_auto_routers_dest_nodes_in_1_vc_free),
    .auto_routers_dest_nodes_in_0_flit_0_valid(router_sink_domain_1_auto_routers_dest_nodes_in_0_flit_0_valid),
    .auto_routers_dest_nodes_in_0_flit_0_bits_head(router_sink_domain_1_auto_routers_dest_nodes_in_0_flit_0_bits_head),
    .auto_routers_dest_nodes_in_0_flit_0_bits_tail(router_sink_domain_1_auto_routers_dest_nodes_in_0_flit_0_bits_tail),
    .auto_routers_dest_nodes_in_0_flit_0_bits_payload(
      router_sink_domain_1_auto_routers_dest_nodes_in_0_flit_0_bits_payload),
    .auto_routers_dest_nodes_in_0_flit_0_bits_flow_ingress_node(
      router_sink_domain_1_auto_routers_dest_nodes_in_0_flit_0_bits_flow_ingress_node),
    .auto_routers_dest_nodes_in_0_flit_0_bits_flow_egress_node(
      router_sink_domain_1_auto_routers_dest_nodes_in_0_flit_0_bits_flow_egress_node),
    .auto_routers_dest_nodes_in_0_flit_0_bits_virt_channel_id(
      router_sink_domain_1_auto_routers_dest_nodes_in_0_flit_0_bits_virt_channel_id),
    .auto_routers_dest_nodes_in_0_credit_return(router_sink_domain_1_auto_routers_dest_nodes_in_0_credit_return),
    .auto_routers_dest_nodes_in_0_vc_free(router_sink_domain_1_auto_routers_dest_nodes_in_0_vc_free),
    .auto_clock_in_clock(router_sink_domain_1_auto_clock_in_clock),
    .auto_clock_in_reset(router_sink_domain_1_auto_clock_in_reset)
  );
  ClockSinkDomain_2 router_sink_domain_2 ( // @[NoC.scala 38:40]
    .auto_routers_debug_out_va_stall_0(router_sink_domain_2_auto_routers_debug_out_va_stall_0),
    .auto_routers_debug_out_va_stall_1(router_sink_domain_2_auto_routers_debug_out_va_stall_1),
    .auto_routers_debug_out_sa_stall_0(router_sink_domain_2_auto_routers_debug_out_sa_stall_0),
    .auto_routers_debug_out_sa_stall_1(router_sink_domain_2_auto_routers_debug_out_sa_stall_1),
    .auto_routers_egress_nodes_out_flit_valid(router_sink_domain_2_auto_routers_egress_nodes_out_flit_valid),
    .auto_routers_egress_nodes_out_flit_bits_head(router_sink_domain_2_auto_routers_egress_nodes_out_flit_bits_head),
    .auto_routers_egress_nodes_out_flit_bits_tail(router_sink_domain_2_auto_routers_egress_nodes_out_flit_bits_tail),
    .auto_routers_egress_nodes_out_flit_bits_payload(
      router_sink_domain_2_auto_routers_egress_nodes_out_flit_bits_payload),
    .auto_routers_egress_nodes_out_flit_bits_ingress_id(
      router_sink_domain_2_auto_routers_egress_nodes_out_flit_bits_ingress_id),
    .auto_routers_ingress_nodes_in_flit_ready(router_sink_domain_2_auto_routers_ingress_nodes_in_flit_ready),
    .auto_routers_ingress_nodes_in_flit_valid(router_sink_domain_2_auto_routers_ingress_nodes_in_flit_valid),
    .auto_routers_ingress_nodes_in_flit_bits_head(router_sink_domain_2_auto_routers_ingress_nodes_in_flit_bits_head),
    .auto_routers_ingress_nodes_in_flit_bits_tail(router_sink_domain_2_auto_routers_ingress_nodes_in_flit_bits_tail),
    .auto_routers_ingress_nodes_in_flit_bits_payload(
      router_sink_domain_2_auto_routers_ingress_nodes_in_flit_bits_payload),
    .auto_routers_ingress_nodes_in_flit_bits_egress_id(
      router_sink_domain_2_auto_routers_ingress_nodes_in_flit_bits_egress_id),
    .auto_routers_source_nodes_out_1_flit_0_valid(router_sink_domain_2_auto_routers_source_nodes_out_1_flit_0_valid),
    .auto_routers_source_nodes_out_1_flit_0_bits_head(
      router_sink_domain_2_auto_routers_source_nodes_out_1_flit_0_bits_head),
    .auto_routers_source_nodes_out_1_flit_0_bits_tail(
      router_sink_domain_2_auto_routers_source_nodes_out_1_flit_0_bits_tail),
    .auto_routers_source_nodes_out_1_flit_0_bits_payload(
      router_sink_domain_2_auto_routers_source_nodes_out_1_flit_0_bits_payload),
    .auto_routers_source_nodes_out_1_flit_0_bits_flow_ingress_node(
      router_sink_domain_2_auto_routers_source_nodes_out_1_flit_0_bits_flow_ingress_node),
    .auto_routers_source_nodes_out_1_flit_0_bits_flow_egress_node(
      router_sink_domain_2_auto_routers_source_nodes_out_1_flit_0_bits_flow_egress_node),
    .auto_routers_source_nodes_out_1_flit_0_bits_virt_channel_id(
      router_sink_domain_2_auto_routers_source_nodes_out_1_flit_0_bits_virt_channel_id),
    .auto_routers_source_nodes_out_1_credit_return(router_sink_domain_2_auto_routers_source_nodes_out_1_credit_return),
    .auto_routers_source_nodes_out_1_vc_free(router_sink_domain_2_auto_routers_source_nodes_out_1_vc_free),
    .auto_routers_source_nodes_out_0_flit_0_valid(router_sink_domain_2_auto_routers_source_nodes_out_0_flit_0_valid),
    .auto_routers_source_nodes_out_0_flit_0_bits_head(
      router_sink_domain_2_auto_routers_source_nodes_out_0_flit_0_bits_head),
    .auto_routers_source_nodes_out_0_flit_0_bits_tail(
      router_sink_domain_2_auto_routers_source_nodes_out_0_flit_0_bits_tail),
    .auto_routers_source_nodes_out_0_flit_0_bits_payload(
      router_sink_domain_2_auto_routers_source_nodes_out_0_flit_0_bits_payload),
    .auto_routers_source_nodes_out_0_flit_0_bits_flow_ingress_node(
      router_sink_domain_2_auto_routers_source_nodes_out_0_flit_0_bits_flow_ingress_node),
    .auto_routers_source_nodes_out_0_flit_0_bits_flow_egress_node(
      router_sink_domain_2_auto_routers_source_nodes_out_0_flit_0_bits_flow_egress_node),
    .auto_routers_source_nodes_out_0_flit_0_bits_virt_channel_id(
      router_sink_domain_2_auto_routers_source_nodes_out_0_flit_0_bits_virt_channel_id),
    .auto_routers_source_nodes_out_0_credit_return(router_sink_domain_2_auto_routers_source_nodes_out_0_credit_return),
    .auto_routers_source_nodes_out_0_vc_free(router_sink_domain_2_auto_routers_source_nodes_out_0_vc_free),
    .auto_routers_dest_nodes_in_1_flit_0_valid(router_sink_domain_2_auto_routers_dest_nodes_in_1_flit_0_valid),
    .auto_routers_dest_nodes_in_1_flit_0_bits_head(router_sink_domain_2_auto_routers_dest_nodes_in_1_flit_0_bits_head),
    .auto_routers_dest_nodes_in_1_flit_0_bits_tail(router_sink_domain_2_auto_routers_dest_nodes_in_1_flit_0_bits_tail),
    .auto_routers_dest_nodes_in_1_flit_0_bits_payload(
      router_sink_domain_2_auto_routers_dest_nodes_in_1_flit_0_bits_payload),
    .auto_routers_dest_nodes_in_1_flit_0_bits_flow_ingress_node(
      router_sink_domain_2_auto_routers_dest_nodes_in_1_flit_0_bits_flow_ingress_node),
    .auto_routers_dest_nodes_in_1_flit_0_bits_flow_egress_node(
      router_sink_domain_2_auto_routers_dest_nodes_in_1_flit_0_bits_flow_egress_node),
    .auto_routers_dest_nodes_in_1_flit_0_bits_virt_channel_id(
      router_sink_domain_2_auto_routers_dest_nodes_in_1_flit_0_bits_virt_channel_id),
    .auto_routers_dest_nodes_in_1_credit_return(router_sink_domain_2_auto_routers_dest_nodes_in_1_credit_return),
    .auto_routers_dest_nodes_in_1_vc_free(router_sink_domain_2_auto_routers_dest_nodes_in_1_vc_free),
    .auto_routers_dest_nodes_in_0_flit_0_valid(router_sink_domain_2_auto_routers_dest_nodes_in_0_flit_0_valid),
    .auto_routers_dest_nodes_in_0_flit_0_bits_head(router_sink_domain_2_auto_routers_dest_nodes_in_0_flit_0_bits_head),
    .auto_routers_dest_nodes_in_0_flit_0_bits_tail(router_sink_domain_2_auto_routers_dest_nodes_in_0_flit_0_bits_tail),
    .auto_routers_dest_nodes_in_0_flit_0_bits_payload(
      router_sink_domain_2_auto_routers_dest_nodes_in_0_flit_0_bits_payload),
    .auto_routers_dest_nodes_in_0_flit_0_bits_flow_ingress_node(
      router_sink_domain_2_auto_routers_dest_nodes_in_0_flit_0_bits_flow_ingress_node),
    .auto_routers_dest_nodes_in_0_flit_0_bits_flow_egress_node(
      router_sink_domain_2_auto_routers_dest_nodes_in_0_flit_0_bits_flow_egress_node),
    .auto_routers_dest_nodes_in_0_flit_0_bits_virt_channel_id(
      router_sink_domain_2_auto_routers_dest_nodes_in_0_flit_0_bits_virt_channel_id),
    .auto_routers_dest_nodes_in_0_credit_return(router_sink_domain_2_auto_routers_dest_nodes_in_0_credit_return),
    .auto_routers_dest_nodes_in_0_vc_free(router_sink_domain_2_auto_routers_dest_nodes_in_0_vc_free),
    .auto_clock_in_clock(router_sink_domain_2_auto_clock_in_clock),
    .auto_clock_in_reset(router_sink_domain_2_auto_clock_in_reset)
  );
  ClockSinkDomain_3 router_sink_domain_3 ( // @[NoC.scala 38:40]
    .auto_routers_debug_out_va_stall_0(router_sink_domain_3_auto_routers_debug_out_va_stall_0),
    .auto_routers_debug_out_va_stall_1(router_sink_domain_3_auto_routers_debug_out_va_stall_1),
    .auto_routers_debug_out_sa_stall_0(router_sink_domain_3_auto_routers_debug_out_sa_stall_0),
    .auto_routers_debug_out_sa_stall_1(router_sink_domain_3_auto_routers_debug_out_sa_stall_1),
    .auto_routers_egress_nodes_out_flit_valid(router_sink_domain_3_auto_routers_egress_nodes_out_flit_valid),
    .auto_routers_egress_nodes_out_flit_bits_head(router_sink_domain_3_auto_routers_egress_nodes_out_flit_bits_head),
    .auto_routers_egress_nodes_out_flit_bits_tail(router_sink_domain_3_auto_routers_egress_nodes_out_flit_bits_tail),
    .auto_routers_egress_nodes_out_flit_bits_payload(
      router_sink_domain_3_auto_routers_egress_nodes_out_flit_bits_payload),
    .auto_routers_egress_nodes_out_flit_bits_ingress_id(
      router_sink_domain_3_auto_routers_egress_nodes_out_flit_bits_ingress_id),
    .auto_routers_ingress_nodes_in_flit_ready(router_sink_domain_3_auto_routers_ingress_nodes_in_flit_ready),
    .auto_routers_ingress_nodes_in_flit_valid(router_sink_domain_3_auto_routers_ingress_nodes_in_flit_valid),
    .auto_routers_ingress_nodes_in_flit_bits_head(router_sink_domain_3_auto_routers_ingress_nodes_in_flit_bits_head),
    .auto_routers_ingress_nodes_in_flit_bits_tail(router_sink_domain_3_auto_routers_ingress_nodes_in_flit_bits_tail),
    .auto_routers_ingress_nodes_in_flit_bits_payload(
      router_sink_domain_3_auto_routers_ingress_nodes_in_flit_bits_payload),
    .auto_routers_ingress_nodes_in_flit_bits_egress_id(
      router_sink_domain_3_auto_routers_ingress_nodes_in_flit_bits_egress_id),
    .auto_routers_source_nodes_out_1_flit_0_valid(router_sink_domain_3_auto_routers_source_nodes_out_1_flit_0_valid),
    .auto_routers_source_nodes_out_1_flit_0_bits_head(
      router_sink_domain_3_auto_routers_source_nodes_out_1_flit_0_bits_head),
    .auto_routers_source_nodes_out_1_flit_0_bits_tail(
      router_sink_domain_3_auto_routers_source_nodes_out_1_flit_0_bits_tail),
    .auto_routers_source_nodes_out_1_flit_0_bits_payload(
      router_sink_domain_3_auto_routers_source_nodes_out_1_flit_0_bits_payload),
    .auto_routers_source_nodes_out_1_flit_0_bits_flow_ingress_node(
      router_sink_domain_3_auto_routers_source_nodes_out_1_flit_0_bits_flow_ingress_node),
    .auto_routers_source_nodes_out_1_flit_0_bits_flow_egress_node(
      router_sink_domain_3_auto_routers_source_nodes_out_1_flit_0_bits_flow_egress_node),
    .auto_routers_source_nodes_out_1_flit_0_bits_virt_channel_id(
      router_sink_domain_3_auto_routers_source_nodes_out_1_flit_0_bits_virt_channel_id),
    .auto_routers_source_nodes_out_1_credit_return(router_sink_domain_3_auto_routers_source_nodes_out_1_credit_return),
    .auto_routers_source_nodes_out_1_vc_free(router_sink_domain_3_auto_routers_source_nodes_out_1_vc_free),
    .auto_routers_source_nodes_out_0_flit_0_valid(router_sink_domain_3_auto_routers_source_nodes_out_0_flit_0_valid),
    .auto_routers_source_nodes_out_0_flit_0_bits_head(
      router_sink_domain_3_auto_routers_source_nodes_out_0_flit_0_bits_head),
    .auto_routers_source_nodes_out_0_flit_0_bits_tail(
      router_sink_domain_3_auto_routers_source_nodes_out_0_flit_0_bits_tail),
    .auto_routers_source_nodes_out_0_flit_0_bits_payload(
      router_sink_domain_3_auto_routers_source_nodes_out_0_flit_0_bits_payload),
    .auto_routers_source_nodes_out_0_flit_0_bits_flow_ingress_node(
      router_sink_domain_3_auto_routers_source_nodes_out_0_flit_0_bits_flow_ingress_node),
    .auto_routers_source_nodes_out_0_flit_0_bits_flow_egress_node(
      router_sink_domain_3_auto_routers_source_nodes_out_0_flit_0_bits_flow_egress_node),
    .auto_routers_source_nodes_out_0_flit_0_bits_virt_channel_id(
      router_sink_domain_3_auto_routers_source_nodes_out_0_flit_0_bits_virt_channel_id),
    .auto_routers_source_nodes_out_0_credit_return(router_sink_domain_3_auto_routers_source_nodes_out_0_credit_return),
    .auto_routers_source_nodes_out_0_vc_free(router_sink_domain_3_auto_routers_source_nodes_out_0_vc_free),
    .auto_routers_dest_nodes_in_1_flit_0_valid(router_sink_domain_3_auto_routers_dest_nodes_in_1_flit_0_valid),
    .auto_routers_dest_nodes_in_1_flit_0_bits_head(router_sink_domain_3_auto_routers_dest_nodes_in_1_flit_0_bits_head),
    .auto_routers_dest_nodes_in_1_flit_0_bits_tail(router_sink_domain_3_auto_routers_dest_nodes_in_1_flit_0_bits_tail),
    .auto_routers_dest_nodes_in_1_flit_0_bits_payload(
      router_sink_domain_3_auto_routers_dest_nodes_in_1_flit_0_bits_payload),
    .auto_routers_dest_nodes_in_1_flit_0_bits_flow_ingress_node(
      router_sink_domain_3_auto_routers_dest_nodes_in_1_flit_0_bits_flow_ingress_node),
    .auto_routers_dest_nodes_in_1_flit_0_bits_flow_egress_node(
      router_sink_domain_3_auto_routers_dest_nodes_in_1_flit_0_bits_flow_egress_node),
    .auto_routers_dest_nodes_in_1_flit_0_bits_virt_channel_id(
      router_sink_domain_3_auto_routers_dest_nodes_in_1_flit_0_bits_virt_channel_id),
    .auto_routers_dest_nodes_in_1_credit_return(router_sink_domain_3_auto_routers_dest_nodes_in_1_credit_return),
    .auto_routers_dest_nodes_in_1_vc_free(router_sink_domain_3_auto_routers_dest_nodes_in_1_vc_free),
    .auto_routers_dest_nodes_in_0_flit_0_valid(router_sink_domain_3_auto_routers_dest_nodes_in_0_flit_0_valid),
    .auto_routers_dest_nodes_in_0_flit_0_bits_head(router_sink_domain_3_auto_routers_dest_nodes_in_0_flit_0_bits_head),
    .auto_routers_dest_nodes_in_0_flit_0_bits_tail(router_sink_domain_3_auto_routers_dest_nodes_in_0_flit_0_bits_tail),
    .auto_routers_dest_nodes_in_0_flit_0_bits_payload(
      router_sink_domain_3_auto_routers_dest_nodes_in_0_flit_0_bits_payload),
    .auto_routers_dest_nodes_in_0_flit_0_bits_flow_ingress_node(
      router_sink_domain_3_auto_routers_dest_nodes_in_0_flit_0_bits_flow_ingress_node),
    .auto_routers_dest_nodes_in_0_flit_0_bits_flow_egress_node(
      router_sink_domain_3_auto_routers_dest_nodes_in_0_flit_0_bits_flow_egress_node),
    .auto_routers_dest_nodes_in_0_flit_0_bits_virt_channel_id(
      router_sink_domain_3_auto_routers_dest_nodes_in_0_flit_0_bits_virt_channel_id),
    .auto_routers_dest_nodes_in_0_credit_return(router_sink_domain_3_auto_routers_dest_nodes_in_0_credit_return),
    .auto_routers_dest_nodes_in_0_vc_free(router_sink_domain_3_auto_routers_dest_nodes_in_0_vc_free),
    .auto_clock_in_clock(router_sink_domain_3_auto_clock_in_clock),
    .auto_clock_in_reset(router_sink_domain_3_auto_clock_in_reset)
  );
  assign io_ingress_3_flit_ready = router_sink_domain_3_auto_routers_ingress_nodes_in_flit_ready; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign io_ingress_2_flit_ready = router_sink_domain_2_auto_routers_ingress_nodes_in_flit_ready; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign io_ingress_1_flit_ready = router_sink_domain_1_auto_routers_ingress_nodes_in_flit_ready; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign io_ingress_0_flit_ready = router_sink_domain_auto_routers_ingress_nodes_in_flit_ready; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign io_egress_3_flit_valid = router_sink_domain_3_auto_routers_egress_nodes_out_flit_valid; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign io_egress_3_flit_bits_head = router_sink_domain_3_auto_routers_egress_nodes_out_flit_bits_head; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign io_egress_3_flit_bits_tail = router_sink_domain_3_auto_routers_egress_nodes_out_flit_bits_tail; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign io_egress_3_flit_bits_payload = router_sink_domain_3_auto_routers_egress_nodes_out_flit_bits_payload; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign io_egress_3_flit_bits_ingress_id = router_sink_domain_3_auto_routers_egress_nodes_out_flit_bits_ingress_id; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign io_egress_2_flit_valid = router_sink_domain_2_auto_routers_egress_nodes_out_flit_valid; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign io_egress_2_flit_bits_head = router_sink_domain_2_auto_routers_egress_nodes_out_flit_bits_head; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign io_egress_2_flit_bits_tail = router_sink_domain_2_auto_routers_egress_nodes_out_flit_bits_tail; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign io_egress_2_flit_bits_payload = router_sink_domain_2_auto_routers_egress_nodes_out_flit_bits_payload; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign io_egress_2_flit_bits_ingress_id = router_sink_domain_2_auto_routers_egress_nodes_out_flit_bits_ingress_id; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign io_egress_1_flit_valid = router_sink_domain_1_auto_routers_egress_nodes_out_flit_valid; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign io_egress_1_flit_bits_head = router_sink_domain_1_auto_routers_egress_nodes_out_flit_bits_head; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign io_egress_1_flit_bits_tail = router_sink_domain_1_auto_routers_egress_nodes_out_flit_bits_tail; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign io_egress_1_flit_bits_payload = router_sink_domain_1_auto_routers_egress_nodes_out_flit_bits_payload; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign io_egress_1_flit_bits_ingress_id = router_sink_domain_1_auto_routers_egress_nodes_out_flit_bits_ingress_id; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign io_egress_0_flit_valid = router_sink_domain_auto_routers_egress_nodes_out_flit_valid; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign io_egress_0_flit_bits_head = router_sink_domain_auto_routers_egress_nodes_out_flit_bits_head; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign io_egress_0_flit_bits_tail = router_sink_domain_auto_routers_egress_nodes_out_flit_bits_tail; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign io_egress_0_flit_bits_payload = router_sink_domain_auto_routers_egress_nodes_out_flit_bits_payload; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign io_egress_0_flit_bits_ingress_id = router_sink_domain_auto_routers_egress_nodes_out_flit_bits_ingress_id; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign router_sink_domain_auto_routers_ingress_nodes_in_flit_valid = io_ingress_0_flit_valid; // @[Nodes.scala 1212:84 NoC.scala 145:78]
  assign router_sink_domain_auto_routers_ingress_nodes_in_flit_bits_head = io_ingress_0_flit_bits_head; // @[Nodes.scala 1212:84 NoC.scala 145:78]
  assign router_sink_domain_auto_routers_ingress_nodes_in_flit_bits_tail = io_ingress_0_flit_bits_tail; // @[Nodes.scala 1212:84 NoC.scala 145:78]
  assign router_sink_domain_auto_routers_ingress_nodes_in_flit_bits_payload = io_ingress_0_flit_bits_payload; // @[Nodes.scala 1212:84 NoC.scala 145:78]
  assign router_sink_domain_auto_routers_ingress_nodes_in_flit_bits_egress_id = io_ingress_0_flit_bits_egress_id; // @[Nodes.scala 1212:84 NoC.scala 145:78]
  assign router_sink_domain_auto_routers_source_nodes_out_1_credit_return =
    router_sink_domain_3_auto_routers_dest_nodes_in_0_credit_return; // @[LazyModule.scala 355:16]
  assign router_sink_domain_auto_routers_source_nodes_out_1_vc_free =
    router_sink_domain_3_auto_routers_dest_nodes_in_0_vc_free; // @[LazyModule.scala 355:16]
  assign router_sink_domain_auto_routers_source_nodes_out_0_credit_return =
    router_sink_domain_1_auto_routers_dest_nodes_in_0_credit_return; // @[LazyModule.scala 355:16]
  assign router_sink_domain_auto_routers_source_nodes_out_0_vc_free =
    router_sink_domain_1_auto_routers_dest_nodes_in_0_vc_free; // @[LazyModule.scala 355:16]
  assign router_sink_domain_auto_routers_dest_nodes_in_1_flit_0_valid =
    router_sink_domain_3_auto_routers_source_nodes_out_0_flit_0_valid; // @[LazyModule.scala 353:16]
  assign router_sink_domain_auto_routers_dest_nodes_in_1_flit_0_bits_head =
    router_sink_domain_3_auto_routers_source_nodes_out_0_flit_0_bits_head; // @[LazyModule.scala 353:16]
  assign router_sink_domain_auto_routers_dest_nodes_in_1_flit_0_bits_tail =
    router_sink_domain_3_auto_routers_source_nodes_out_0_flit_0_bits_tail; // @[LazyModule.scala 353:16]
  assign router_sink_domain_auto_routers_dest_nodes_in_1_flit_0_bits_payload =
    router_sink_domain_3_auto_routers_source_nodes_out_0_flit_0_bits_payload; // @[LazyModule.scala 353:16]
  assign router_sink_domain_auto_routers_dest_nodes_in_1_flit_0_bits_flow_ingress_node =
    router_sink_domain_3_auto_routers_source_nodes_out_0_flit_0_bits_flow_ingress_node; // @[LazyModule.scala 353:16]
  assign router_sink_domain_auto_routers_dest_nodes_in_1_flit_0_bits_flow_egress_node =
    router_sink_domain_3_auto_routers_source_nodes_out_0_flit_0_bits_flow_egress_node; // @[LazyModule.scala 353:16]
  assign router_sink_domain_auto_routers_dest_nodes_in_1_flit_0_bits_virt_channel_id =
    router_sink_domain_3_auto_routers_source_nodes_out_0_flit_0_bits_virt_channel_id; // @[LazyModule.scala 353:16]
  assign router_sink_domain_auto_routers_dest_nodes_in_0_flit_0_valid =
    router_sink_domain_1_auto_routers_source_nodes_out_0_flit_0_valid; // @[LazyModule.scala 353:16]
  assign router_sink_domain_auto_routers_dest_nodes_in_0_flit_0_bits_head =
    router_sink_domain_1_auto_routers_source_nodes_out_0_flit_0_bits_head; // @[LazyModule.scala 353:16]
  assign router_sink_domain_auto_routers_dest_nodes_in_0_flit_0_bits_tail =
    router_sink_domain_1_auto_routers_source_nodes_out_0_flit_0_bits_tail; // @[LazyModule.scala 353:16]
  assign router_sink_domain_auto_routers_dest_nodes_in_0_flit_0_bits_payload =
    router_sink_domain_1_auto_routers_source_nodes_out_0_flit_0_bits_payload; // @[LazyModule.scala 353:16]
  assign router_sink_domain_auto_routers_dest_nodes_in_0_flit_0_bits_flow_ingress_node =
    router_sink_domain_1_auto_routers_source_nodes_out_0_flit_0_bits_flow_ingress_node; // @[LazyModule.scala 353:16]
  assign router_sink_domain_auto_routers_dest_nodes_in_0_flit_0_bits_flow_egress_node =
    router_sink_domain_1_auto_routers_source_nodes_out_0_flit_0_bits_flow_egress_node; // @[LazyModule.scala 353:16]
  assign router_sink_domain_auto_routers_dest_nodes_in_0_flit_0_bits_virt_channel_id =
    router_sink_domain_1_auto_routers_source_nodes_out_0_flit_0_bits_virt_channel_id; // @[LazyModule.scala 353:16]
  assign router_sink_domain_auto_clock_in_clock = io_router_clocks_0_clock; // @[Nodes.scala 1212:84 NoC.scala 147:88]
  assign router_sink_domain_auto_clock_in_reset = io_router_clocks_0_reset; // @[Nodes.scala 1212:84 NoC.scala 147:88]
  assign router_sink_domain_1_auto_routers_ingress_nodes_in_flit_valid = io_ingress_1_flit_valid; // @[Nodes.scala 1212:84 NoC.scala 145:78]
  assign router_sink_domain_1_auto_routers_ingress_nodes_in_flit_bits_head = io_ingress_1_flit_bits_head; // @[Nodes.scala 1212:84 NoC.scala 145:78]
  assign router_sink_domain_1_auto_routers_ingress_nodes_in_flit_bits_tail = io_ingress_1_flit_bits_tail; // @[Nodes.scala 1212:84 NoC.scala 145:78]
  assign router_sink_domain_1_auto_routers_ingress_nodes_in_flit_bits_payload = io_ingress_1_flit_bits_payload; // @[Nodes.scala 1212:84 NoC.scala 145:78]
  assign router_sink_domain_1_auto_routers_ingress_nodes_in_flit_bits_egress_id = io_ingress_1_flit_bits_egress_id; // @[Nodes.scala 1212:84 NoC.scala 145:78]
  assign router_sink_domain_1_auto_routers_source_nodes_out_1_credit_return =
    router_sink_domain_2_auto_routers_dest_nodes_in_0_credit_return; // @[LazyModule.scala 355:16]
  assign router_sink_domain_1_auto_routers_source_nodes_out_1_vc_free =
    router_sink_domain_2_auto_routers_dest_nodes_in_0_vc_free; // @[LazyModule.scala 355:16]
  assign router_sink_domain_1_auto_routers_source_nodes_out_0_credit_return =
    router_sink_domain_auto_routers_dest_nodes_in_0_credit_return; // @[LazyModule.scala 353:16]
  assign router_sink_domain_1_auto_routers_source_nodes_out_0_vc_free =
    router_sink_domain_auto_routers_dest_nodes_in_0_vc_free; // @[LazyModule.scala 353:16]
  assign router_sink_domain_1_auto_routers_dest_nodes_in_1_flit_0_valid =
    router_sink_domain_2_auto_routers_source_nodes_out_0_flit_0_valid; // @[LazyModule.scala 353:16]
  assign router_sink_domain_1_auto_routers_dest_nodes_in_1_flit_0_bits_head =
    router_sink_domain_2_auto_routers_source_nodes_out_0_flit_0_bits_head; // @[LazyModule.scala 353:16]
  assign router_sink_domain_1_auto_routers_dest_nodes_in_1_flit_0_bits_tail =
    router_sink_domain_2_auto_routers_source_nodes_out_0_flit_0_bits_tail; // @[LazyModule.scala 353:16]
  assign router_sink_domain_1_auto_routers_dest_nodes_in_1_flit_0_bits_payload =
    router_sink_domain_2_auto_routers_source_nodes_out_0_flit_0_bits_payload; // @[LazyModule.scala 353:16]
  assign router_sink_domain_1_auto_routers_dest_nodes_in_1_flit_0_bits_flow_ingress_node =
    router_sink_domain_2_auto_routers_source_nodes_out_0_flit_0_bits_flow_ingress_node; // @[LazyModule.scala 353:16]
  assign router_sink_domain_1_auto_routers_dest_nodes_in_1_flit_0_bits_flow_egress_node =
    router_sink_domain_2_auto_routers_source_nodes_out_0_flit_0_bits_flow_egress_node; // @[LazyModule.scala 353:16]
  assign router_sink_domain_1_auto_routers_dest_nodes_in_1_flit_0_bits_virt_channel_id =
    router_sink_domain_2_auto_routers_source_nodes_out_0_flit_0_bits_virt_channel_id; // @[LazyModule.scala 353:16]
  assign router_sink_domain_1_auto_routers_dest_nodes_in_0_flit_0_valid =
    router_sink_domain_auto_routers_source_nodes_out_0_flit_0_valid; // @[LazyModule.scala 355:16]
  assign router_sink_domain_1_auto_routers_dest_nodes_in_0_flit_0_bits_head =
    router_sink_domain_auto_routers_source_nodes_out_0_flit_0_bits_head; // @[LazyModule.scala 355:16]
  assign router_sink_domain_1_auto_routers_dest_nodes_in_0_flit_0_bits_tail =
    router_sink_domain_auto_routers_source_nodes_out_0_flit_0_bits_tail; // @[LazyModule.scala 355:16]
  assign router_sink_domain_1_auto_routers_dest_nodes_in_0_flit_0_bits_payload =
    router_sink_domain_auto_routers_source_nodes_out_0_flit_0_bits_payload; // @[LazyModule.scala 355:16]
  assign router_sink_domain_1_auto_routers_dest_nodes_in_0_flit_0_bits_flow_ingress_node =
    router_sink_domain_auto_routers_source_nodes_out_0_flit_0_bits_flow_ingress_node; // @[LazyModule.scala 355:16]
  assign router_sink_domain_1_auto_routers_dest_nodes_in_0_flit_0_bits_flow_egress_node =
    router_sink_domain_auto_routers_source_nodes_out_0_flit_0_bits_flow_egress_node; // @[LazyModule.scala 355:16]
  assign router_sink_domain_1_auto_routers_dest_nodes_in_0_flit_0_bits_virt_channel_id =
    router_sink_domain_auto_routers_source_nodes_out_0_flit_0_bits_virt_channel_id; // @[LazyModule.scala 355:16]
  assign router_sink_domain_1_auto_clock_in_clock = io_router_clocks_1_clock; // @[Nodes.scala 1212:84 NoC.scala 147:88]
  assign router_sink_domain_1_auto_clock_in_reset = io_router_clocks_1_reset; // @[Nodes.scala 1212:84 NoC.scala 147:88]
  assign router_sink_domain_2_auto_routers_ingress_nodes_in_flit_valid = io_ingress_2_flit_valid; // @[Nodes.scala 1212:84 NoC.scala 145:78]
  assign router_sink_domain_2_auto_routers_ingress_nodes_in_flit_bits_head = io_ingress_2_flit_bits_head; // @[Nodes.scala 1212:84 NoC.scala 145:78]
  assign router_sink_domain_2_auto_routers_ingress_nodes_in_flit_bits_tail = io_ingress_2_flit_bits_tail; // @[Nodes.scala 1212:84 NoC.scala 145:78]
  assign router_sink_domain_2_auto_routers_ingress_nodes_in_flit_bits_payload = io_ingress_2_flit_bits_payload; // @[Nodes.scala 1212:84 NoC.scala 145:78]
  assign router_sink_domain_2_auto_routers_ingress_nodes_in_flit_bits_egress_id = io_ingress_2_flit_bits_egress_id; // @[Nodes.scala 1212:84 NoC.scala 145:78]
  assign router_sink_domain_2_auto_routers_source_nodes_out_1_credit_return =
    router_sink_domain_3_auto_routers_dest_nodes_in_1_credit_return; // @[LazyModule.scala 355:16]
  assign router_sink_domain_2_auto_routers_source_nodes_out_1_vc_free =
    router_sink_domain_3_auto_routers_dest_nodes_in_1_vc_free; // @[LazyModule.scala 355:16]
  assign router_sink_domain_2_auto_routers_source_nodes_out_0_credit_return =
    router_sink_domain_1_auto_routers_dest_nodes_in_1_credit_return; // @[LazyModule.scala 353:16]
  assign router_sink_domain_2_auto_routers_source_nodes_out_0_vc_free =
    router_sink_domain_1_auto_routers_dest_nodes_in_1_vc_free; // @[LazyModule.scala 353:16]
  assign router_sink_domain_2_auto_routers_dest_nodes_in_1_flit_0_valid =
    router_sink_domain_3_auto_routers_source_nodes_out_1_flit_0_valid; // @[LazyModule.scala 353:16]
  assign router_sink_domain_2_auto_routers_dest_nodes_in_1_flit_0_bits_head =
    router_sink_domain_3_auto_routers_source_nodes_out_1_flit_0_bits_head; // @[LazyModule.scala 353:16]
  assign router_sink_domain_2_auto_routers_dest_nodes_in_1_flit_0_bits_tail =
    router_sink_domain_3_auto_routers_source_nodes_out_1_flit_0_bits_tail; // @[LazyModule.scala 353:16]
  assign router_sink_domain_2_auto_routers_dest_nodes_in_1_flit_0_bits_payload =
    router_sink_domain_3_auto_routers_source_nodes_out_1_flit_0_bits_payload; // @[LazyModule.scala 353:16]
  assign router_sink_domain_2_auto_routers_dest_nodes_in_1_flit_0_bits_flow_ingress_node =
    router_sink_domain_3_auto_routers_source_nodes_out_1_flit_0_bits_flow_ingress_node; // @[LazyModule.scala 353:16]
  assign router_sink_domain_2_auto_routers_dest_nodes_in_1_flit_0_bits_flow_egress_node =
    router_sink_domain_3_auto_routers_source_nodes_out_1_flit_0_bits_flow_egress_node; // @[LazyModule.scala 353:16]
  assign router_sink_domain_2_auto_routers_dest_nodes_in_1_flit_0_bits_virt_channel_id =
    router_sink_domain_3_auto_routers_source_nodes_out_1_flit_0_bits_virt_channel_id; // @[LazyModule.scala 353:16]
  assign router_sink_domain_2_auto_routers_dest_nodes_in_0_flit_0_valid =
    router_sink_domain_1_auto_routers_source_nodes_out_1_flit_0_valid; // @[LazyModule.scala 355:16]
  assign router_sink_domain_2_auto_routers_dest_nodes_in_0_flit_0_bits_head =
    router_sink_domain_1_auto_routers_source_nodes_out_1_flit_0_bits_head; // @[LazyModule.scala 355:16]
  assign router_sink_domain_2_auto_routers_dest_nodes_in_0_flit_0_bits_tail =
    router_sink_domain_1_auto_routers_source_nodes_out_1_flit_0_bits_tail; // @[LazyModule.scala 355:16]
  assign router_sink_domain_2_auto_routers_dest_nodes_in_0_flit_0_bits_payload =
    router_sink_domain_1_auto_routers_source_nodes_out_1_flit_0_bits_payload; // @[LazyModule.scala 355:16]
  assign router_sink_domain_2_auto_routers_dest_nodes_in_0_flit_0_bits_flow_ingress_node =
    router_sink_domain_1_auto_routers_source_nodes_out_1_flit_0_bits_flow_ingress_node; // @[LazyModule.scala 355:16]
  assign router_sink_domain_2_auto_routers_dest_nodes_in_0_flit_0_bits_flow_egress_node =
    router_sink_domain_1_auto_routers_source_nodes_out_1_flit_0_bits_flow_egress_node; // @[LazyModule.scala 355:16]
  assign router_sink_domain_2_auto_routers_dest_nodes_in_0_flit_0_bits_virt_channel_id =
    router_sink_domain_1_auto_routers_source_nodes_out_1_flit_0_bits_virt_channel_id; // @[LazyModule.scala 355:16]
  assign router_sink_domain_2_auto_clock_in_clock = io_router_clocks_2_clock; // @[Nodes.scala 1212:84 NoC.scala 147:88]
  assign router_sink_domain_2_auto_clock_in_reset = io_router_clocks_2_reset; // @[Nodes.scala 1212:84 NoC.scala 147:88]
  assign router_sink_domain_3_auto_routers_ingress_nodes_in_flit_valid = io_ingress_3_flit_valid; // @[Nodes.scala 1212:84 NoC.scala 145:78]
  assign router_sink_domain_3_auto_routers_ingress_nodes_in_flit_bits_head = io_ingress_3_flit_bits_head; // @[Nodes.scala 1212:84 NoC.scala 145:78]
  assign router_sink_domain_3_auto_routers_ingress_nodes_in_flit_bits_tail = io_ingress_3_flit_bits_tail; // @[Nodes.scala 1212:84 NoC.scala 145:78]
  assign router_sink_domain_3_auto_routers_ingress_nodes_in_flit_bits_payload = io_ingress_3_flit_bits_payload; // @[Nodes.scala 1212:84 NoC.scala 145:78]
  assign router_sink_domain_3_auto_routers_ingress_nodes_in_flit_bits_egress_id = io_ingress_3_flit_bits_egress_id; // @[Nodes.scala 1212:84 NoC.scala 145:78]
  assign router_sink_domain_3_auto_routers_source_nodes_out_1_credit_return =
    router_sink_domain_2_auto_routers_dest_nodes_in_1_credit_return; // @[LazyModule.scala 353:16]
  assign router_sink_domain_3_auto_routers_source_nodes_out_1_vc_free =
    router_sink_domain_2_auto_routers_dest_nodes_in_1_vc_free; // @[LazyModule.scala 353:16]
  assign router_sink_domain_3_auto_routers_source_nodes_out_0_credit_return =
    router_sink_domain_auto_routers_dest_nodes_in_1_credit_return; // @[LazyModule.scala 353:16]
  assign router_sink_domain_3_auto_routers_source_nodes_out_0_vc_free =
    router_sink_domain_auto_routers_dest_nodes_in_1_vc_free; // @[LazyModule.scala 353:16]
  assign router_sink_domain_3_auto_routers_dest_nodes_in_1_flit_0_valid =
    router_sink_domain_2_auto_routers_source_nodes_out_1_flit_0_valid; // @[LazyModule.scala 355:16]
  assign router_sink_domain_3_auto_routers_dest_nodes_in_1_flit_0_bits_head =
    router_sink_domain_2_auto_routers_source_nodes_out_1_flit_0_bits_head; // @[LazyModule.scala 355:16]
  assign router_sink_domain_3_auto_routers_dest_nodes_in_1_flit_0_bits_tail =
    router_sink_domain_2_auto_routers_source_nodes_out_1_flit_0_bits_tail; // @[LazyModule.scala 355:16]
  assign router_sink_domain_3_auto_routers_dest_nodes_in_1_flit_0_bits_payload =
    router_sink_domain_2_auto_routers_source_nodes_out_1_flit_0_bits_payload; // @[LazyModule.scala 355:16]
  assign router_sink_domain_3_auto_routers_dest_nodes_in_1_flit_0_bits_flow_ingress_node =
    router_sink_domain_2_auto_routers_source_nodes_out_1_flit_0_bits_flow_ingress_node; // @[LazyModule.scala 355:16]
  assign router_sink_domain_3_auto_routers_dest_nodes_in_1_flit_0_bits_flow_egress_node =
    router_sink_domain_2_auto_routers_source_nodes_out_1_flit_0_bits_flow_egress_node; // @[LazyModule.scala 355:16]
  assign router_sink_domain_3_auto_routers_dest_nodes_in_1_flit_0_bits_virt_channel_id =
    router_sink_domain_2_auto_routers_source_nodes_out_1_flit_0_bits_virt_channel_id; // @[LazyModule.scala 355:16]
  assign router_sink_domain_3_auto_routers_dest_nodes_in_0_flit_0_valid =
    router_sink_domain_auto_routers_source_nodes_out_1_flit_0_valid; // @[LazyModule.scala 355:16]
  assign router_sink_domain_3_auto_routers_dest_nodes_in_0_flit_0_bits_head =
    router_sink_domain_auto_routers_source_nodes_out_1_flit_0_bits_head; // @[LazyModule.scala 355:16]
  assign router_sink_domain_3_auto_routers_dest_nodes_in_0_flit_0_bits_tail =
    router_sink_domain_auto_routers_source_nodes_out_1_flit_0_bits_tail; // @[LazyModule.scala 355:16]
  assign router_sink_domain_3_auto_routers_dest_nodes_in_0_flit_0_bits_payload =
    router_sink_domain_auto_routers_source_nodes_out_1_flit_0_bits_payload; // @[LazyModule.scala 355:16]
  assign router_sink_domain_3_auto_routers_dest_nodes_in_0_flit_0_bits_flow_ingress_node =
    router_sink_domain_auto_routers_source_nodes_out_1_flit_0_bits_flow_ingress_node; // @[LazyModule.scala 355:16]
  assign router_sink_domain_3_auto_routers_dest_nodes_in_0_flit_0_bits_flow_egress_node =
    router_sink_domain_auto_routers_source_nodes_out_1_flit_0_bits_flow_egress_node; // @[LazyModule.scala 355:16]
  assign router_sink_domain_3_auto_routers_dest_nodes_in_0_flit_0_bits_virt_channel_id =
    router_sink_domain_auto_routers_source_nodes_out_1_flit_0_bits_virt_channel_id; // @[LazyModule.scala 355:16]
  assign router_sink_domain_3_auto_clock_in_clock = io_router_clocks_3_clock; // @[Nodes.scala 1212:84 NoC.scala 147:88]
  assign router_sink_domain_3_auto_clock_in_reset = io_router_clocks_3_reset; // @[Nodes.scala 1212:84 NoC.scala 147:88]
  always @(posedge clock) begin
    if (reset) begin // @[NoC.scala 160:37]
      debug_va_stall_ctr <= 64'h0; // @[NoC.scala 160:37]
    end else begin
      debug_va_stall_ctr <= _debug_va_stall_ctr_T_23; // @[NoC.scala 163:24]
    end
    if (reset) begin // @[NoC.scala 161:37]
      debug_sa_stall_ctr <= 64'h0; // @[NoC.scala 161:37]
    end else begin
      debug_sa_stall_ctr <= _debug_sa_stall_ctr_T_23; // @[NoC.scala 164:24]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  debug_va_stall_ctr = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  debug_sa_stall_ctr = _RAND_1[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MaxPeriodFibonacciLFSR(
  input   clock,
  input   reset,
  output  io_out_0,
  output  io_out_1,
  output  io_out_2,
  output  io_out_3,
  output  io_out_4,
  output  io_out_5,
  output  io_out_6,
  output  io_out_7,
  output  io_out_8,
  output  io_out_9,
  output  io_out_10,
  output  io_out_11,
  output  io_out_12,
  output  io_out_13,
  output  io_out_14,
  output  io_out_15,
  output  io_out_16,
  output  io_out_17,
  output  io_out_18,
  output  io_out_19
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
`endif // RANDOMIZE_REG_INIT
  reg  state_0; // @[PRNG.scala 55:49]
  reg  state_1; // @[PRNG.scala 55:49]
  reg  state_2; // @[PRNG.scala 55:49]
  reg  state_3; // @[PRNG.scala 55:49]
  reg  state_4; // @[PRNG.scala 55:49]
  reg  state_5; // @[PRNG.scala 55:49]
  reg  state_6; // @[PRNG.scala 55:49]
  reg  state_7; // @[PRNG.scala 55:49]
  reg  state_8; // @[PRNG.scala 55:49]
  reg  state_9; // @[PRNG.scala 55:49]
  reg  state_10; // @[PRNG.scala 55:49]
  reg  state_11; // @[PRNG.scala 55:49]
  reg  state_12; // @[PRNG.scala 55:49]
  reg  state_13; // @[PRNG.scala 55:49]
  reg  state_14; // @[PRNG.scala 55:49]
  reg  state_15; // @[PRNG.scala 55:49]
  reg  state_16; // @[PRNG.scala 55:49]
  reg  state_17; // @[PRNG.scala 55:49]
  reg  state_18; // @[PRNG.scala 55:49]
  reg  state_19; // @[PRNG.scala 55:49]
  wire  _T = state_19 ^ state_16; // @[LFSR.scala 15:41]
  assign io_out_0 = state_0; // @[PRNG.scala 78:10]
  assign io_out_1 = state_1; // @[PRNG.scala 78:10]
  assign io_out_2 = state_2; // @[PRNG.scala 78:10]
  assign io_out_3 = state_3; // @[PRNG.scala 78:10]
  assign io_out_4 = state_4; // @[PRNG.scala 78:10]
  assign io_out_5 = state_5; // @[PRNG.scala 78:10]
  assign io_out_6 = state_6; // @[PRNG.scala 78:10]
  assign io_out_7 = state_7; // @[PRNG.scala 78:10]
  assign io_out_8 = state_8; // @[PRNG.scala 78:10]
  assign io_out_9 = state_9; // @[PRNG.scala 78:10]
  assign io_out_10 = state_10; // @[PRNG.scala 78:10]
  assign io_out_11 = state_11; // @[PRNG.scala 78:10]
  assign io_out_12 = state_12; // @[PRNG.scala 78:10]
  assign io_out_13 = state_13; // @[PRNG.scala 78:10]
  assign io_out_14 = state_14; // @[PRNG.scala 78:10]
  assign io_out_15 = state_15; // @[PRNG.scala 78:10]
  assign io_out_16 = state_16; // @[PRNG.scala 78:10]
  assign io_out_17 = state_17; // @[PRNG.scala 78:10]
  assign io_out_18 = state_18; // @[PRNG.scala 78:10]
  assign io_out_19 = state_19; // @[PRNG.scala 78:10]
  always @(posedge clock) begin
    state_0 <= reset | _T; // @[PRNG.scala 55:{49,49}]
    if (reset) begin // @[PRNG.scala 55:49]
      state_1 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_1 <= state_0;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_2 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_2 <= state_1;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_3 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_3 <= state_2;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_4 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_4 <= state_3;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_5 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_5 <= state_4;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_6 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_6 <= state_5;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_7 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_7 <= state_6;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_8 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_8 <= state_7;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_9 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_9 <= state_8;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_10 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_10 <= state_9;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_11 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_11 <= state_10;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_12 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_12 <= state_11;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_13 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_13 <= state_12;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_14 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_14 <= state_13;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_15 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_15 <= state_14;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_16 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_16 <= state_15;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_17 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_17 <= state_16;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_18 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_18 <= state_17;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_19 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_19 <= state_18;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  state_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  state_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  state_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  state_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  state_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  state_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  state_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  state_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  state_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  state_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  state_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  state_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  state_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  state_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  state_15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  state_16 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  state_17 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  state_18 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  state_19 = _RAND_19[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module InputGen(
  input         clock,
  input         reset,
  input         io_out_ready,
  output        io_out_valid,
  output        io_out_bits_head,
  output        io_out_bits_tail,
  output [63:0] io_out_bits_payload,
  output [1:0]  io_out_bits_egress_id,
  input         io_rob_ready,
  input  [6:0]  io_rob_idx,
  input  [31:0] io_tsc,
  output        io_fire,
  output [3:0]  io_n_flits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  packet_remaining_prng_clock; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_reset; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_0; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_1; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_2; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_3; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_4; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_5; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_6; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_7; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_8; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_9; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_10; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_11; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_12; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_13; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_14; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_15; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_16; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_17; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_18; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_19; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_clock; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_reset; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_0; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_1; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_2; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_3; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_4; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_5; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_6; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_7; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_8; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_9; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_10; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_11; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_12; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_13; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_14; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_15; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_16; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_17; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_18; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_19; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_clock; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_reset; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_0; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_1; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_2; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_3; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_4; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_5; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_6; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_7; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_8; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_9; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_10; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_11; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_12; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_13; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_14; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_15; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_16; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_17; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_18; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_19; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_clock; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_reset; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_0; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_1; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_2; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_3; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_4; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_5; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_6; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_7; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_8; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_9; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_10; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_11; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_12; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_13; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_14; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_15; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_16; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_17; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_18; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_19; // @[PRNG.scala 91:22]
  reg [3:0] flits_left; // @[TestHarness.scala 71:27]
  reg [3:0] flits_fired; // @[TestHarness.scala 72:28]
  reg [1:0] egress; // @[TestHarness.scala 73:19]
  reg [31:0] payload_tsc; // @[TestHarness.scala 74:20]
  reg [15:0] payload_rob_idx; // @[TestHarness.scala 74:20]
  wire  can_fire = flits_left == 4'h0 & io_rob_ready; // @[TestHarness.scala 76:39]
  wire [9:0] packet_remaining_lo = {packet_remaining_prng_io_out_9,packet_remaining_prng_io_out_8,
    packet_remaining_prng_io_out_7,packet_remaining_prng_io_out_6,packet_remaining_prng_io_out_5,
    packet_remaining_prng_io_out_4,packet_remaining_prng_io_out_3,packet_remaining_prng_io_out_2,
    packet_remaining_prng_io_out_1,packet_remaining_prng_io_out_0}; // @[PRNG.scala 95:17]
  wire [9:0] packet_remaining_hi = {packet_remaining_prng_io_out_19,packet_remaining_prng_io_out_18,
    packet_remaining_prng_io_out_17,packet_remaining_prng_io_out_16,packet_remaining_prng_io_out_15,
    packet_remaining_prng_io_out_14,packet_remaining_prng_io_out_13,packet_remaining_prng_io_out_12,
    packet_remaining_prng_io_out_11,packet_remaining_prng_io_out_10}; // @[PRNG.scala 95:17]
  wire [19:0] _packet_remaining_T = {packet_remaining_hi,packet_remaining_lo}; // @[PRNG.scala 95:17]
  wire [19:0] _GEN_0 = _packet_remaining_T % 20'h8; // @[TestHarness.scala 78:89]
  wire [3:0] packet_remaining = _GEN_0[3:0]; // @[TestHarness.scala 78:89]
  wire [9:0] io_out_bits_egress_id_lo = {io_out_bits_egress_id_prng_io_out_9,io_out_bits_egress_id_prng_io_out_8,
    io_out_bits_egress_id_prng_io_out_7,io_out_bits_egress_id_prng_io_out_6,io_out_bits_egress_id_prng_io_out_5,
    io_out_bits_egress_id_prng_io_out_4,io_out_bits_egress_id_prng_io_out_3,io_out_bits_egress_id_prng_io_out_2,
    io_out_bits_egress_id_prng_io_out_1,io_out_bits_egress_id_prng_io_out_0}; // @[PRNG.scala 95:17]
  wire [9:0] io_out_bits_egress_id_hi = {io_out_bits_egress_id_prng_io_out_19,io_out_bits_egress_id_prng_io_out_18,
    io_out_bits_egress_id_prng_io_out_17,io_out_bits_egress_id_prng_io_out_16,io_out_bits_egress_id_prng_io_out_15,
    io_out_bits_egress_id_prng_io_out_14,io_out_bits_egress_id_prng_io_out_13,io_out_bits_egress_id_prng_io_out_12,
    io_out_bits_egress_id_prng_io_out_11,io_out_bits_egress_id_prng_io_out_10}; // @[PRNG.scala 95:17]
  wire [19:0] _io_out_bits_egress_id_T = {io_out_bits_egress_id_hi,io_out_bits_egress_id_lo}; // @[PRNG.scala 95:17]
  wire [19:0] _GEN_5 = _io_out_bits_egress_id_T % 20'h4; // @[TestHarness.scala 84:92]
  wire [1:0] _GEN_1 = 2'h1 == _GEN_5[1:0] ? 2'h1 : 2'h0; // @[TestHarness.scala 84:{25,25}]
  wire [1:0] _GEN_2 = 2'h2 == _GEN_5[1:0] ? 2'h2 : _GEN_1; // @[TestHarness.scala 84:{25,25}]
  wire [1:0] _GEN_3 = 2'h3 == _GEN_5[1:0] ? 2'h3 : _GEN_2; // @[TestHarness.scala 84:{25,25}]
  wire [31:0] out_payload_tsc = flits_left != 4'h0 ? payload_tsc : io_tsc; // @[TestHarness.scala 100:29 105:17 87:19]
  wire [15:0] out_payload_rob_idx = flits_left != 4'h0 ? payload_rob_idx : {{9'd0}, io_rob_idx}; // @[TestHarness.scala 100:29 105:17 88:23]
  wire [47:0] io_out_bits_payload_hi = {out_payload_tsc,out_payload_rob_idx}; // @[TestHarness.scala 86:38]
  wire [3:0] _GEN_18 = flits_left != 4'h0 ? flits_fired : 4'h0; // @[TestHarness.scala 100:29 106:29 89:27]
  wire [15:0] out_payload_flits_fired = {{12'd0}, _GEN_18}; // @[TestHarness.scala 85:25]
  wire  _io_fire_T = io_out_ready & io_out_valid; // @[Decoupled.scala 51:35]
  wire [3:0] _GEN_4 = io_fire & ~io_out_bits_tail ? packet_remaining : flits_left; // @[TestHarness.scala 94:39 95:16 71:27]
  wire [3:0] _GEN_9 = io_fire & ~io_out_bits_tail ? 4'h1 : flits_fired; // @[TestHarness.scala 94:39 98:17 72:28]
  wire [3:0] _flits_fired_T_1 = flits_fired + 4'h1; // @[TestHarness.scala 109:34]
  wire [3:0] _flits_left_T_1 = flits_left - 4'h1; // @[TestHarness.scala 110:32]
  MaxPeriodFibonacciLFSR packet_remaining_prng ( // @[PRNG.scala 91:22]
    .clock(packet_remaining_prng_clock),
    .reset(packet_remaining_prng_reset),
    .io_out_0(packet_remaining_prng_io_out_0),
    .io_out_1(packet_remaining_prng_io_out_1),
    .io_out_2(packet_remaining_prng_io_out_2),
    .io_out_3(packet_remaining_prng_io_out_3),
    .io_out_4(packet_remaining_prng_io_out_4),
    .io_out_5(packet_remaining_prng_io_out_5),
    .io_out_6(packet_remaining_prng_io_out_6),
    .io_out_7(packet_remaining_prng_io_out_7),
    .io_out_8(packet_remaining_prng_io_out_8),
    .io_out_9(packet_remaining_prng_io_out_9),
    .io_out_10(packet_remaining_prng_io_out_10),
    .io_out_11(packet_remaining_prng_io_out_11),
    .io_out_12(packet_remaining_prng_io_out_12),
    .io_out_13(packet_remaining_prng_io_out_13),
    .io_out_14(packet_remaining_prng_io_out_14),
    .io_out_15(packet_remaining_prng_io_out_15),
    .io_out_16(packet_remaining_prng_io_out_16),
    .io_out_17(packet_remaining_prng_io_out_17),
    .io_out_18(packet_remaining_prng_io_out_18),
    .io_out_19(packet_remaining_prng_io_out_19)
  );
  MaxPeriodFibonacciLFSR random_flit_delay_prng ( // @[PRNG.scala 91:22]
    .clock(random_flit_delay_prng_clock),
    .reset(random_flit_delay_prng_reset),
    .io_out_0(random_flit_delay_prng_io_out_0),
    .io_out_1(random_flit_delay_prng_io_out_1),
    .io_out_2(random_flit_delay_prng_io_out_2),
    .io_out_3(random_flit_delay_prng_io_out_3),
    .io_out_4(random_flit_delay_prng_io_out_4),
    .io_out_5(random_flit_delay_prng_io_out_5),
    .io_out_6(random_flit_delay_prng_io_out_6),
    .io_out_7(random_flit_delay_prng_io_out_7),
    .io_out_8(random_flit_delay_prng_io_out_8),
    .io_out_9(random_flit_delay_prng_io_out_9),
    .io_out_10(random_flit_delay_prng_io_out_10),
    .io_out_11(random_flit_delay_prng_io_out_11),
    .io_out_12(random_flit_delay_prng_io_out_12),
    .io_out_13(random_flit_delay_prng_io_out_13),
    .io_out_14(random_flit_delay_prng_io_out_14),
    .io_out_15(random_flit_delay_prng_io_out_15),
    .io_out_16(random_flit_delay_prng_io_out_16),
    .io_out_17(random_flit_delay_prng_io_out_17),
    .io_out_18(random_flit_delay_prng_io_out_18),
    .io_out_19(random_flit_delay_prng_io_out_19)
  );
  MaxPeriodFibonacciLFSR random_packet_delay_prng ( // @[PRNG.scala 91:22]
    .clock(random_packet_delay_prng_clock),
    .reset(random_packet_delay_prng_reset),
    .io_out_0(random_packet_delay_prng_io_out_0),
    .io_out_1(random_packet_delay_prng_io_out_1),
    .io_out_2(random_packet_delay_prng_io_out_2),
    .io_out_3(random_packet_delay_prng_io_out_3),
    .io_out_4(random_packet_delay_prng_io_out_4),
    .io_out_5(random_packet_delay_prng_io_out_5),
    .io_out_6(random_packet_delay_prng_io_out_6),
    .io_out_7(random_packet_delay_prng_io_out_7),
    .io_out_8(random_packet_delay_prng_io_out_8),
    .io_out_9(random_packet_delay_prng_io_out_9),
    .io_out_10(random_packet_delay_prng_io_out_10),
    .io_out_11(random_packet_delay_prng_io_out_11),
    .io_out_12(random_packet_delay_prng_io_out_12),
    .io_out_13(random_packet_delay_prng_io_out_13),
    .io_out_14(random_packet_delay_prng_io_out_14),
    .io_out_15(random_packet_delay_prng_io_out_15),
    .io_out_16(random_packet_delay_prng_io_out_16),
    .io_out_17(random_packet_delay_prng_io_out_17),
    .io_out_18(random_packet_delay_prng_io_out_18),
    .io_out_19(random_packet_delay_prng_io_out_19)
  );
  MaxPeriodFibonacciLFSR io_out_bits_egress_id_prng ( // @[PRNG.scala 91:22]
    .clock(io_out_bits_egress_id_prng_clock),
    .reset(io_out_bits_egress_id_prng_reset),
    .io_out_0(io_out_bits_egress_id_prng_io_out_0),
    .io_out_1(io_out_bits_egress_id_prng_io_out_1),
    .io_out_2(io_out_bits_egress_id_prng_io_out_2),
    .io_out_3(io_out_bits_egress_id_prng_io_out_3),
    .io_out_4(io_out_bits_egress_id_prng_io_out_4),
    .io_out_5(io_out_bits_egress_id_prng_io_out_5),
    .io_out_6(io_out_bits_egress_id_prng_io_out_6),
    .io_out_7(io_out_bits_egress_id_prng_io_out_7),
    .io_out_8(io_out_bits_egress_id_prng_io_out_8),
    .io_out_9(io_out_bits_egress_id_prng_io_out_9),
    .io_out_10(io_out_bits_egress_id_prng_io_out_10),
    .io_out_11(io_out_bits_egress_id_prng_io_out_11),
    .io_out_12(io_out_bits_egress_id_prng_io_out_12),
    .io_out_13(io_out_bits_egress_id_prng_io_out_13),
    .io_out_14(io_out_bits_egress_id_prng_io_out_14),
    .io_out_15(io_out_bits_egress_id_prng_io_out_15),
    .io_out_16(io_out_bits_egress_id_prng_io_out_16),
    .io_out_17(io_out_bits_egress_id_prng_io_out_17),
    .io_out_18(io_out_bits_egress_id_prng_io_out_18),
    .io_out_19(io_out_bits_egress_id_prng_io_out_19)
  );
  assign io_out_valid = flits_left != 4'h0 | can_fire; // @[TestHarness.scala 100:29 101:18 81:16]
  assign io_out_bits_head = flits_left != 4'h0 ? 1'h0 : 1'h1; // @[TestHarness.scala 100:29 102:22 82:20]
  assign io_out_bits_tail = flits_left != 4'h0 ? flits_left == 4'h1 : packet_remaining == 4'h0; // @[TestHarness.scala 100:29 103:22 83:20]
  assign io_out_bits_payload = {io_out_bits_payload_hi,out_payload_flits_fired}; // @[TestHarness.scala 86:38]
  assign io_out_bits_egress_id = flits_left != 4'h0 ? egress : _GEN_3; // @[TestHarness.scala 100:29 104:27 84:25]
  assign io_fire = can_fire & _io_fire_T; // @[TestHarness.scala 92:23]
  assign io_n_flits = packet_remaining + 4'h1; // @[TestHarness.scala 91:34]
  assign packet_remaining_prng_clock = clock;
  assign packet_remaining_prng_reset = reset;
  assign random_flit_delay_prng_clock = clock;
  assign random_flit_delay_prng_reset = reset;
  assign random_packet_delay_prng_clock = clock;
  assign random_packet_delay_prng_reset = reset;
  assign io_out_bits_egress_id_prng_clock = clock;
  assign io_out_bits_egress_id_prng_reset = reset;
  always @(posedge clock) begin
    if (reset) begin // @[TestHarness.scala 71:27]
      flits_left <= 4'h0; // @[TestHarness.scala 71:27]
    end else if (flits_left != 4'h0) begin // @[TestHarness.scala 100:29]
      if (_io_fire_T) begin // @[TestHarness.scala 108:26]
        flits_left <= _flits_left_T_1; // @[TestHarness.scala 110:18]
      end else begin
        flits_left <= _GEN_4;
      end
    end else begin
      flits_left <= _GEN_4;
    end
    if (reset) begin // @[TestHarness.scala 72:28]
      flits_fired <= 4'h0; // @[TestHarness.scala 72:28]
    end else if (flits_left != 4'h0) begin // @[TestHarness.scala 100:29]
      if (_io_fire_T) begin // @[TestHarness.scala 108:26]
        flits_fired <= _flits_fired_T_1; // @[TestHarness.scala 109:19]
      end else begin
        flits_fired <= _GEN_9;
      end
    end else begin
      flits_fired <= _GEN_9;
    end
    if (io_fire & ~io_out_bits_tail) begin // @[TestHarness.scala 94:39]
      egress <= io_out_bits_egress_id; // @[TestHarness.scala 97:12]
    end
    if (io_fire & ~io_out_bits_tail) begin // @[TestHarness.scala 94:39]
      if (!(flits_left != 4'h0)) begin // @[TestHarness.scala 100:29]
        payload_tsc <= io_tsc; // @[TestHarness.scala 87:19]
      end
    end
    if (io_fire & ~io_out_bits_tail) begin // @[TestHarness.scala 94:39]
      if (!(flits_left != 4'h0)) begin // @[TestHarness.scala 100:29]
        payload_rob_idx <= {{9'd0}, io_rob_idx}; // @[TestHarness.scala 88:23]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  flits_left = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  flits_fired = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  egress = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  payload_tsc = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  payload_rob_idx = _RAND_4[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_52(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_head,
  input         io_enq_bits_tail,
  input  [63:0] io_enq_bits_payload,
  input  [1:0]  io_enq_bits_egress_id,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_head,
  output        io_deq_bits_tail,
  output [63:0] io_deq_bits_payload,
  output [1:0]  io_deq_bits_egress_id
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg  ram_head [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_head_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_head_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_head_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_tail [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_tail_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_tail_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_tail_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_en; // @[Decoupled.scala 273:95]
  reg [63:0] ram_payload [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_payload_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_payload_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [63:0] ram_payload_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [63:0] ram_payload_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_payload_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_payload_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_payload_MPORT_en; // @[Decoupled.scala 273:95]
  reg [1:0] ram_egress_id [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_egress_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_egress_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [1:0] ram_egress_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_egress_id_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_egress_id_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_egress_id_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_egress_id_MPORT_en; // @[Decoupled.scala 273:95]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 278:28]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  wire  _GEN_12 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 318:26 280:27 318:35]
  wire  do_enq = empty ? _GEN_12 : _do_enq_T; // @[Decoupled.scala 315:17 280:27]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 315:17 317:14 281:27]
  assign ram_head_io_deq_bits_MPORT_en = 1'h1;
  assign ram_head_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_head_io_deq_bits_MPORT_data = ram_head[ram_head_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_head_MPORT_data = io_enq_bits_head;
  assign ram_head_MPORT_addr = 1'h0;
  assign ram_head_MPORT_mask = 1'h1;
  assign ram_head_MPORT_en = empty ? _GEN_12 : _do_enq_T;
  assign ram_tail_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tail_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tail_io_deq_bits_MPORT_data = ram_tail[ram_tail_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_tail_MPORT_data = io_enq_bits_tail;
  assign ram_tail_MPORT_addr = 1'h0;
  assign ram_tail_MPORT_mask = 1'h1;
  assign ram_tail_MPORT_en = empty ? _GEN_12 : _do_enq_T;
  assign ram_payload_io_deq_bits_MPORT_en = 1'h1;
  assign ram_payload_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_payload_io_deq_bits_MPORT_data = ram_payload[ram_payload_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_payload_MPORT_data = io_enq_bits_payload;
  assign ram_payload_MPORT_addr = 1'h0;
  assign ram_payload_MPORT_mask = 1'h1;
  assign ram_payload_MPORT_en = empty ? _GEN_12 : _do_enq_T;
  assign ram_egress_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_egress_id_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_egress_id_io_deq_bits_MPORT_data = ram_egress_id[ram_egress_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_egress_id_MPORT_data = io_enq_bits_egress_id;
  assign ram_egress_id_MPORT_addr = 1'h0;
  assign ram_egress_id_MPORT_mask = 1'h1;
  assign ram_egress_id_MPORT_en = empty ? _GEN_12 : _do_enq_T;
  assign io_enq_ready = io_deq_ready | empty; // @[Decoupled.scala 303:16 323:{24,39}]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 302:16 314:{24,39}]
  assign io_deq_bits_head = empty ? io_enq_bits_head : ram_head_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_tail = empty ? io_enq_bits_tail : ram_tail_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_payload = empty ? io_enq_bits_payload : ram_payload_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_egress_id = empty ? io_enq_bits_egress_id : ram_egress_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  always @(posedge clock) begin
    if (ram_head_MPORT_en & ram_head_MPORT_mask) begin
      ram_head[ram_head_MPORT_addr] <= ram_head_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_tail_MPORT_en & ram_tail_MPORT_mask) begin
      ram_tail[ram_tail_MPORT_addr] <= ram_tail_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_payload_MPORT_en & ram_payload_MPORT_mask) begin
      ram_payload[ram_payload_MPORT_addr] <= ram_payload_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_egress_id_MPORT_en & ram_egress_id_MPORT_mask) begin
      ram_egress_id[ram_egress_id_MPORT_addr] <= ram_egress_id_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      if (empty) begin // @[Decoupled.scala 315:17]
        if (io_deq_ready) begin // @[Decoupled.scala 318:26]
          maybe_full <= 1'h0; // @[Decoupled.scala 318:35]
        end else begin
          maybe_full <= _do_enq_T; // @[Decoupled.scala 280:27]
        end
      end else begin
        maybe_full <= _do_enq_T; // @[Decoupled.scala 280:27]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_head[initvar] = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tail[initvar] = _RAND_1[0:0];
  _RAND_2 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload[initvar] = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_egress_id[initvar] = _RAND_3[1:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  maybe_full = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module NoCTester(
  input         clock,
  input         reset,
  input         io_to_noc_3_flit_ready,
  output        io_to_noc_3_flit_valid,
  output        io_to_noc_3_flit_bits_head,
  output        io_to_noc_3_flit_bits_tail,
  output [63:0] io_to_noc_3_flit_bits_payload,
  output [1:0]  io_to_noc_3_flit_bits_egress_id,
  input         io_to_noc_2_flit_ready,
  output        io_to_noc_2_flit_valid,
  output        io_to_noc_2_flit_bits_head,
  output        io_to_noc_2_flit_bits_tail,
  output [63:0] io_to_noc_2_flit_bits_payload,
  output [1:0]  io_to_noc_2_flit_bits_egress_id,
  input         io_to_noc_1_flit_ready,
  output        io_to_noc_1_flit_valid,
  output        io_to_noc_1_flit_bits_head,
  output        io_to_noc_1_flit_bits_tail,
  output [63:0] io_to_noc_1_flit_bits_payload,
  output [1:0]  io_to_noc_1_flit_bits_egress_id,
  input         io_to_noc_0_flit_ready,
  output        io_to_noc_0_flit_valid,
  output        io_to_noc_0_flit_bits_head,
  output        io_to_noc_0_flit_bits_tail,
  output [63:0] io_to_noc_0_flit_bits_payload,
  output [1:0]  io_to_noc_0_flit_bits_egress_id,
  output        io_from_noc_3_flit_ready,
  input         io_from_noc_3_flit_valid,
  input         io_from_noc_3_flit_bits_head,
  input         io_from_noc_3_flit_bits_tail,
  input  [63:0] io_from_noc_3_flit_bits_payload,
  input  [1:0]  io_from_noc_3_flit_bits_ingress_id,
  output        io_from_noc_2_flit_ready,
  input         io_from_noc_2_flit_valid,
  input         io_from_noc_2_flit_bits_head,
  input         io_from_noc_2_flit_bits_tail,
  input  [63:0] io_from_noc_2_flit_bits_payload,
  input  [1:0]  io_from_noc_2_flit_bits_ingress_id,
  output        io_from_noc_1_flit_ready,
  input         io_from_noc_1_flit_valid,
  input         io_from_noc_1_flit_bits_head,
  input         io_from_noc_1_flit_bits_tail,
  input  [63:0] io_from_noc_1_flit_bits_payload,
  input  [1:0]  io_from_noc_1_flit_bits_ingress_id,
  output        io_from_noc_0_flit_ready,
  input         io_from_noc_0_flit_valid,
  input         io_from_noc_0_flit_bits_head,
  input         io_from_noc_0_flit_bits_tail,
  input  [63:0] io_from_noc_0_flit_bits_payload,
  input  [1:0]  io_from_noc_0_flit_bits_ingress_id,
  output        io_success
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [127:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [63:0] _RAND_901;
  reg [63:0] _RAND_902;
  reg [63:0] _RAND_903;
  reg [63:0] _RAND_904;
  reg [63:0] _RAND_905;
  reg [63:0] _RAND_906;
  reg [63:0] _RAND_907;
  reg [63:0] _RAND_908;
  reg [63:0] _RAND_909;
  reg [63:0] _RAND_910;
  reg [63:0] _RAND_911;
  reg [63:0] _RAND_912;
  reg [63:0] _RAND_913;
  reg [63:0] _RAND_914;
  reg [63:0] _RAND_915;
  reg [63:0] _RAND_916;
  reg [63:0] _RAND_917;
  reg [63:0] _RAND_918;
  reg [63:0] _RAND_919;
  reg [63:0] _RAND_920;
  reg [63:0] _RAND_921;
  reg [63:0] _RAND_922;
  reg [63:0] _RAND_923;
  reg [63:0] _RAND_924;
  reg [63:0] _RAND_925;
  reg [63:0] _RAND_926;
  reg [63:0] _RAND_927;
  reg [63:0] _RAND_928;
  reg [63:0] _RAND_929;
  reg [63:0] _RAND_930;
  reg [63:0] _RAND_931;
  reg [63:0] _RAND_932;
  reg [63:0] _RAND_933;
  reg [63:0] _RAND_934;
  reg [63:0] _RAND_935;
  reg [63:0] _RAND_936;
  reg [63:0] _RAND_937;
  reg [63:0] _RAND_938;
  reg [63:0] _RAND_939;
  reg [63:0] _RAND_940;
  reg [63:0] _RAND_941;
  reg [63:0] _RAND_942;
  reg [63:0] _RAND_943;
  reg [63:0] _RAND_944;
  reg [63:0] _RAND_945;
  reg [63:0] _RAND_946;
  reg [63:0] _RAND_947;
  reg [63:0] _RAND_948;
  reg [63:0] _RAND_949;
  reg [63:0] _RAND_950;
  reg [63:0] _RAND_951;
  reg [63:0] _RAND_952;
  reg [63:0] _RAND_953;
  reg [63:0] _RAND_954;
  reg [63:0] _RAND_955;
  reg [63:0] _RAND_956;
  reg [63:0] _RAND_957;
  reg [63:0] _RAND_958;
  reg [63:0] _RAND_959;
  reg [63:0] _RAND_960;
  reg [63:0] _RAND_961;
  reg [63:0] _RAND_962;
  reg [63:0] _RAND_963;
  reg [63:0] _RAND_964;
  reg [63:0] _RAND_965;
  reg [63:0] _RAND_966;
  reg [63:0] _RAND_967;
  reg [63:0] _RAND_968;
  reg [63:0] _RAND_969;
  reg [63:0] _RAND_970;
  reg [63:0] _RAND_971;
  reg [63:0] _RAND_972;
  reg [63:0] _RAND_973;
  reg [63:0] _RAND_974;
  reg [63:0] _RAND_975;
  reg [63:0] _RAND_976;
  reg [63:0] _RAND_977;
  reg [63:0] _RAND_978;
  reg [63:0] _RAND_979;
  reg [63:0] _RAND_980;
  reg [63:0] _RAND_981;
  reg [63:0] _RAND_982;
  reg [63:0] _RAND_983;
  reg [63:0] _RAND_984;
  reg [63:0] _RAND_985;
  reg [63:0] _RAND_986;
  reg [63:0] _RAND_987;
  reg [63:0] _RAND_988;
  reg [63:0] _RAND_989;
  reg [63:0] _RAND_990;
  reg [63:0] _RAND_991;
  reg [63:0] _RAND_992;
  reg [63:0] _RAND_993;
  reg [63:0] _RAND_994;
  reg [63:0] _RAND_995;
  reg [63:0] _RAND_996;
  reg [63:0] _RAND_997;
  reg [63:0] _RAND_998;
  reg [63:0] _RAND_999;
  reg [63:0] _RAND_1000;
  reg [63:0] _RAND_1001;
  reg [63:0] _RAND_1002;
  reg [63:0] _RAND_1003;
  reg [63:0] _RAND_1004;
  reg [63:0] _RAND_1005;
  reg [63:0] _RAND_1006;
  reg [63:0] _RAND_1007;
  reg [63:0] _RAND_1008;
  reg [63:0] _RAND_1009;
  reg [63:0] _RAND_1010;
  reg [63:0] _RAND_1011;
  reg [63:0] _RAND_1012;
  reg [63:0] _RAND_1013;
  reg [63:0] _RAND_1014;
  reg [63:0] _RAND_1015;
  reg [63:0] _RAND_1016;
  reg [63:0] _RAND_1017;
  reg [63:0] _RAND_1018;
  reg [63:0] _RAND_1019;
  reg [63:0] _RAND_1020;
  reg [63:0] _RAND_1021;
  reg [63:0] _RAND_1022;
  reg [63:0] _RAND_1023;
  reg [63:0] _RAND_1024;
  reg [63:0] _RAND_1025;
  reg [63:0] _RAND_1026;
  reg [63:0] _RAND_1027;
  reg [63:0] _RAND_1028;
  reg [31:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
`endif // RANDOMIZE_REG_INIT
  wire  igen_clock; // @[TestHarness.scala 171:22]
  wire  igen_reset; // @[TestHarness.scala 171:22]
  wire  igen_io_out_ready; // @[TestHarness.scala 171:22]
  wire  igen_io_out_valid; // @[TestHarness.scala 171:22]
  wire  igen_io_out_bits_head; // @[TestHarness.scala 171:22]
  wire  igen_io_out_bits_tail; // @[TestHarness.scala 171:22]
  wire [63:0] igen_io_out_bits_payload; // @[TestHarness.scala 171:22]
  wire [1:0] igen_io_out_bits_egress_id; // @[TestHarness.scala 171:22]
  wire  igen_io_rob_ready; // @[TestHarness.scala 171:22]
  wire [6:0] igen_io_rob_idx; // @[TestHarness.scala 171:22]
  wire [31:0] igen_io_tsc; // @[TestHarness.scala 171:22]
  wire  igen_io_fire; // @[TestHarness.scala 171:22]
  wire [3:0] igen_io_n_flits; // @[TestHarness.scala 171:22]
  wire  io_to_noc_0_flit_q_clock; // @[Decoupled.scala 375:21]
  wire  io_to_noc_0_flit_q_reset; // @[Decoupled.scala 375:21]
  wire  io_to_noc_0_flit_q_io_enq_ready; // @[Decoupled.scala 375:21]
  wire  io_to_noc_0_flit_q_io_enq_valid; // @[Decoupled.scala 375:21]
  wire  io_to_noc_0_flit_q_io_enq_bits_head; // @[Decoupled.scala 375:21]
  wire  io_to_noc_0_flit_q_io_enq_bits_tail; // @[Decoupled.scala 375:21]
  wire [63:0] io_to_noc_0_flit_q_io_enq_bits_payload; // @[Decoupled.scala 375:21]
  wire [1:0] io_to_noc_0_flit_q_io_enq_bits_egress_id; // @[Decoupled.scala 375:21]
  wire  io_to_noc_0_flit_q_io_deq_ready; // @[Decoupled.scala 375:21]
  wire  io_to_noc_0_flit_q_io_deq_valid; // @[Decoupled.scala 375:21]
  wire  io_to_noc_0_flit_q_io_deq_bits_head; // @[Decoupled.scala 375:21]
  wire  io_to_noc_0_flit_q_io_deq_bits_tail; // @[Decoupled.scala 375:21]
  wire [63:0] io_to_noc_0_flit_q_io_deq_bits_payload; // @[Decoupled.scala 375:21]
  wire [1:0] io_to_noc_0_flit_q_io_deq_bits_egress_id; // @[Decoupled.scala 375:21]
  wire  igen_1_clock; // @[TestHarness.scala 171:22]
  wire  igen_1_reset; // @[TestHarness.scala 171:22]
  wire  igen_1_io_out_ready; // @[TestHarness.scala 171:22]
  wire  igen_1_io_out_valid; // @[TestHarness.scala 171:22]
  wire  igen_1_io_out_bits_head; // @[TestHarness.scala 171:22]
  wire  igen_1_io_out_bits_tail; // @[TestHarness.scala 171:22]
  wire [63:0] igen_1_io_out_bits_payload; // @[TestHarness.scala 171:22]
  wire [1:0] igen_1_io_out_bits_egress_id; // @[TestHarness.scala 171:22]
  wire  igen_1_io_rob_ready; // @[TestHarness.scala 171:22]
  wire [6:0] igen_1_io_rob_idx; // @[TestHarness.scala 171:22]
  wire [31:0] igen_1_io_tsc; // @[TestHarness.scala 171:22]
  wire  igen_1_io_fire; // @[TestHarness.scala 171:22]
  wire [3:0] igen_1_io_n_flits; // @[TestHarness.scala 171:22]
  wire  io_to_noc_1_flit_q_clock; // @[Decoupled.scala 375:21]
  wire  io_to_noc_1_flit_q_reset; // @[Decoupled.scala 375:21]
  wire  io_to_noc_1_flit_q_io_enq_ready; // @[Decoupled.scala 375:21]
  wire  io_to_noc_1_flit_q_io_enq_valid; // @[Decoupled.scala 375:21]
  wire  io_to_noc_1_flit_q_io_enq_bits_head; // @[Decoupled.scala 375:21]
  wire  io_to_noc_1_flit_q_io_enq_bits_tail; // @[Decoupled.scala 375:21]
  wire [63:0] io_to_noc_1_flit_q_io_enq_bits_payload; // @[Decoupled.scala 375:21]
  wire [1:0] io_to_noc_1_flit_q_io_enq_bits_egress_id; // @[Decoupled.scala 375:21]
  wire  io_to_noc_1_flit_q_io_deq_ready; // @[Decoupled.scala 375:21]
  wire  io_to_noc_1_flit_q_io_deq_valid; // @[Decoupled.scala 375:21]
  wire  io_to_noc_1_flit_q_io_deq_bits_head; // @[Decoupled.scala 375:21]
  wire  io_to_noc_1_flit_q_io_deq_bits_tail; // @[Decoupled.scala 375:21]
  wire [63:0] io_to_noc_1_flit_q_io_deq_bits_payload; // @[Decoupled.scala 375:21]
  wire [1:0] io_to_noc_1_flit_q_io_deq_bits_egress_id; // @[Decoupled.scala 375:21]
  wire  igen_2_clock; // @[TestHarness.scala 171:22]
  wire  igen_2_reset; // @[TestHarness.scala 171:22]
  wire  igen_2_io_out_ready; // @[TestHarness.scala 171:22]
  wire  igen_2_io_out_valid; // @[TestHarness.scala 171:22]
  wire  igen_2_io_out_bits_head; // @[TestHarness.scala 171:22]
  wire  igen_2_io_out_bits_tail; // @[TestHarness.scala 171:22]
  wire [63:0] igen_2_io_out_bits_payload; // @[TestHarness.scala 171:22]
  wire [1:0] igen_2_io_out_bits_egress_id; // @[TestHarness.scala 171:22]
  wire  igen_2_io_rob_ready; // @[TestHarness.scala 171:22]
  wire [6:0] igen_2_io_rob_idx; // @[TestHarness.scala 171:22]
  wire [31:0] igen_2_io_tsc; // @[TestHarness.scala 171:22]
  wire  igen_2_io_fire; // @[TestHarness.scala 171:22]
  wire [3:0] igen_2_io_n_flits; // @[TestHarness.scala 171:22]
  wire  io_to_noc_2_flit_q_clock; // @[Decoupled.scala 375:21]
  wire  io_to_noc_2_flit_q_reset; // @[Decoupled.scala 375:21]
  wire  io_to_noc_2_flit_q_io_enq_ready; // @[Decoupled.scala 375:21]
  wire  io_to_noc_2_flit_q_io_enq_valid; // @[Decoupled.scala 375:21]
  wire  io_to_noc_2_flit_q_io_enq_bits_head; // @[Decoupled.scala 375:21]
  wire  io_to_noc_2_flit_q_io_enq_bits_tail; // @[Decoupled.scala 375:21]
  wire [63:0] io_to_noc_2_flit_q_io_enq_bits_payload; // @[Decoupled.scala 375:21]
  wire [1:0] io_to_noc_2_flit_q_io_enq_bits_egress_id; // @[Decoupled.scala 375:21]
  wire  io_to_noc_2_flit_q_io_deq_ready; // @[Decoupled.scala 375:21]
  wire  io_to_noc_2_flit_q_io_deq_valid; // @[Decoupled.scala 375:21]
  wire  io_to_noc_2_flit_q_io_deq_bits_head; // @[Decoupled.scala 375:21]
  wire  io_to_noc_2_flit_q_io_deq_bits_tail; // @[Decoupled.scala 375:21]
  wire [63:0] io_to_noc_2_flit_q_io_deq_bits_payload; // @[Decoupled.scala 375:21]
  wire [1:0] io_to_noc_2_flit_q_io_deq_bits_egress_id; // @[Decoupled.scala 375:21]
  wire  igen_3_clock; // @[TestHarness.scala 171:22]
  wire  igen_3_reset; // @[TestHarness.scala 171:22]
  wire  igen_3_io_out_ready; // @[TestHarness.scala 171:22]
  wire  igen_3_io_out_valid; // @[TestHarness.scala 171:22]
  wire  igen_3_io_out_bits_head; // @[TestHarness.scala 171:22]
  wire  igen_3_io_out_bits_tail; // @[TestHarness.scala 171:22]
  wire [63:0] igen_3_io_out_bits_payload; // @[TestHarness.scala 171:22]
  wire [1:0] igen_3_io_out_bits_egress_id; // @[TestHarness.scala 171:22]
  wire  igen_3_io_rob_ready; // @[TestHarness.scala 171:22]
  wire [6:0] igen_3_io_rob_idx; // @[TestHarness.scala 171:22]
  wire [31:0] igen_3_io_tsc; // @[TestHarness.scala 171:22]
  wire  igen_3_io_fire; // @[TestHarness.scala 171:22]
  wire [3:0] igen_3_io_n_flits; // @[TestHarness.scala 171:22]
  wire  io_to_noc_3_flit_q_clock; // @[Decoupled.scala 375:21]
  wire  io_to_noc_3_flit_q_reset; // @[Decoupled.scala 375:21]
  wire  io_to_noc_3_flit_q_io_enq_ready; // @[Decoupled.scala 375:21]
  wire  io_to_noc_3_flit_q_io_enq_valid; // @[Decoupled.scala 375:21]
  wire  io_to_noc_3_flit_q_io_enq_bits_head; // @[Decoupled.scala 375:21]
  wire  io_to_noc_3_flit_q_io_enq_bits_tail; // @[Decoupled.scala 375:21]
  wire [63:0] io_to_noc_3_flit_q_io_enq_bits_payload; // @[Decoupled.scala 375:21]
  wire [1:0] io_to_noc_3_flit_q_io_enq_bits_egress_id; // @[Decoupled.scala 375:21]
  wire  io_to_noc_3_flit_q_io_deq_ready; // @[Decoupled.scala 375:21]
  wire  io_to_noc_3_flit_q_io_deq_valid; // @[Decoupled.scala 375:21]
  wire  io_to_noc_3_flit_q_io_deq_bits_head; // @[Decoupled.scala 375:21]
  wire  io_to_noc_3_flit_q_io_deq_bits_tail; // @[Decoupled.scala 375:21]
  wire [63:0] io_to_noc_3_flit_q_io_deq_bits_payload; // @[Decoupled.scala 375:21]
  wire [1:0] io_to_noc_3_flit_q_io_deq_bits_egress_id; // @[Decoupled.scala 375:21]
  wire  plusarg_reader_out; // @[PlusArg.scala 80:11]
  wire  io_from_noc_0_flit_ready_prng_clock; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_reset; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_0; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_1; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_2; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_3; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_4; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_5; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_6; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_7; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_8; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_9; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_10; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_11; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_12; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_13; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_14; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_15; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_16; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_17; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_18; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_19; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_clock; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_reset; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_io_out_0; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_io_out_1; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_io_out_2; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_io_out_3; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_io_out_4; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_io_out_5; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_io_out_6; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_io_out_7; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_io_out_8; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_io_out_9; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_io_out_10; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_io_out_11; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_io_out_12; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_io_out_13; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_io_out_14; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_io_out_15; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_io_out_16; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_io_out_17; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_io_out_18; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_io_out_19; // @[PRNG.scala 91:22]
  wire  io_from_noc_2_flit_ready_prng_clock; // @[PRNG.scala 91:22]
  wire  io_from_noc_2_flit_ready_prng_reset; // @[PRNG.scala 91:22]
  wire  io_from_noc_2_flit_ready_prng_io_out_0; // @[PRNG.scala 91:22]
  wire  io_from_noc_2_flit_ready_prng_io_out_1; // @[PRNG.scala 91:22]
  wire  io_from_noc_2_flit_ready_prng_io_out_2; // @[PRNG.scala 91:22]
  wire  io_from_noc_2_flit_ready_prng_io_out_3; // @[PRNG.scala 91:22]
  wire  io_from_noc_2_flit_ready_prng_io_out_4; // @[PRNG.scala 91:22]
  wire  io_from_noc_2_flit_ready_prng_io_out_5; // @[PRNG.scala 91:22]
  wire  io_from_noc_2_flit_ready_prng_io_out_6; // @[PRNG.scala 91:22]
  wire  io_from_noc_2_flit_ready_prng_io_out_7; // @[PRNG.scala 91:22]
  wire  io_from_noc_2_flit_ready_prng_io_out_8; // @[PRNG.scala 91:22]
  wire  io_from_noc_2_flit_ready_prng_io_out_9; // @[PRNG.scala 91:22]
  wire  io_from_noc_2_flit_ready_prng_io_out_10; // @[PRNG.scala 91:22]
  wire  io_from_noc_2_flit_ready_prng_io_out_11; // @[PRNG.scala 91:22]
  wire  io_from_noc_2_flit_ready_prng_io_out_12; // @[PRNG.scala 91:22]
  wire  io_from_noc_2_flit_ready_prng_io_out_13; // @[PRNG.scala 91:22]
  wire  io_from_noc_2_flit_ready_prng_io_out_14; // @[PRNG.scala 91:22]
  wire  io_from_noc_2_flit_ready_prng_io_out_15; // @[PRNG.scala 91:22]
  wire  io_from_noc_2_flit_ready_prng_io_out_16; // @[PRNG.scala 91:22]
  wire  io_from_noc_2_flit_ready_prng_io_out_17; // @[PRNG.scala 91:22]
  wire  io_from_noc_2_flit_ready_prng_io_out_18; // @[PRNG.scala 91:22]
  wire  io_from_noc_2_flit_ready_prng_io_out_19; // @[PRNG.scala 91:22]
  wire  io_from_noc_3_flit_ready_prng_clock; // @[PRNG.scala 91:22]
  wire  io_from_noc_3_flit_ready_prng_reset; // @[PRNG.scala 91:22]
  wire  io_from_noc_3_flit_ready_prng_io_out_0; // @[PRNG.scala 91:22]
  wire  io_from_noc_3_flit_ready_prng_io_out_1; // @[PRNG.scala 91:22]
  wire  io_from_noc_3_flit_ready_prng_io_out_2; // @[PRNG.scala 91:22]
  wire  io_from_noc_3_flit_ready_prng_io_out_3; // @[PRNG.scala 91:22]
  wire  io_from_noc_3_flit_ready_prng_io_out_4; // @[PRNG.scala 91:22]
  wire  io_from_noc_3_flit_ready_prng_io_out_5; // @[PRNG.scala 91:22]
  wire  io_from_noc_3_flit_ready_prng_io_out_6; // @[PRNG.scala 91:22]
  wire  io_from_noc_3_flit_ready_prng_io_out_7; // @[PRNG.scala 91:22]
  wire  io_from_noc_3_flit_ready_prng_io_out_8; // @[PRNG.scala 91:22]
  wire  io_from_noc_3_flit_ready_prng_io_out_9; // @[PRNG.scala 91:22]
  wire  io_from_noc_3_flit_ready_prng_io_out_10; // @[PRNG.scala 91:22]
  wire  io_from_noc_3_flit_ready_prng_io_out_11; // @[PRNG.scala 91:22]
  wire  io_from_noc_3_flit_ready_prng_io_out_12; // @[PRNG.scala 91:22]
  wire  io_from_noc_3_flit_ready_prng_io_out_13; // @[PRNG.scala 91:22]
  wire  io_from_noc_3_flit_ready_prng_io_out_14; // @[PRNG.scala 91:22]
  wire  io_from_noc_3_flit_ready_prng_io_out_15; // @[PRNG.scala 91:22]
  wire  io_from_noc_3_flit_ready_prng_io_out_16; // @[PRNG.scala 91:22]
  wire  io_from_noc_3_flit_ready_prng_io_out_17; // @[PRNG.scala 91:22]
  wire  io_from_noc_3_flit_ready_prng_io_out_18; // @[PRNG.scala 91:22]
  wire  io_from_noc_3_flit_ready_prng_io_out_19; // @[PRNG.scala 91:22]
  reg [31:0] txs; // @[TestHarness.scala 136:20]
  reg [31:0] flits; // @[TestHarness.scala 137:22]
  reg [31:0] tsc; // @[TestHarness.scala 141:20]
  wire [31:0] _tsc_T_1 = tsc + 32'h1; // @[TestHarness.scala 142:14]
  reg [10:0] idle_counter; // @[TestHarness.scala 144:29]
  wire [10:0] _idle_counter_T_1 = idle_counter + 11'h1; // @[TestHarness.scala 146:46]
  reg [127:0] rob_valids; // @[TestHarness.scala 156:27]
  wire [127:0] _T_5 = ~rob_valids; // @[TestHarness.scala 161:59]
  wire [6:0] _sels_0_T_128 = _T_5[126] ? 7'h7e : 7'h7f; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_129 = _T_5[125] ? 7'h7d : _sels_0_T_128; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_130 = _T_5[124] ? 7'h7c : _sels_0_T_129; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_131 = _T_5[123] ? 7'h7b : _sels_0_T_130; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_132 = _T_5[122] ? 7'h7a : _sels_0_T_131; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_133 = _T_5[121] ? 7'h79 : _sels_0_T_132; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_134 = _T_5[120] ? 7'h78 : _sels_0_T_133; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_135 = _T_5[119] ? 7'h77 : _sels_0_T_134; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_136 = _T_5[118] ? 7'h76 : _sels_0_T_135; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_137 = _T_5[117] ? 7'h75 : _sels_0_T_136; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_138 = _T_5[116] ? 7'h74 : _sels_0_T_137; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_139 = _T_5[115] ? 7'h73 : _sels_0_T_138; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_140 = _T_5[114] ? 7'h72 : _sels_0_T_139; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_141 = _T_5[113] ? 7'h71 : _sels_0_T_140; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_142 = _T_5[112] ? 7'h70 : _sels_0_T_141; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_143 = _T_5[111] ? 7'h6f : _sels_0_T_142; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_144 = _T_5[110] ? 7'h6e : _sels_0_T_143; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_145 = _T_5[109] ? 7'h6d : _sels_0_T_144; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_146 = _T_5[108] ? 7'h6c : _sels_0_T_145; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_147 = _T_5[107] ? 7'h6b : _sels_0_T_146; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_148 = _T_5[106] ? 7'h6a : _sels_0_T_147; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_149 = _T_5[105] ? 7'h69 : _sels_0_T_148; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_150 = _T_5[104] ? 7'h68 : _sels_0_T_149; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_151 = _T_5[103] ? 7'h67 : _sels_0_T_150; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_152 = _T_5[102] ? 7'h66 : _sels_0_T_151; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_153 = _T_5[101] ? 7'h65 : _sels_0_T_152; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_154 = _T_5[100] ? 7'h64 : _sels_0_T_153; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_155 = _T_5[99] ? 7'h63 : _sels_0_T_154; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_156 = _T_5[98] ? 7'h62 : _sels_0_T_155; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_157 = _T_5[97] ? 7'h61 : _sels_0_T_156; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_158 = _T_5[96] ? 7'h60 : _sels_0_T_157; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_159 = _T_5[95] ? 7'h5f : _sels_0_T_158; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_160 = _T_5[94] ? 7'h5e : _sels_0_T_159; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_161 = _T_5[93] ? 7'h5d : _sels_0_T_160; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_162 = _T_5[92] ? 7'h5c : _sels_0_T_161; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_163 = _T_5[91] ? 7'h5b : _sels_0_T_162; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_164 = _T_5[90] ? 7'h5a : _sels_0_T_163; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_165 = _T_5[89] ? 7'h59 : _sels_0_T_164; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_166 = _T_5[88] ? 7'h58 : _sels_0_T_165; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_167 = _T_5[87] ? 7'h57 : _sels_0_T_166; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_168 = _T_5[86] ? 7'h56 : _sels_0_T_167; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_169 = _T_5[85] ? 7'h55 : _sels_0_T_168; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_170 = _T_5[84] ? 7'h54 : _sels_0_T_169; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_171 = _T_5[83] ? 7'h53 : _sels_0_T_170; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_172 = _T_5[82] ? 7'h52 : _sels_0_T_171; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_173 = _T_5[81] ? 7'h51 : _sels_0_T_172; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_174 = _T_5[80] ? 7'h50 : _sels_0_T_173; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_175 = _T_5[79] ? 7'h4f : _sels_0_T_174; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_176 = _T_5[78] ? 7'h4e : _sels_0_T_175; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_177 = _T_5[77] ? 7'h4d : _sels_0_T_176; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_178 = _T_5[76] ? 7'h4c : _sels_0_T_177; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_179 = _T_5[75] ? 7'h4b : _sels_0_T_178; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_180 = _T_5[74] ? 7'h4a : _sels_0_T_179; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_181 = _T_5[73] ? 7'h49 : _sels_0_T_180; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_182 = _T_5[72] ? 7'h48 : _sels_0_T_181; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_183 = _T_5[71] ? 7'h47 : _sels_0_T_182; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_184 = _T_5[70] ? 7'h46 : _sels_0_T_183; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_185 = _T_5[69] ? 7'h45 : _sels_0_T_184; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_186 = _T_5[68] ? 7'h44 : _sels_0_T_185; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_187 = _T_5[67] ? 7'h43 : _sels_0_T_186; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_188 = _T_5[66] ? 7'h42 : _sels_0_T_187; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_189 = _T_5[65] ? 7'h41 : _sels_0_T_188; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_190 = _T_5[64] ? 7'h40 : _sels_0_T_189; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_191 = _T_5[63] ? 7'h3f : _sels_0_T_190; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_192 = _T_5[62] ? 7'h3e : _sels_0_T_191; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_193 = _T_5[61] ? 7'h3d : _sels_0_T_192; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_194 = _T_5[60] ? 7'h3c : _sels_0_T_193; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_195 = _T_5[59] ? 7'h3b : _sels_0_T_194; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_196 = _T_5[58] ? 7'h3a : _sels_0_T_195; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_197 = _T_5[57] ? 7'h39 : _sels_0_T_196; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_198 = _T_5[56] ? 7'h38 : _sels_0_T_197; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_199 = _T_5[55] ? 7'h37 : _sels_0_T_198; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_200 = _T_5[54] ? 7'h36 : _sels_0_T_199; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_201 = _T_5[53] ? 7'h35 : _sels_0_T_200; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_202 = _T_5[52] ? 7'h34 : _sels_0_T_201; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_203 = _T_5[51] ? 7'h33 : _sels_0_T_202; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_204 = _T_5[50] ? 7'h32 : _sels_0_T_203; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_205 = _T_5[49] ? 7'h31 : _sels_0_T_204; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_206 = _T_5[48] ? 7'h30 : _sels_0_T_205; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_207 = _T_5[47] ? 7'h2f : _sels_0_T_206; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_208 = _T_5[46] ? 7'h2e : _sels_0_T_207; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_209 = _T_5[45] ? 7'h2d : _sels_0_T_208; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_210 = _T_5[44] ? 7'h2c : _sels_0_T_209; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_211 = _T_5[43] ? 7'h2b : _sels_0_T_210; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_212 = _T_5[42] ? 7'h2a : _sels_0_T_211; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_213 = _T_5[41] ? 7'h29 : _sels_0_T_212; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_214 = _T_5[40] ? 7'h28 : _sels_0_T_213; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_215 = _T_5[39] ? 7'h27 : _sels_0_T_214; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_216 = _T_5[38] ? 7'h26 : _sels_0_T_215; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_217 = _T_5[37] ? 7'h25 : _sels_0_T_216; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_218 = _T_5[36] ? 7'h24 : _sels_0_T_217; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_219 = _T_5[35] ? 7'h23 : _sels_0_T_218; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_220 = _T_5[34] ? 7'h22 : _sels_0_T_219; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_221 = _T_5[33] ? 7'h21 : _sels_0_T_220; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_222 = _T_5[32] ? 7'h20 : _sels_0_T_221; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_223 = _T_5[31] ? 7'h1f : _sels_0_T_222; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_224 = _T_5[30] ? 7'h1e : _sels_0_T_223; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_225 = _T_5[29] ? 7'h1d : _sels_0_T_224; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_226 = _T_5[28] ? 7'h1c : _sels_0_T_225; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_227 = _T_5[27] ? 7'h1b : _sels_0_T_226; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_228 = _T_5[26] ? 7'h1a : _sels_0_T_227; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_229 = _T_5[25] ? 7'h19 : _sels_0_T_228; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_230 = _T_5[24] ? 7'h18 : _sels_0_T_229; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_231 = _T_5[23] ? 7'h17 : _sels_0_T_230; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_232 = _T_5[22] ? 7'h16 : _sels_0_T_231; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_233 = _T_5[21] ? 7'h15 : _sels_0_T_232; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_234 = _T_5[20] ? 7'h14 : _sels_0_T_233; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_235 = _T_5[19] ? 7'h13 : _sels_0_T_234; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_236 = _T_5[18] ? 7'h12 : _sels_0_T_235; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_237 = _T_5[17] ? 7'h11 : _sels_0_T_236; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_238 = _T_5[16] ? 7'h10 : _sels_0_T_237; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_239 = _T_5[15] ? 7'hf : _sels_0_T_238; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_240 = _T_5[14] ? 7'he : _sels_0_T_239; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_241 = _T_5[13] ? 7'hd : _sels_0_T_240; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_242 = _T_5[12] ? 7'hc : _sels_0_T_241; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_243 = _T_5[11] ? 7'hb : _sels_0_T_242; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_244 = _T_5[10] ? 7'ha : _sels_0_T_243; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_245 = _T_5[9] ? 7'h9 : _sels_0_T_244; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_246 = _T_5[8] ? 7'h8 : _sels_0_T_245; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_247 = _T_5[7] ? 7'h7 : _sels_0_T_246; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_248 = _T_5[6] ? 7'h6 : _sels_0_T_247; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_249 = _T_5[5] ? 7'h5 : _sels_0_T_248; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_250 = _T_5[4] ? 7'h4 : _sels_0_T_249; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_251 = _T_5[3] ? 7'h3 : _sels_0_T_250; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_252 = _T_5[2] ? 7'h2 : _sels_0_T_251; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_253 = _T_5[1] ? 7'h1 : _sels_0_T_252; // @[Mux.scala 47:70]
  wire [6:0] rob_alloc_ids_0 = _T_5[0] ? 7'h0 : _sels_0_T_253; // @[Mux.scala 47:70]
  wire [127:0] _GEN_7169 = {{127'd0}, igen_io_fire}; // @[TestHarness.scala 187:45]
  wire [127:0] _T_32 = _GEN_7169 << rob_alloc_ids_0; // @[TestHarness.scala 187:45]
  wire [127:0] _T_6 = 128'h1 << rob_alloc_ids_0; // @[TestHarness.scala 31:27]
  wire [127:0] _T_7 = ~_T_6; // @[TestHarness.scala 31:21]
  wire [127:0] _T_8 = _T_5 & _T_7; // @[TestHarness.scala 31:19]
  wire [6:0] _sels_1_T_128 = _T_8[126] ? 7'h7e : 7'h7f; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_129 = _T_8[125] ? 7'h7d : _sels_1_T_128; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_130 = _T_8[124] ? 7'h7c : _sels_1_T_129; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_131 = _T_8[123] ? 7'h7b : _sels_1_T_130; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_132 = _T_8[122] ? 7'h7a : _sels_1_T_131; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_133 = _T_8[121] ? 7'h79 : _sels_1_T_132; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_134 = _T_8[120] ? 7'h78 : _sels_1_T_133; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_135 = _T_8[119] ? 7'h77 : _sels_1_T_134; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_136 = _T_8[118] ? 7'h76 : _sels_1_T_135; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_137 = _T_8[117] ? 7'h75 : _sels_1_T_136; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_138 = _T_8[116] ? 7'h74 : _sels_1_T_137; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_139 = _T_8[115] ? 7'h73 : _sels_1_T_138; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_140 = _T_8[114] ? 7'h72 : _sels_1_T_139; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_141 = _T_8[113] ? 7'h71 : _sels_1_T_140; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_142 = _T_8[112] ? 7'h70 : _sels_1_T_141; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_143 = _T_8[111] ? 7'h6f : _sels_1_T_142; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_144 = _T_8[110] ? 7'h6e : _sels_1_T_143; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_145 = _T_8[109] ? 7'h6d : _sels_1_T_144; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_146 = _T_8[108] ? 7'h6c : _sels_1_T_145; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_147 = _T_8[107] ? 7'h6b : _sels_1_T_146; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_148 = _T_8[106] ? 7'h6a : _sels_1_T_147; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_149 = _T_8[105] ? 7'h69 : _sels_1_T_148; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_150 = _T_8[104] ? 7'h68 : _sels_1_T_149; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_151 = _T_8[103] ? 7'h67 : _sels_1_T_150; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_152 = _T_8[102] ? 7'h66 : _sels_1_T_151; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_153 = _T_8[101] ? 7'h65 : _sels_1_T_152; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_154 = _T_8[100] ? 7'h64 : _sels_1_T_153; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_155 = _T_8[99] ? 7'h63 : _sels_1_T_154; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_156 = _T_8[98] ? 7'h62 : _sels_1_T_155; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_157 = _T_8[97] ? 7'h61 : _sels_1_T_156; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_158 = _T_8[96] ? 7'h60 : _sels_1_T_157; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_159 = _T_8[95] ? 7'h5f : _sels_1_T_158; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_160 = _T_8[94] ? 7'h5e : _sels_1_T_159; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_161 = _T_8[93] ? 7'h5d : _sels_1_T_160; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_162 = _T_8[92] ? 7'h5c : _sels_1_T_161; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_163 = _T_8[91] ? 7'h5b : _sels_1_T_162; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_164 = _T_8[90] ? 7'h5a : _sels_1_T_163; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_165 = _T_8[89] ? 7'h59 : _sels_1_T_164; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_166 = _T_8[88] ? 7'h58 : _sels_1_T_165; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_167 = _T_8[87] ? 7'h57 : _sels_1_T_166; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_168 = _T_8[86] ? 7'h56 : _sels_1_T_167; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_169 = _T_8[85] ? 7'h55 : _sels_1_T_168; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_170 = _T_8[84] ? 7'h54 : _sels_1_T_169; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_171 = _T_8[83] ? 7'h53 : _sels_1_T_170; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_172 = _T_8[82] ? 7'h52 : _sels_1_T_171; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_173 = _T_8[81] ? 7'h51 : _sels_1_T_172; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_174 = _T_8[80] ? 7'h50 : _sels_1_T_173; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_175 = _T_8[79] ? 7'h4f : _sels_1_T_174; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_176 = _T_8[78] ? 7'h4e : _sels_1_T_175; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_177 = _T_8[77] ? 7'h4d : _sels_1_T_176; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_178 = _T_8[76] ? 7'h4c : _sels_1_T_177; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_179 = _T_8[75] ? 7'h4b : _sels_1_T_178; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_180 = _T_8[74] ? 7'h4a : _sels_1_T_179; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_181 = _T_8[73] ? 7'h49 : _sels_1_T_180; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_182 = _T_8[72] ? 7'h48 : _sels_1_T_181; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_183 = _T_8[71] ? 7'h47 : _sels_1_T_182; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_184 = _T_8[70] ? 7'h46 : _sels_1_T_183; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_185 = _T_8[69] ? 7'h45 : _sels_1_T_184; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_186 = _T_8[68] ? 7'h44 : _sels_1_T_185; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_187 = _T_8[67] ? 7'h43 : _sels_1_T_186; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_188 = _T_8[66] ? 7'h42 : _sels_1_T_187; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_189 = _T_8[65] ? 7'h41 : _sels_1_T_188; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_190 = _T_8[64] ? 7'h40 : _sels_1_T_189; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_191 = _T_8[63] ? 7'h3f : _sels_1_T_190; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_192 = _T_8[62] ? 7'h3e : _sels_1_T_191; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_193 = _T_8[61] ? 7'h3d : _sels_1_T_192; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_194 = _T_8[60] ? 7'h3c : _sels_1_T_193; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_195 = _T_8[59] ? 7'h3b : _sels_1_T_194; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_196 = _T_8[58] ? 7'h3a : _sels_1_T_195; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_197 = _T_8[57] ? 7'h39 : _sels_1_T_196; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_198 = _T_8[56] ? 7'h38 : _sels_1_T_197; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_199 = _T_8[55] ? 7'h37 : _sels_1_T_198; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_200 = _T_8[54] ? 7'h36 : _sels_1_T_199; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_201 = _T_8[53] ? 7'h35 : _sels_1_T_200; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_202 = _T_8[52] ? 7'h34 : _sels_1_T_201; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_203 = _T_8[51] ? 7'h33 : _sels_1_T_202; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_204 = _T_8[50] ? 7'h32 : _sels_1_T_203; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_205 = _T_8[49] ? 7'h31 : _sels_1_T_204; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_206 = _T_8[48] ? 7'h30 : _sels_1_T_205; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_207 = _T_8[47] ? 7'h2f : _sels_1_T_206; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_208 = _T_8[46] ? 7'h2e : _sels_1_T_207; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_209 = _T_8[45] ? 7'h2d : _sels_1_T_208; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_210 = _T_8[44] ? 7'h2c : _sels_1_T_209; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_211 = _T_8[43] ? 7'h2b : _sels_1_T_210; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_212 = _T_8[42] ? 7'h2a : _sels_1_T_211; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_213 = _T_8[41] ? 7'h29 : _sels_1_T_212; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_214 = _T_8[40] ? 7'h28 : _sels_1_T_213; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_215 = _T_8[39] ? 7'h27 : _sels_1_T_214; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_216 = _T_8[38] ? 7'h26 : _sels_1_T_215; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_217 = _T_8[37] ? 7'h25 : _sels_1_T_216; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_218 = _T_8[36] ? 7'h24 : _sels_1_T_217; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_219 = _T_8[35] ? 7'h23 : _sels_1_T_218; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_220 = _T_8[34] ? 7'h22 : _sels_1_T_219; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_221 = _T_8[33] ? 7'h21 : _sels_1_T_220; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_222 = _T_8[32] ? 7'h20 : _sels_1_T_221; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_223 = _T_8[31] ? 7'h1f : _sels_1_T_222; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_224 = _T_8[30] ? 7'h1e : _sels_1_T_223; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_225 = _T_8[29] ? 7'h1d : _sels_1_T_224; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_226 = _T_8[28] ? 7'h1c : _sels_1_T_225; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_227 = _T_8[27] ? 7'h1b : _sels_1_T_226; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_228 = _T_8[26] ? 7'h1a : _sels_1_T_227; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_229 = _T_8[25] ? 7'h19 : _sels_1_T_228; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_230 = _T_8[24] ? 7'h18 : _sels_1_T_229; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_231 = _T_8[23] ? 7'h17 : _sels_1_T_230; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_232 = _T_8[22] ? 7'h16 : _sels_1_T_231; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_233 = _T_8[21] ? 7'h15 : _sels_1_T_232; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_234 = _T_8[20] ? 7'h14 : _sels_1_T_233; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_235 = _T_8[19] ? 7'h13 : _sels_1_T_234; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_236 = _T_8[18] ? 7'h12 : _sels_1_T_235; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_237 = _T_8[17] ? 7'h11 : _sels_1_T_236; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_238 = _T_8[16] ? 7'h10 : _sels_1_T_237; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_239 = _T_8[15] ? 7'hf : _sels_1_T_238; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_240 = _T_8[14] ? 7'he : _sels_1_T_239; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_241 = _T_8[13] ? 7'hd : _sels_1_T_240; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_242 = _T_8[12] ? 7'hc : _sels_1_T_241; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_243 = _T_8[11] ? 7'hb : _sels_1_T_242; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_244 = _T_8[10] ? 7'ha : _sels_1_T_243; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_245 = _T_8[9] ? 7'h9 : _sels_1_T_244; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_246 = _T_8[8] ? 7'h8 : _sels_1_T_245; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_247 = _T_8[7] ? 7'h7 : _sels_1_T_246; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_248 = _T_8[6] ? 7'h6 : _sels_1_T_247; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_249 = _T_8[5] ? 7'h5 : _sels_1_T_248; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_250 = _T_8[4] ? 7'h4 : _sels_1_T_249; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_251 = _T_8[3] ? 7'h3 : _sels_1_T_250; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_252 = _T_8[2] ? 7'h2 : _sels_1_T_251; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_253 = _T_8[1] ? 7'h1 : _sels_1_T_252; // @[Mux.scala 47:70]
  wire [6:0] rob_alloc_ids_1 = _T_8[0] ? 7'h0 : _sels_1_T_253; // @[Mux.scala 47:70]
  wire [127:0] _GEN_7170 = {{127'd0}, igen_1_io_fire}; // @[TestHarness.scala 187:45]
  wire [127:0] _T_46 = _GEN_7170 << rob_alloc_ids_1; // @[TestHarness.scala 187:45]
  wire [127:0] _T_47 = _T_32 | _T_46; // @[TestHarness.scala 187:29]
  wire [127:0] _T_9 = 128'h1 << rob_alloc_ids_1; // @[TestHarness.scala 31:27]
  wire [127:0] _T_10 = ~_T_9; // @[TestHarness.scala 31:21]
  wire [127:0] _T_11 = _T_8 & _T_10; // @[TestHarness.scala 31:19]
  wire [6:0] _sels_2_T_128 = _T_11[126] ? 7'h7e : 7'h7f; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_129 = _T_11[125] ? 7'h7d : _sels_2_T_128; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_130 = _T_11[124] ? 7'h7c : _sels_2_T_129; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_131 = _T_11[123] ? 7'h7b : _sels_2_T_130; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_132 = _T_11[122] ? 7'h7a : _sels_2_T_131; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_133 = _T_11[121] ? 7'h79 : _sels_2_T_132; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_134 = _T_11[120] ? 7'h78 : _sels_2_T_133; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_135 = _T_11[119] ? 7'h77 : _sels_2_T_134; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_136 = _T_11[118] ? 7'h76 : _sels_2_T_135; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_137 = _T_11[117] ? 7'h75 : _sels_2_T_136; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_138 = _T_11[116] ? 7'h74 : _sels_2_T_137; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_139 = _T_11[115] ? 7'h73 : _sels_2_T_138; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_140 = _T_11[114] ? 7'h72 : _sels_2_T_139; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_141 = _T_11[113] ? 7'h71 : _sels_2_T_140; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_142 = _T_11[112] ? 7'h70 : _sels_2_T_141; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_143 = _T_11[111] ? 7'h6f : _sels_2_T_142; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_144 = _T_11[110] ? 7'h6e : _sels_2_T_143; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_145 = _T_11[109] ? 7'h6d : _sels_2_T_144; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_146 = _T_11[108] ? 7'h6c : _sels_2_T_145; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_147 = _T_11[107] ? 7'h6b : _sels_2_T_146; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_148 = _T_11[106] ? 7'h6a : _sels_2_T_147; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_149 = _T_11[105] ? 7'h69 : _sels_2_T_148; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_150 = _T_11[104] ? 7'h68 : _sels_2_T_149; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_151 = _T_11[103] ? 7'h67 : _sels_2_T_150; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_152 = _T_11[102] ? 7'h66 : _sels_2_T_151; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_153 = _T_11[101] ? 7'h65 : _sels_2_T_152; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_154 = _T_11[100] ? 7'h64 : _sels_2_T_153; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_155 = _T_11[99] ? 7'h63 : _sels_2_T_154; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_156 = _T_11[98] ? 7'h62 : _sels_2_T_155; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_157 = _T_11[97] ? 7'h61 : _sels_2_T_156; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_158 = _T_11[96] ? 7'h60 : _sels_2_T_157; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_159 = _T_11[95] ? 7'h5f : _sels_2_T_158; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_160 = _T_11[94] ? 7'h5e : _sels_2_T_159; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_161 = _T_11[93] ? 7'h5d : _sels_2_T_160; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_162 = _T_11[92] ? 7'h5c : _sels_2_T_161; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_163 = _T_11[91] ? 7'h5b : _sels_2_T_162; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_164 = _T_11[90] ? 7'h5a : _sels_2_T_163; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_165 = _T_11[89] ? 7'h59 : _sels_2_T_164; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_166 = _T_11[88] ? 7'h58 : _sels_2_T_165; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_167 = _T_11[87] ? 7'h57 : _sels_2_T_166; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_168 = _T_11[86] ? 7'h56 : _sels_2_T_167; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_169 = _T_11[85] ? 7'h55 : _sels_2_T_168; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_170 = _T_11[84] ? 7'h54 : _sels_2_T_169; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_171 = _T_11[83] ? 7'h53 : _sels_2_T_170; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_172 = _T_11[82] ? 7'h52 : _sels_2_T_171; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_173 = _T_11[81] ? 7'h51 : _sels_2_T_172; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_174 = _T_11[80] ? 7'h50 : _sels_2_T_173; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_175 = _T_11[79] ? 7'h4f : _sels_2_T_174; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_176 = _T_11[78] ? 7'h4e : _sels_2_T_175; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_177 = _T_11[77] ? 7'h4d : _sels_2_T_176; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_178 = _T_11[76] ? 7'h4c : _sels_2_T_177; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_179 = _T_11[75] ? 7'h4b : _sels_2_T_178; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_180 = _T_11[74] ? 7'h4a : _sels_2_T_179; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_181 = _T_11[73] ? 7'h49 : _sels_2_T_180; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_182 = _T_11[72] ? 7'h48 : _sels_2_T_181; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_183 = _T_11[71] ? 7'h47 : _sels_2_T_182; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_184 = _T_11[70] ? 7'h46 : _sels_2_T_183; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_185 = _T_11[69] ? 7'h45 : _sels_2_T_184; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_186 = _T_11[68] ? 7'h44 : _sels_2_T_185; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_187 = _T_11[67] ? 7'h43 : _sels_2_T_186; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_188 = _T_11[66] ? 7'h42 : _sels_2_T_187; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_189 = _T_11[65] ? 7'h41 : _sels_2_T_188; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_190 = _T_11[64] ? 7'h40 : _sels_2_T_189; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_191 = _T_11[63] ? 7'h3f : _sels_2_T_190; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_192 = _T_11[62] ? 7'h3e : _sels_2_T_191; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_193 = _T_11[61] ? 7'h3d : _sels_2_T_192; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_194 = _T_11[60] ? 7'h3c : _sels_2_T_193; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_195 = _T_11[59] ? 7'h3b : _sels_2_T_194; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_196 = _T_11[58] ? 7'h3a : _sels_2_T_195; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_197 = _T_11[57] ? 7'h39 : _sels_2_T_196; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_198 = _T_11[56] ? 7'h38 : _sels_2_T_197; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_199 = _T_11[55] ? 7'h37 : _sels_2_T_198; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_200 = _T_11[54] ? 7'h36 : _sels_2_T_199; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_201 = _T_11[53] ? 7'h35 : _sels_2_T_200; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_202 = _T_11[52] ? 7'h34 : _sels_2_T_201; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_203 = _T_11[51] ? 7'h33 : _sels_2_T_202; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_204 = _T_11[50] ? 7'h32 : _sels_2_T_203; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_205 = _T_11[49] ? 7'h31 : _sels_2_T_204; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_206 = _T_11[48] ? 7'h30 : _sels_2_T_205; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_207 = _T_11[47] ? 7'h2f : _sels_2_T_206; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_208 = _T_11[46] ? 7'h2e : _sels_2_T_207; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_209 = _T_11[45] ? 7'h2d : _sels_2_T_208; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_210 = _T_11[44] ? 7'h2c : _sels_2_T_209; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_211 = _T_11[43] ? 7'h2b : _sels_2_T_210; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_212 = _T_11[42] ? 7'h2a : _sels_2_T_211; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_213 = _T_11[41] ? 7'h29 : _sels_2_T_212; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_214 = _T_11[40] ? 7'h28 : _sels_2_T_213; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_215 = _T_11[39] ? 7'h27 : _sels_2_T_214; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_216 = _T_11[38] ? 7'h26 : _sels_2_T_215; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_217 = _T_11[37] ? 7'h25 : _sels_2_T_216; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_218 = _T_11[36] ? 7'h24 : _sels_2_T_217; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_219 = _T_11[35] ? 7'h23 : _sels_2_T_218; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_220 = _T_11[34] ? 7'h22 : _sels_2_T_219; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_221 = _T_11[33] ? 7'h21 : _sels_2_T_220; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_222 = _T_11[32] ? 7'h20 : _sels_2_T_221; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_223 = _T_11[31] ? 7'h1f : _sels_2_T_222; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_224 = _T_11[30] ? 7'h1e : _sels_2_T_223; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_225 = _T_11[29] ? 7'h1d : _sels_2_T_224; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_226 = _T_11[28] ? 7'h1c : _sels_2_T_225; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_227 = _T_11[27] ? 7'h1b : _sels_2_T_226; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_228 = _T_11[26] ? 7'h1a : _sels_2_T_227; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_229 = _T_11[25] ? 7'h19 : _sels_2_T_228; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_230 = _T_11[24] ? 7'h18 : _sels_2_T_229; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_231 = _T_11[23] ? 7'h17 : _sels_2_T_230; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_232 = _T_11[22] ? 7'h16 : _sels_2_T_231; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_233 = _T_11[21] ? 7'h15 : _sels_2_T_232; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_234 = _T_11[20] ? 7'h14 : _sels_2_T_233; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_235 = _T_11[19] ? 7'h13 : _sels_2_T_234; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_236 = _T_11[18] ? 7'h12 : _sels_2_T_235; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_237 = _T_11[17] ? 7'h11 : _sels_2_T_236; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_238 = _T_11[16] ? 7'h10 : _sels_2_T_237; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_239 = _T_11[15] ? 7'hf : _sels_2_T_238; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_240 = _T_11[14] ? 7'he : _sels_2_T_239; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_241 = _T_11[13] ? 7'hd : _sels_2_T_240; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_242 = _T_11[12] ? 7'hc : _sels_2_T_241; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_243 = _T_11[11] ? 7'hb : _sels_2_T_242; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_244 = _T_11[10] ? 7'ha : _sels_2_T_243; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_245 = _T_11[9] ? 7'h9 : _sels_2_T_244; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_246 = _T_11[8] ? 7'h8 : _sels_2_T_245; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_247 = _T_11[7] ? 7'h7 : _sels_2_T_246; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_248 = _T_11[6] ? 7'h6 : _sels_2_T_247; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_249 = _T_11[5] ? 7'h5 : _sels_2_T_248; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_250 = _T_11[4] ? 7'h4 : _sels_2_T_249; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_251 = _T_11[3] ? 7'h3 : _sels_2_T_250; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_252 = _T_11[2] ? 7'h2 : _sels_2_T_251; // @[Mux.scala 47:70]
  wire [6:0] _sels_2_T_253 = _T_11[1] ? 7'h1 : _sels_2_T_252; // @[Mux.scala 47:70]
  wire [6:0] rob_alloc_ids_2 = _T_11[0] ? 7'h0 : _sels_2_T_253; // @[Mux.scala 47:70]
  wire [127:0] _GEN_7171 = {{127'd0}, igen_2_io_fire}; // @[TestHarness.scala 187:45]
  wire [127:0] _T_60 = _GEN_7171 << rob_alloc_ids_2; // @[TestHarness.scala 187:45]
  wire [127:0] _T_61 = _T_47 | _T_60; // @[TestHarness.scala 187:29]
  wire [127:0] _T_12 = 128'h1 << rob_alloc_ids_2; // @[TestHarness.scala 31:27]
  wire [127:0] _T_13 = ~_T_12; // @[TestHarness.scala 31:21]
  wire [127:0] _T_14 = _T_11 & _T_13; // @[TestHarness.scala 31:19]
  wire [6:0] _sels_3_T_128 = _T_14[126] ? 7'h7e : 7'h7f; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_129 = _T_14[125] ? 7'h7d : _sels_3_T_128; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_130 = _T_14[124] ? 7'h7c : _sels_3_T_129; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_131 = _T_14[123] ? 7'h7b : _sels_3_T_130; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_132 = _T_14[122] ? 7'h7a : _sels_3_T_131; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_133 = _T_14[121] ? 7'h79 : _sels_3_T_132; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_134 = _T_14[120] ? 7'h78 : _sels_3_T_133; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_135 = _T_14[119] ? 7'h77 : _sels_3_T_134; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_136 = _T_14[118] ? 7'h76 : _sels_3_T_135; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_137 = _T_14[117] ? 7'h75 : _sels_3_T_136; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_138 = _T_14[116] ? 7'h74 : _sels_3_T_137; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_139 = _T_14[115] ? 7'h73 : _sels_3_T_138; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_140 = _T_14[114] ? 7'h72 : _sels_3_T_139; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_141 = _T_14[113] ? 7'h71 : _sels_3_T_140; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_142 = _T_14[112] ? 7'h70 : _sels_3_T_141; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_143 = _T_14[111] ? 7'h6f : _sels_3_T_142; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_144 = _T_14[110] ? 7'h6e : _sels_3_T_143; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_145 = _T_14[109] ? 7'h6d : _sels_3_T_144; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_146 = _T_14[108] ? 7'h6c : _sels_3_T_145; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_147 = _T_14[107] ? 7'h6b : _sels_3_T_146; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_148 = _T_14[106] ? 7'h6a : _sels_3_T_147; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_149 = _T_14[105] ? 7'h69 : _sels_3_T_148; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_150 = _T_14[104] ? 7'h68 : _sels_3_T_149; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_151 = _T_14[103] ? 7'h67 : _sels_3_T_150; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_152 = _T_14[102] ? 7'h66 : _sels_3_T_151; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_153 = _T_14[101] ? 7'h65 : _sels_3_T_152; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_154 = _T_14[100] ? 7'h64 : _sels_3_T_153; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_155 = _T_14[99] ? 7'h63 : _sels_3_T_154; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_156 = _T_14[98] ? 7'h62 : _sels_3_T_155; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_157 = _T_14[97] ? 7'h61 : _sels_3_T_156; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_158 = _T_14[96] ? 7'h60 : _sels_3_T_157; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_159 = _T_14[95] ? 7'h5f : _sels_3_T_158; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_160 = _T_14[94] ? 7'h5e : _sels_3_T_159; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_161 = _T_14[93] ? 7'h5d : _sels_3_T_160; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_162 = _T_14[92] ? 7'h5c : _sels_3_T_161; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_163 = _T_14[91] ? 7'h5b : _sels_3_T_162; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_164 = _T_14[90] ? 7'h5a : _sels_3_T_163; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_165 = _T_14[89] ? 7'h59 : _sels_3_T_164; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_166 = _T_14[88] ? 7'h58 : _sels_3_T_165; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_167 = _T_14[87] ? 7'h57 : _sels_3_T_166; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_168 = _T_14[86] ? 7'h56 : _sels_3_T_167; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_169 = _T_14[85] ? 7'h55 : _sels_3_T_168; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_170 = _T_14[84] ? 7'h54 : _sels_3_T_169; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_171 = _T_14[83] ? 7'h53 : _sels_3_T_170; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_172 = _T_14[82] ? 7'h52 : _sels_3_T_171; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_173 = _T_14[81] ? 7'h51 : _sels_3_T_172; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_174 = _T_14[80] ? 7'h50 : _sels_3_T_173; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_175 = _T_14[79] ? 7'h4f : _sels_3_T_174; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_176 = _T_14[78] ? 7'h4e : _sels_3_T_175; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_177 = _T_14[77] ? 7'h4d : _sels_3_T_176; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_178 = _T_14[76] ? 7'h4c : _sels_3_T_177; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_179 = _T_14[75] ? 7'h4b : _sels_3_T_178; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_180 = _T_14[74] ? 7'h4a : _sels_3_T_179; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_181 = _T_14[73] ? 7'h49 : _sels_3_T_180; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_182 = _T_14[72] ? 7'h48 : _sels_3_T_181; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_183 = _T_14[71] ? 7'h47 : _sels_3_T_182; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_184 = _T_14[70] ? 7'h46 : _sels_3_T_183; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_185 = _T_14[69] ? 7'h45 : _sels_3_T_184; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_186 = _T_14[68] ? 7'h44 : _sels_3_T_185; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_187 = _T_14[67] ? 7'h43 : _sels_3_T_186; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_188 = _T_14[66] ? 7'h42 : _sels_3_T_187; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_189 = _T_14[65] ? 7'h41 : _sels_3_T_188; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_190 = _T_14[64] ? 7'h40 : _sels_3_T_189; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_191 = _T_14[63] ? 7'h3f : _sels_3_T_190; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_192 = _T_14[62] ? 7'h3e : _sels_3_T_191; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_193 = _T_14[61] ? 7'h3d : _sels_3_T_192; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_194 = _T_14[60] ? 7'h3c : _sels_3_T_193; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_195 = _T_14[59] ? 7'h3b : _sels_3_T_194; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_196 = _T_14[58] ? 7'h3a : _sels_3_T_195; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_197 = _T_14[57] ? 7'h39 : _sels_3_T_196; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_198 = _T_14[56] ? 7'h38 : _sels_3_T_197; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_199 = _T_14[55] ? 7'h37 : _sels_3_T_198; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_200 = _T_14[54] ? 7'h36 : _sels_3_T_199; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_201 = _T_14[53] ? 7'h35 : _sels_3_T_200; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_202 = _T_14[52] ? 7'h34 : _sels_3_T_201; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_203 = _T_14[51] ? 7'h33 : _sels_3_T_202; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_204 = _T_14[50] ? 7'h32 : _sels_3_T_203; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_205 = _T_14[49] ? 7'h31 : _sels_3_T_204; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_206 = _T_14[48] ? 7'h30 : _sels_3_T_205; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_207 = _T_14[47] ? 7'h2f : _sels_3_T_206; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_208 = _T_14[46] ? 7'h2e : _sels_3_T_207; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_209 = _T_14[45] ? 7'h2d : _sels_3_T_208; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_210 = _T_14[44] ? 7'h2c : _sels_3_T_209; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_211 = _T_14[43] ? 7'h2b : _sels_3_T_210; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_212 = _T_14[42] ? 7'h2a : _sels_3_T_211; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_213 = _T_14[41] ? 7'h29 : _sels_3_T_212; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_214 = _T_14[40] ? 7'h28 : _sels_3_T_213; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_215 = _T_14[39] ? 7'h27 : _sels_3_T_214; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_216 = _T_14[38] ? 7'h26 : _sels_3_T_215; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_217 = _T_14[37] ? 7'h25 : _sels_3_T_216; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_218 = _T_14[36] ? 7'h24 : _sels_3_T_217; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_219 = _T_14[35] ? 7'h23 : _sels_3_T_218; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_220 = _T_14[34] ? 7'h22 : _sels_3_T_219; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_221 = _T_14[33] ? 7'h21 : _sels_3_T_220; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_222 = _T_14[32] ? 7'h20 : _sels_3_T_221; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_223 = _T_14[31] ? 7'h1f : _sels_3_T_222; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_224 = _T_14[30] ? 7'h1e : _sels_3_T_223; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_225 = _T_14[29] ? 7'h1d : _sels_3_T_224; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_226 = _T_14[28] ? 7'h1c : _sels_3_T_225; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_227 = _T_14[27] ? 7'h1b : _sels_3_T_226; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_228 = _T_14[26] ? 7'h1a : _sels_3_T_227; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_229 = _T_14[25] ? 7'h19 : _sels_3_T_228; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_230 = _T_14[24] ? 7'h18 : _sels_3_T_229; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_231 = _T_14[23] ? 7'h17 : _sels_3_T_230; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_232 = _T_14[22] ? 7'h16 : _sels_3_T_231; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_233 = _T_14[21] ? 7'h15 : _sels_3_T_232; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_234 = _T_14[20] ? 7'h14 : _sels_3_T_233; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_235 = _T_14[19] ? 7'h13 : _sels_3_T_234; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_236 = _T_14[18] ? 7'h12 : _sels_3_T_235; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_237 = _T_14[17] ? 7'h11 : _sels_3_T_236; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_238 = _T_14[16] ? 7'h10 : _sels_3_T_237; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_239 = _T_14[15] ? 7'hf : _sels_3_T_238; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_240 = _T_14[14] ? 7'he : _sels_3_T_239; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_241 = _T_14[13] ? 7'hd : _sels_3_T_240; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_242 = _T_14[12] ? 7'hc : _sels_3_T_241; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_243 = _T_14[11] ? 7'hb : _sels_3_T_242; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_244 = _T_14[10] ? 7'ha : _sels_3_T_243; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_245 = _T_14[9] ? 7'h9 : _sels_3_T_244; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_246 = _T_14[8] ? 7'h8 : _sels_3_T_245; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_247 = _T_14[7] ? 7'h7 : _sels_3_T_246; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_248 = _T_14[6] ? 7'h6 : _sels_3_T_247; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_249 = _T_14[5] ? 7'h5 : _sels_3_T_248; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_250 = _T_14[4] ? 7'h4 : _sels_3_T_249; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_251 = _T_14[3] ? 7'h3 : _sels_3_T_250; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_252 = _T_14[2] ? 7'h2 : _sels_3_T_251; // @[Mux.scala 47:70]
  wire [6:0] _sels_3_T_253 = _T_14[1] ? 7'h1 : _sels_3_T_252; // @[Mux.scala 47:70]
  wire [6:0] rob_alloc_ids_3 = _T_14[0] ? 7'h0 : _sels_3_T_253; // @[Mux.scala 47:70]
  wire [127:0] _GEN_7172 = {{127'd0}, igen_3_io_fire}; // @[TestHarness.scala 187:45]
  wire [127:0] _T_74 = _GEN_7172 << rob_alloc_ids_3; // @[TestHarness.scala 187:45]
  wire [127:0] rob_allocs = _T_61 | _T_74; // @[TestHarness.scala 187:29]
  wire  _T_118 = io_from_noc_0_flit_ready & io_from_noc_0_flit_valid; // @[Decoupled.scala 51:35]
  wire  _T_119 = _T_118 & io_from_noc_0_flit_bits_tail; // @[TestHarness.scala 218:45]
  wire [15:0] out_payload_rob_idx = io_from_noc_0_flit_bits_payload[31:16]; // @[TestHarness.scala 194:51]
  wire [65535:0] _GEN_7173 = {{65535'd0}, _T_119}; // @[TestHarness.scala 218:66]
  wire [65535:0] _T_120 = _GEN_7173 << out_payload_rob_idx; // @[TestHarness.scala 218:66]
  wire  _T_165 = io_from_noc_1_flit_ready & io_from_noc_1_flit_valid; // @[Decoupled.scala 51:35]
  wire  _T_166 = _T_165 & io_from_noc_1_flit_bits_tail; // @[TestHarness.scala 218:45]
  wire [15:0] out_payload_1_rob_idx = io_from_noc_1_flit_bits_payload[31:16]; // @[TestHarness.scala 194:51]
  wire [65535:0] _GEN_7174 = {{65535'd0}, _T_166}; // @[TestHarness.scala 218:66]
  wire [65535:0] _T_167 = _GEN_7174 << out_payload_1_rob_idx; // @[TestHarness.scala 218:66]
  wire [65535:0] _T_168 = _T_120 | _T_167; // @[TestHarness.scala 218:27]
  wire  _T_212 = io_from_noc_2_flit_ready & io_from_noc_2_flit_valid; // @[Decoupled.scala 51:35]
  wire  _T_213 = _T_212 & io_from_noc_2_flit_bits_tail; // @[TestHarness.scala 218:45]
  wire [15:0] out_payload_2_rob_idx = io_from_noc_2_flit_bits_payload[31:16]; // @[TestHarness.scala 194:51]
  wire [65535:0] _GEN_7175 = {{65535'd0}, _T_213}; // @[TestHarness.scala 218:66]
  wire [65535:0] _T_214 = _GEN_7175 << out_payload_2_rob_idx; // @[TestHarness.scala 218:66]
  wire [65535:0] _T_215 = _T_168 | _T_214; // @[TestHarness.scala 218:27]
  wire  _T_259 = io_from_noc_3_flit_ready & io_from_noc_3_flit_valid; // @[Decoupled.scala 51:35]
  wire  _T_260 = _T_259 & io_from_noc_3_flit_bits_tail; // @[TestHarness.scala 218:45]
  wire [15:0] out_payload_3_rob_idx = io_from_noc_3_flit_bits_payload[31:16]; // @[TestHarness.scala 194:51]
  wire [65535:0] _GEN_7176 = {{65535'd0}, _T_260}; // @[TestHarness.scala 218:66]
  wire [65535:0] _T_261 = _GEN_7176 << out_payload_3_rob_idx; // @[TestHarness.scala 218:66]
  wire [65535:0] rob_frees = _T_215 | _T_261; // @[TestHarness.scala 218:27]
  wire  idle = rob_allocs == 128'h0 & rob_frees == 65536'h0; // @[TestHarness.scala 223:30]
  wire  _T_3 = ~reset; // @[TestHarness.scala 148:9]
  reg [31:0] rob_payload_0_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_0_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_0_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_1_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_1_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_1_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_2_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_2_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_2_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_3_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_3_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_3_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_4_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_4_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_4_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_5_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_5_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_5_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_6_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_6_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_6_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_7_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_7_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_7_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_8_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_8_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_8_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_9_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_9_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_9_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_10_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_10_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_10_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_11_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_11_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_11_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_12_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_12_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_12_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_13_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_13_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_13_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_14_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_14_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_14_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_15_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_15_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_15_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_16_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_16_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_16_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_17_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_17_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_17_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_18_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_18_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_18_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_19_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_19_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_19_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_20_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_20_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_20_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_21_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_21_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_21_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_22_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_22_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_22_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_23_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_23_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_23_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_24_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_24_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_24_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_25_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_25_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_25_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_26_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_26_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_26_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_27_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_27_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_27_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_28_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_28_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_28_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_29_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_29_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_29_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_30_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_30_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_30_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_31_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_31_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_31_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_32_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_32_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_32_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_33_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_33_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_33_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_34_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_34_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_34_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_35_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_35_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_35_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_36_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_36_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_36_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_37_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_37_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_37_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_38_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_38_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_38_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_39_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_39_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_39_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_40_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_40_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_40_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_41_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_41_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_41_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_42_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_42_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_42_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_43_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_43_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_43_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_44_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_44_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_44_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_45_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_45_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_45_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_46_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_46_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_46_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_47_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_47_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_47_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_48_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_48_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_48_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_49_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_49_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_49_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_50_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_50_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_50_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_51_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_51_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_51_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_52_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_52_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_52_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_53_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_53_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_53_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_54_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_54_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_54_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_55_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_55_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_55_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_56_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_56_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_56_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_57_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_57_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_57_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_58_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_58_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_58_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_59_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_59_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_59_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_60_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_60_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_60_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_61_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_61_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_61_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_62_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_62_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_62_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_63_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_63_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_63_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_64_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_64_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_64_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_65_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_65_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_65_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_66_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_66_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_66_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_67_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_67_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_67_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_68_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_68_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_68_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_69_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_69_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_69_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_70_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_70_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_70_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_71_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_71_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_71_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_72_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_72_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_72_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_73_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_73_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_73_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_74_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_74_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_74_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_75_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_75_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_75_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_76_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_76_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_76_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_77_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_77_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_77_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_78_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_78_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_78_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_79_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_79_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_79_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_80_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_80_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_80_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_81_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_81_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_81_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_82_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_82_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_82_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_83_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_83_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_83_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_84_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_84_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_84_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_85_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_85_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_85_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_86_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_86_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_86_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_87_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_87_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_87_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_88_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_88_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_88_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_89_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_89_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_89_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_90_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_90_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_90_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_91_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_91_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_91_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_92_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_92_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_92_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_93_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_93_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_93_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_94_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_94_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_94_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_95_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_95_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_95_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_96_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_96_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_96_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_97_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_97_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_97_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_98_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_98_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_98_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_99_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_99_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_99_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_100_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_100_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_100_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_101_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_101_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_101_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_102_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_102_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_102_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_103_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_103_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_103_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_104_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_104_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_104_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_105_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_105_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_105_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_106_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_106_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_106_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_107_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_107_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_107_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_108_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_108_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_108_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_109_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_109_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_109_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_110_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_110_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_110_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_111_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_111_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_111_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_112_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_112_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_112_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_113_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_113_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_113_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_114_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_114_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_114_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_115_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_115_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_115_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_116_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_116_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_116_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_117_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_117_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_117_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_118_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_118_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_118_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_119_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_119_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_119_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_120_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_120_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_120_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_121_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_121_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_121_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_122_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_122_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_122_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_123_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_123_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_123_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_124_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_124_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_124_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_125_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_125_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_125_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_126_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_126_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_126_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_127_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_127_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_127_flits_fired; // @[TestHarness.scala 150:24]
  reg [1:0] rob_egress_id_0; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_1; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_2; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_3; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_4; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_5; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_6; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_7; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_8; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_9; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_10; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_11; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_12; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_13; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_14; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_15; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_16; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_17; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_18; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_19; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_20; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_21; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_22; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_23; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_24; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_25; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_26; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_27; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_28; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_29; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_30; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_31; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_32; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_33; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_34; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_35; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_36; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_37; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_38; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_39; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_40; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_41; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_42; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_43; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_44; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_45; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_46; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_47; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_48; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_49; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_50; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_51; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_52; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_53; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_54; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_55; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_56; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_57; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_58; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_59; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_60; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_61; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_62; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_63; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_64; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_65; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_66; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_67; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_68; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_69; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_70; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_71; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_72; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_73; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_74; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_75; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_76; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_77; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_78; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_79; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_80; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_81; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_82; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_83; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_84; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_85; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_86; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_87; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_88; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_89; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_90; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_91; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_92; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_93; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_94; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_95; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_96; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_97; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_98; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_99; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_100; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_101; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_102; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_103; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_104; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_105; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_106; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_107; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_108; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_109; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_110; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_111; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_112; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_113; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_114; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_115; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_116; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_117; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_118; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_119; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_120; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_121; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_122; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_123; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_124; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_125; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_126; // @[TestHarness.scala 151:26]
  reg [1:0] rob_egress_id_127; // @[TestHarness.scala 151:26]
  reg [1:0] rob_ingress_id_0; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_1; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_2; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_3; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_4; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_5; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_6; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_7; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_8; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_9; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_10; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_11; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_12; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_13; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_14; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_15; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_16; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_17; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_18; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_19; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_20; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_21; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_22; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_23; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_24; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_25; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_26; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_27; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_28; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_29; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_30; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_31; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_32; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_33; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_34; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_35; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_36; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_37; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_38; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_39; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_40; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_41; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_42; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_43; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_44; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_45; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_46; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_47; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_48; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_49; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_50; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_51; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_52; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_53; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_54; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_55; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_56; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_57; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_58; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_59; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_60; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_61; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_62; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_63; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_64; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_65; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_66; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_67; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_68; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_69; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_70; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_71; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_72; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_73; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_74; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_75; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_76; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_77; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_78; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_79; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_80; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_81; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_82; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_83; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_84; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_85; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_86; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_87; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_88; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_89; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_90; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_91; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_92; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_93; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_94; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_95; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_96; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_97; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_98; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_99; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_100; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_101; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_102; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_103; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_104; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_105; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_106; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_107; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_108; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_109; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_110; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_111; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_112; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_113; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_114; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_115; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_116; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_117; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_118; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_119; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_120; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_121; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_122; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_123; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_124; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_125; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_126; // @[TestHarness.scala 152:27]
  reg [1:0] rob_ingress_id_127; // @[TestHarness.scala 152:27]
  reg [3:0] rob_n_flits_0; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_1; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_2; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_3; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_4; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_5; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_6; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_7; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_8; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_9; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_10; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_11; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_12; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_13; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_14; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_15; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_16; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_17; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_18; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_19; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_20; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_21; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_22; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_23; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_24; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_25; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_26; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_27; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_28; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_29; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_30; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_31; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_32; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_33; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_34; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_35; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_36; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_37; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_38; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_39; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_40; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_41; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_42; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_43; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_44; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_45; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_46; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_47; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_48; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_49; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_50; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_51; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_52; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_53; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_54; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_55; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_56; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_57; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_58; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_59; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_60; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_61; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_62; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_63; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_64; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_65; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_66; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_67; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_68; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_69; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_70; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_71; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_72; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_73; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_74; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_75; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_76; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_77; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_78; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_79; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_80; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_81; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_82; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_83; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_84; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_85; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_86; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_87; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_88; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_89; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_90; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_91; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_92; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_93; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_94; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_95; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_96; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_97; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_98; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_99; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_100; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_101; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_102; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_103; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_104; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_105; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_106; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_107; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_108; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_109; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_110; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_111; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_112; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_113; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_114; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_115; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_116; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_117; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_118; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_119; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_120; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_121; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_122; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_123; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_124; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_125; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_126; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_127; // @[TestHarness.scala 153:24]
  reg [3:0] rob_flits_returned_0; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_1; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_2; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_3; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_4; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_5; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_6; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_7; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_8; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_9; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_10; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_11; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_12; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_13; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_14; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_15; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_16; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_17; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_18; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_19; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_20; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_21; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_22; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_23; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_24; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_25; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_26; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_27; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_28; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_29; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_30; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_31; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_32; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_33; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_34; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_35; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_36; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_37; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_38; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_39; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_40; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_41; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_42; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_43; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_44; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_45; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_46; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_47; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_48; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_49; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_50; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_51; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_52; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_53; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_54; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_55; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_56; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_57; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_58; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_59; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_60; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_61; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_62; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_63; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_64; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_65; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_66; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_67; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_68; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_69; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_70; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_71; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_72; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_73; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_74; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_75; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_76; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_77; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_78; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_79; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_80; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_81; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_82; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_83; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_84; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_85; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_86; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_87; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_88; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_89; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_90; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_91; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_92; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_93; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_94; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_95; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_96; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_97; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_98; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_99; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_100; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_101; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_102; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_103; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_104; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_105; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_106; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_107; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_108; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_109; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_110; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_111; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_112; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_113; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_114; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_115; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_116; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_117; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_118; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_119; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_120; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_121; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_122; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_123; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_124; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_125; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_126; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_127; // @[TestHarness.scala 154:31]
  reg [63:0] rob_tscs_0; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_1; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_2; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_3; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_4; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_5; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_6; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_7; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_8; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_9; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_10; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_11; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_12; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_13; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_14; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_15; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_16; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_17; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_18; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_19; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_20; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_21; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_22; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_23; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_24; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_25; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_26; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_27; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_28; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_29; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_30; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_31; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_32; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_33; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_34; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_35; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_36; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_37; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_38; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_39; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_40; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_41; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_42; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_43; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_44; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_45; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_46; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_47; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_48; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_49; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_50; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_51; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_52; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_53; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_54; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_55; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_56; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_57; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_58; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_59; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_60; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_61; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_62; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_63; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_64; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_65; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_66; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_67; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_68; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_69; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_70; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_71; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_72; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_73; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_74; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_75; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_76; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_77; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_78; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_79; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_80; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_81; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_82; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_83; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_84; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_85; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_86; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_87; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_88; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_89; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_90; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_91; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_92; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_93; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_94; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_95; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_96; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_97; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_98; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_99; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_100; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_101; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_102; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_103; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_104; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_105; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_106; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_107; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_108; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_109; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_110; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_111; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_112; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_113; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_114; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_115; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_116; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_117; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_118; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_119; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_120; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_121; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_122; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_123; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_124; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_125; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_126; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_127; // @[TestHarness.scala 155:21]
  wire  rob_alloc_fires_0 = _T_5 != 128'h0; // @[TestHarness.scala 30:24]
  wire  rob_alloc_fires_1 = _T_8 != 128'h0; // @[TestHarness.scala 30:24]
  wire  rob_alloc_fires_2 = _T_11 != 128'h0; // @[TestHarness.scala 30:24]
  wire  rob_alloc_fires_3 = _T_14 != 128'h0; // @[TestHarness.scala 30:24]
  wire [127:0] _rob_alloc_avail_T = rob_valids >> rob_alloc_ids_0; // @[TestHarness.scala 162:61]
  wire  rob_alloc_avail_0 = ~_rob_alloc_avail_T[0]; // @[TestHarness.scala 162:50]
  wire [127:0] _rob_alloc_avail_T_2 = rob_valids >> rob_alloc_ids_1; // @[TestHarness.scala 162:61]
  wire  rob_alloc_avail_1 = ~_rob_alloc_avail_T_2[0]; // @[TestHarness.scala 162:50]
  wire [127:0] _rob_alloc_avail_T_4 = rob_valids >> rob_alloc_ids_2; // @[TestHarness.scala 162:61]
  wire  rob_alloc_avail_2 = ~_rob_alloc_avail_T_4[0]; // @[TestHarness.scala 162:50]
  wire [127:0] _rob_alloc_avail_T_6 = rob_valids >> rob_alloc_ids_3; // @[TestHarness.scala 162:61]
  wire  rob_alloc_avail_3 = ~_rob_alloc_avail_T_6[0]; // @[TestHarness.scala 162:50]
  wire  success = txs >= 32'hc350 & rob_valids == 128'h0; // @[TestHarness.scala 163:35]
  reg  io_success_REG; // @[TestHarness.scala 164:24]
  wire  _igen_io_rob_ready_T_1 = tsc >= 32'ha; // @[TestHarness.scala 175:11]
  wire  _igen_io_rob_ready_T_2 = rob_alloc_avail_0 & rob_alloc_fires_0 & _igen_io_rob_ready_T_1; // @[TestHarness.scala 174:72]
  wire [63:0] _rob_payload_WIRE_1 = igen_io_out_bits_payload; // @[TestHarness.scala 179:{72,72}]
  wire [31:0] _GEN_1 = 7'h0 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_0_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_2 = 7'h1 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_1_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_3 = 7'h2 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_2_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_4 = 7'h3 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_3_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_5 = 7'h4 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_4_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_6 = 7'h5 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_5_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_7 = 7'h6 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_6_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_8 = 7'h7 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_7_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_9 = 7'h8 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_8_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_10 = 7'h9 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_9_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_11 = 7'ha == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_10_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_12 = 7'hb == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_11_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_13 = 7'hc == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_12_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_14 = 7'hd == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_13_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_15 = 7'he == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_14_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_16 = 7'hf == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_15_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_17 = 7'h10 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_16_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_18 = 7'h11 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_17_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_19 = 7'h12 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_18_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_20 = 7'h13 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_19_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_21 = 7'h14 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_20_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_22 = 7'h15 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_21_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_23 = 7'h16 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_22_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_24 = 7'h17 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_23_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_25 = 7'h18 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_24_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_26 = 7'h19 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_25_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_27 = 7'h1a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_26_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_28 = 7'h1b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_27_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_29 = 7'h1c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_28_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_30 = 7'h1d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_29_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_31 = 7'h1e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_30_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_32 = 7'h1f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_31_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_33 = 7'h20 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_32_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_34 = 7'h21 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_33_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_35 = 7'h22 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_34_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_36 = 7'h23 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_35_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_37 = 7'h24 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_36_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_38 = 7'h25 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_37_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_39 = 7'h26 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_38_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_40 = 7'h27 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_39_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_41 = 7'h28 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_40_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_42 = 7'h29 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_41_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_43 = 7'h2a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_42_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_44 = 7'h2b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_43_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_45 = 7'h2c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_44_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_46 = 7'h2d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_45_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_47 = 7'h2e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_46_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_48 = 7'h2f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_47_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_49 = 7'h30 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_48_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_50 = 7'h31 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_49_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_51 = 7'h32 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_50_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_52 = 7'h33 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_51_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_53 = 7'h34 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_52_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_54 = 7'h35 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_53_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_55 = 7'h36 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_54_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_56 = 7'h37 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_55_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_57 = 7'h38 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_56_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_58 = 7'h39 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_57_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_59 = 7'h3a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_58_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_60 = 7'h3b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_59_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_61 = 7'h3c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_60_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_62 = 7'h3d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_61_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_63 = 7'h3e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_62_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_64 = 7'h3f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_63_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_65 = 7'h40 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_64_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_66 = 7'h41 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_65_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_67 = 7'h42 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_66_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_68 = 7'h43 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_67_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_69 = 7'h44 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_68_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_70 = 7'h45 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_69_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_71 = 7'h46 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_70_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_72 = 7'h47 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_71_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_73 = 7'h48 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_72_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_74 = 7'h49 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_73_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_75 = 7'h4a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_74_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_76 = 7'h4b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_75_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_77 = 7'h4c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_76_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_78 = 7'h4d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_77_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_79 = 7'h4e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_78_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_80 = 7'h4f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_79_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_81 = 7'h50 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_80_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_82 = 7'h51 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_81_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_83 = 7'h52 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_82_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_84 = 7'h53 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_83_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_85 = 7'h54 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_84_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_86 = 7'h55 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_85_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_87 = 7'h56 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_86_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_88 = 7'h57 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_87_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_89 = 7'h58 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_88_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_90 = 7'h59 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_89_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_91 = 7'h5a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_90_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_92 = 7'h5b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_91_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_93 = 7'h5c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_92_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_94 = 7'h5d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_93_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_95 = 7'h5e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_94_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_96 = 7'h5f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_95_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_97 = 7'h60 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_96_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_98 = 7'h61 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_97_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_99 = 7'h62 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_98_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_100 = 7'h63 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_99_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_101 = 7'h64 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_100_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_102 = 7'h65 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_101_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_103 = 7'h66 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_102_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_104 = 7'h67 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_103_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_105 = 7'h68 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_104_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_106 = 7'h69 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_105_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_107 = 7'h6a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_106_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_108 = 7'h6b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_107_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_109 = 7'h6c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_108_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_110 = 7'h6d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_109_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_111 = 7'h6e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_110_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_112 = 7'h6f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_111_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_113 = 7'h70 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_112_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_114 = 7'h71 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_113_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_115 = 7'h72 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_114_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_116 = 7'h73 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_115_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_117 = 7'h74 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_116_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_118 = 7'h75 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_117_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_119 = 7'h76 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_118_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_120 = 7'h77 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_119_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_121 = 7'h78 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_120_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_122 = 7'h79 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_121_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_123 = 7'h7a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_122_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_124 = 7'h7b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_123_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_125 = 7'h7c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_124_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_126 = 7'h7d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_125_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_127 = 7'h7e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_126_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_128 = 7'h7f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_127_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_129 = 7'h0 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_0_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_130 = 7'h1 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_1_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_131 = 7'h2 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_2_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_132 = 7'h3 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_3_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_133 = 7'h4 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_4_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_134 = 7'h5 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_5_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_135 = 7'h6 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_6_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_136 = 7'h7 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_7_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_137 = 7'h8 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_8_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_138 = 7'h9 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_9_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_139 = 7'ha == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_10_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_140 = 7'hb == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_11_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_141 = 7'hc == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_12_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_142 = 7'hd == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_13_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_143 = 7'he == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_14_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_144 = 7'hf == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_15_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_145 = 7'h10 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_16_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_146 = 7'h11 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_17_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_147 = 7'h12 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_18_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_148 = 7'h13 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_19_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_149 = 7'h14 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_20_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_150 = 7'h15 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_21_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_151 = 7'h16 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_22_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_152 = 7'h17 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_23_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_153 = 7'h18 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_24_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_154 = 7'h19 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_25_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_155 = 7'h1a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_26_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_156 = 7'h1b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_27_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_157 = 7'h1c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_28_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_158 = 7'h1d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_29_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_159 = 7'h1e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_30_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_160 = 7'h1f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_31_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_161 = 7'h20 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_32_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_162 = 7'h21 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_33_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_163 = 7'h22 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_34_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_164 = 7'h23 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_35_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_165 = 7'h24 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_36_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_166 = 7'h25 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_37_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_167 = 7'h26 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_38_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_168 = 7'h27 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_39_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_169 = 7'h28 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_40_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_170 = 7'h29 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_41_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_171 = 7'h2a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_42_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_172 = 7'h2b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_43_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_173 = 7'h2c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_44_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_174 = 7'h2d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_45_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_175 = 7'h2e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_46_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_176 = 7'h2f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_47_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_177 = 7'h30 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_48_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_178 = 7'h31 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_49_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_179 = 7'h32 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_50_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_180 = 7'h33 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_51_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_181 = 7'h34 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_52_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_182 = 7'h35 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_53_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_183 = 7'h36 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_54_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_184 = 7'h37 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_55_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_185 = 7'h38 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_56_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_186 = 7'h39 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_57_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_187 = 7'h3a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_58_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_188 = 7'h3b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_59_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_189 = 7'h3c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_60_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_190 = 7'h3d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_61_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_191 = 7'h3e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_62_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_192 = 7'h3f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_63_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_193 = 7'h40 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_64_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_194 = 7'h41 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_65_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_195 = 7'h42 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_66_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_196 = 7'h43 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_67_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_197 = 7'h44 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_68_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_198 = 7'h45 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_69_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_199 = 7'h46 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_70_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_200 = 7'h47 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_71_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_201 = 7'h48 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_72_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_202 = 7'h49 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_73_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_203 = 7'h4a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_74_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_204 = 7'h4b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_75_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_205 = 7'h4c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_76_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_206 = 7'h4d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_77_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_207 = 7'h4e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_78_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_208 = 7'h4f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_79_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_209 = 7'h50 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_80_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_210 = 7'h51 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_81_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_211 = 7'h52 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_82_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_212 = 7'h53 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_83_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_213 = 7'h54 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_84_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_214 = 7'h55 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_85_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_215 = 7'h56 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_86_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_216 = 7'h57 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_87_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_217 = 7'h58 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_88_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_218 = 7'h59 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_89_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_219 = 7'h5a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_90_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_220 = 7'h5b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_91_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_221 = 7'h5c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_92_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_222 = 7'h5d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_93_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_223 = 7'h5e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_94_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_224 = 7'h5f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_95_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_225 = 7'h60 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_96_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_226 = 7'h61 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_97_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_227 = 7'h62 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_98_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_228 = 7'h63 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_99_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_229 = 7'h64 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_100_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_230 = 7'h65 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_101_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_231 = 7'h66 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_102_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_232 = 7'h67 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_103_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_233 = 7'h68 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_104_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_234 = 7'h69 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_105_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_235 = 7'h6a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_106_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_236 = 7'h6b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_107_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_237 = 7'h6c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_108_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_238 = 7'h6d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_109_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_239 = 7'h6e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_110_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_240 = 7'h6f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_111_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_241 = 7'h70 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_112_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_242 = 7'h71 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_113_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_243 = 7'h72 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_114_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_244 = 7'h73 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_115_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_245 = 7'h74 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_116_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_246 = 7'h75 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_117_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_247 = 7'h76 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_118_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_248 = 7'h77 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_119_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_249 = 7'h78 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_120_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_250 = 7'h79 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_121_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_251 = 7'h7a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_122_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_252 = 7'h7b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_123_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_253 = 7'h7c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_124_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_254 = 7'h7d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_125_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_255 = 7'h7e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_126_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_256 = 7'h7f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_127_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_257 = 7'h0 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_0_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_258 = 7'h1 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_1_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_259 = 7'h2 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_2_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_260 = 7'h3 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_3_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_261 = 7'h4 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_4_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_262 = 7'h5 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_5_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_263 = 7'h6 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_6_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_264 = 7'h7 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_7_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_265 = 7'h8 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_8_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_266 = 7'h9 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_9_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_267 = 7'ha == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_10_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_268 = 7'hb == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_11_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_269 = 7'hc == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_12_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_270 = 7'hd == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_13_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_271 = 7'he == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_14_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_272 = 7'hf == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_15_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_273 = 7'h10 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_16_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_274 = 7'h11 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_17_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_275 = 7'h12 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_18_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_276 = 7'h13 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_19_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_277 = 7'h14 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_20_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_278 = 7'h15 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_21_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_279 = 7'h16 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_22_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_280 = 7'h17 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_23_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_281 = 7'h18 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_24_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_282 = 7'h19 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_25_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_283 = 7'h1a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_26_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_284 = 7'h1b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_27_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_285 = 7'h1c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_28_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_286 = 7'h1d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_29_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_287 = 7'h1e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_30_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_288 = 7'h1f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_31_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_289 = 7'h20 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_32_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_290 = 7'h21 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_33_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_291 = 7'h22 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_34_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_292 = 7'h23 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_35_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_293 = 7'h24 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_36_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_294 = 7'h25 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_37_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_295 = 7'h26 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_38_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_296 = 7'h27 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_39_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_297 = 7'h28 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_40_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_298 = 7'h29 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_41_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_299 = 7'h2a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_42_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_300 = 7'h2b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_43_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_301 = 7'h2c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_44_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_302 = 7'h2d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_45_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_303 = 7'h2e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_46_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_304 = 7'h2f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_47_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_305 = 7'h30 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_48_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_306 = 7'h31 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_49_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_307 = 7'h32 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_50_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_308 = 7'h33 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_51_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_309 = 7'h34 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_52_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_310 = 7'h35 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_53_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_311 = 7'h36 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_54_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_312 = 7'h37 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_55_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_313 = 7'h38 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_56_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_314 = 7'h39 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_57_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_315 = 7'h3a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_58_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_316 = 7'h3b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_59_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_317 = 7'h3c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_60_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_318 = 7'h3d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_61_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_319 = 7'h3e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_62_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_320 = 7'h3f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_63_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_321 = 7'h40 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_64_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_322 = 7'h41 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_65_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_323 = 7'h42 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_66_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_324 = 7'h43 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_67_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_325 = 7'h44 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_68_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_326 = 7'h45 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_69_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_327 = 7'h46 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_70_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_328 = 7'h47 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_71_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_329 = 7'h48 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_72_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_330 = 7'h49 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_73_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_331 = 7'h4a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_74_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_332 = 7'h4b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_75_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_333 = 7'h4c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_76_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_334 = 7'h4d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_77_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_335 = 7'h4e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_78_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_336 = 7'h4f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_79_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_337 = 7'h50 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_80_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_338 = 7'h51 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_81_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_339 = 7'h52 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_82_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_340 = 7'h53 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_83_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_341 = 7'h54 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_84_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_342 = 7'h55 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_85_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_343 = 7'h56 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_86_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_344 = 7'h57 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_87_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_345 = 7'h58 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_88_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_346 = 7'h59 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_89_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_347 = 7'h5a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_90_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_348 = 7'h5b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_91_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_349 = 7'h5c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_92_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_350 = 7'h5d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_93_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_351 = 7'h5e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_94_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_352 = 7'h5f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_95_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_353 = 7'h60 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_96_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_354 = 7'h61 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_97_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_355 = 7'h62 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_98_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_356 = 7'h63 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_99_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_357 = 7'h64 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_100_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_358 = 7'h65 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_101_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_359 = 7'h66 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_102_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_360 = 7'h67 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_103_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_361 = 7'h68 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_104_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_362 = 7'h69 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_105_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_363 = 7'h6a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_106_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_364 = 7'h6b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_107_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_365 = 7'h6c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_108_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_366 = 7'h6d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_109_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_367 = 7'h6e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_110_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_368 = 7'h6f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_111_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_369 = 7'h70 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_112_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_370 = 7'h71 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_113_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_371 = 7'h72 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_114_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_372 = 7'h73 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_115_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_373 = 7'h74 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_116_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_374 = 7'h75 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_117_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_375 = 7'h76 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_118_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_376 = 7'h77 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_119_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_377 = 7'h78 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_120_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_378 = 7'h79 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_121_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_379 = 7'h7a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_122_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_380 = 7'h7b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_123_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_381 = 7'h7c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_124_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_382 = 7'h7d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_125_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_383 = 7'h7e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_126_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_384 = 7'h7f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_127_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [1:0] _rob_egress_id_T_23 = igen_io_out_bits_egress_id; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_385 = 7'h0 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_0; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_386 = 7'h1 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_1; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_387 = 7'h2 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_2; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_388 = 7'h3 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_3; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_389 = 7'h4 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_4; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_390 = 7'h5 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_5; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_391 = 7'h6 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_6; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_392 = 7'h7 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_7; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_393 = 7'h8 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_8; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_394 = 7'h9 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_9; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_395 = 7'ha == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_10; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_396 = 7'hb == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_11; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_397 = 7'hc == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_12; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_398 = 7'hd == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_13; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_399 = 7'he == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_14; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_400 = 7'hf == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_15; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_401 = 7'h10 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_16; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_402 = 7'h11 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_17; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_403 = 7'h12 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_18; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_404 = 7'h13 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_19; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_405 = 7'h14 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_20; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_406 = 7'h15 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_21; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_407 = 7'h16 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_22; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_408 = 7'h17 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_23; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_409 = 7'h18 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_24; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_410 = 7'h19 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_25; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_411 = 7'h1a == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_26; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_412 = 7'h1b == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_27; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_413 = 7'h1c == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_28; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_414 = 7'h1d == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_29; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_415 = 7'h1e == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_30; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_416 = 7'h1f == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_31; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_417 = 7'h20 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_32; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_418 = 7'h21 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_33; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_419 = 7'h22 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_34; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_420 = 7'h23 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_35; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_421 = 7'h24 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_36; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_422 = 7'h25 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_37; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_423 = 7'h26 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_38; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_424 = 7'h27 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_39; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_425 = 7'h28 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_40; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_426 = 7'h29 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_41; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_427 = 7'h2a == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_42; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_428 = 7'h2b == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_43; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_429 = 7'h2c == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_44; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_430 = 7'h2d == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_45; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_431 = 7'h2e == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_46; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_432 = 7'h2f == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_47; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_433 = 7'h30 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_48; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_434 = 7'h31 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_49; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_435 = 7'h32 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_50; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_436 = 7'h33 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_51; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_437 = 7'h34 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_52; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_438 = 7'h35 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_53; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_439 = 7'h36 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_54; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_440 = 7'h37 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_55; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_441 = 7'h38 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_56; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_442 = 7'h39 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_57; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_443 = 7'h3a == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_58; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_444 = 7'h3b == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_59; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_445 = 7'h3c == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_60; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_446 = 7'h3d == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_61; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_447 = 7'h3e == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_62; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_448 = 7'h3f == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_63; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_449 = 7'h40 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_64; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_450 = 7'h41 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_65; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_451 = 7'h42 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_66; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_452 = 7'h43 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_67; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_453 = 7'h44 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_68; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_454 = 7'h45 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_69; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_455 = 7'h46 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_70; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_456 = 7'h47 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_71; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_457 = 7'h48 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_72; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_458 = 7'h49 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_73; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_459 = 7'h4a == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_74; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_460 = 7'h4b == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_75; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_461 = 7'h4c == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_76; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_462 = 7'h4d == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_77; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_463 = 7'h4e == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_78; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_464 = 7'h4f == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_79; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_465 = 7'h50 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_80; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_466 = 7'h51 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_81; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_467 = 7'h52 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_82; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_468 = 7'h53 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_83; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_469 = 7'h54 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_84; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_470 = 7'h55 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_85; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_471 = 7'h56 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_86; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_472 = 7'h57 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_87; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_473 = 7'h58 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_88; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_474 = 7'h59 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_89; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_475 = 7'h5a == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_90; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_476 = 7'h5b == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_91; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_477 = 7'h5c == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_92; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_478 = 7'h5d == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_93; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_479 = 7'h5e == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_94; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_480 = 7'h5f == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_95; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_481 = 7'h60 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_96; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_482 = 7'h61 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_97; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_483 = 7'h62 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_98; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_484 = 7'h63 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_99; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_485 = 7'h64 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_100; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_486 = 7'h65 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_101; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_487 = 7'h66 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_102; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_488 = 7'h67 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_103; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_489 = 7'h68 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_104; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_490 = 7'h69 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_105; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_491 = 7'h6a == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_106; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_492 = 7'h6b == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_107; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_493 = 7'h6c == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_108; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_494 = 7'h6d == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_109; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_495 = 7'h6e == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_110; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_496 = 7'h6f == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_111; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_497 = 7'h70 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_112; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_498 = 7'h71 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_113; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_499 = 7'h72 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_114; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_500 = 7'h73 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_115; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_501 = 7'h74 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_116; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_502 = 7'h75 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_117; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_503 = 7'h76 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_118; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_504 = 7'h77 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_119; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_505 = 7'h78 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_120; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_506 = 7'h79 == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_121; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_507 = 7'h7a == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_122; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_508 = 7'h7b == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_123; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_509 = 7'h7c == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_124; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_510 = 7'h7d == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_125; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_511 = 7'h7e == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_126; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_512 = 7'h7f == rob_alloc_ids_0 ? _rob_egress_id_T_23 : rob_egress_id_127; // @[TestHarness.scala 151:26 180:{36,36}]
  wire [1:0] _GEN_513 = 7'h0 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_0; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_514 = 7'h1 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_1; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_515 = 7'h2 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_2; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_516 = 7'h3 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_3; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_517 = 7'h4 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_4; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_518 = 7'h5 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_5; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_519 = 7'h6 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_6; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_520 = 7'h7 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_7; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_521 = 7'h8 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_8; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_522 = 7'h9 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_9; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_523 = 7'ha == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_10; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_524 = 7'hb == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_11; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_525 = 7'hc == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_12; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_526 = 7'hd == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_13; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_527 = 7'he == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_14; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_528 = 7'hf == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_15; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_529 = 7'h10 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_16; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_530 = 7'h11 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_17; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_531 = 7'h12 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_18; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_532 = 7'h13 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_19; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_533 = 7'h14 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_20; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_534 = 7'h15 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_21; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_535 = 7'h16 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_22; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_536 = 7'h17 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_23; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_537 = 7'h18 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_24; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_538 = 7'h19 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_25; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_539 = 7'h1a == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_26; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_540 = 7'h1b == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_27; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_541 = 7'h1c == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_28; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_542 = 7'h1d == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_29; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_543 = 7'h1e == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_30; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_544 = 7'h1f == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_31; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_545 = 7'h20 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_32; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_546 = 7'h21 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_33; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_547 = 7'h22 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_34; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_548 = 7'h23 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_35; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_549 = 7'h24 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_36; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_550 = 7'h25 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_37; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_551 = 7'h26 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_38; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_552 = 7'h27 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_39; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_553 = 7'h28 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_40; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_554 = 7'h29 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_41; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_555 = 7'h2a == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_42; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_556 = 7'h2b == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_43; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_557 = 7'h2c == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_44; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_558 = 7'h2d == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_45; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_559 = 7'h2e == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_46; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_560 = 7'h2f == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_47; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_561 = 7'h30 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_48; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_562 = 7'h31 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_49; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_563 = 7'h32 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_50; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_564 = 7'h33 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_51; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_565 = 7'h34 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_52; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_566 = 7'h35 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_53; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_567 = 7'h36 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_54; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_568 = 7'h37 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_55; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_569 = 7'h38 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_56; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_570 = 7'h39 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_57; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_571 = 7'h3a == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_58; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_572 = 7'h3b == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_59; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_573 = 7'h3c == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_60; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_574 = 7'h3d == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_61; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_575 = 7'h3e == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_62; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_576 = 7'h3f == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_63; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_577 = 7'h40 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_64; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_578 = 7'h41 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_65; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_579 = 7'h42 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_66; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_580 = 7'h43 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_67; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_581 = 7'h44 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_68; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_582 = 7'h45 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_69; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_583 = 7'h46 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_70; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_584 = 7'h47 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_71; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_585 = 7'h48 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_72; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_586 = 7'h49 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_73; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_587 = 7'h4a == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_74; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_588 = 7'h4b == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_75; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_589 = 7'h4c == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_76; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_590 = 7'h4d == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_77; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_591 = 7'h4e == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_78; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_592 = 7'h4f == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_79; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_593 = 7'h50 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_80; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_594 = 7'h51 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_81; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_595 = 7'h52 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_82; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_596 = 7'h53 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_83; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_597 = 7'h54 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_84; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_598 = 7'h55 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_85; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_599 = 7'h56 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_86; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_600 = 7'h57 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_87; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_601 = 7'h58 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_88; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_602 = 7'h59 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_89; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_603 = 7'h5a == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_90; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_604 = 7'h5b == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_91; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_605 = 7'h5c == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_92; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_606 = 7'h5d == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_93; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_607 = 7'h5e == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_94; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_608 = 7'h5f == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_95; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_609 = 7'h60 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_96; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_610 = 7'h61 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_97; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_611 = 7'h62 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_98; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_612 = 7'h63 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_99; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_613 = 7'h64 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_100; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_614 = 7'h65 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_101; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_615 = 7'h66 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_102; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_616 = 7'h67 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_103; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_617 = 7'h68 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_104; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_618 = 7'h69 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_105; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_619 = 7'h6a == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_106; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_620 = 7'h6b == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_107; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_621 = 7'h6c == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_108; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_622 = 7'h6d == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_109; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_623 = 7'h6e == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_110; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_624 = 7'h6f == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_111; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_625 = 7'h70 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_112; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_626 = 7'h71 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_113; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_627 = 7'h72 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_114; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_628 = 7'h73 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_115; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_629 = 7'h74 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_116; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_630 = 7'h75 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_117; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_631 = 7'h76 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_118; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_632 = 7'h77 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_119; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_633 = 7'h78 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_120; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_634 = 7'h79 == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_121; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_635 = 7'h7a == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_122; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_636 = 7'h7b == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_123; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_637 = 7'h7c == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_124; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_638 = 7'h7d == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_125; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_639 = 7'h7e == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_126; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [1:0] _GEN_640 = 7'h7f == rob_alloc_ids_0 ? 2'h0 : rob_ingress_id_127; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [3:0] _rob_n_flits_T_27 = igen_io_n_flits; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_641 = 7'h0 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_0; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_642 = 7'h1 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_1; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_643 = 7'h2 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_2; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_644 = 7'h3 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_3; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_645 = 7'h4 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_4; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_646 = 7'h5 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_5; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_647 = 7'h6 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_6; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_648 = 7'h7 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_7; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_649 = 7'h8 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_8; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_650 = 7'h9 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_9; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_651 = 7'ha == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_10; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_652 = 7'hb == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_11; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_653 = 7'hc == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_12; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_654 = 7'hd == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_13; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_655 = 7'he == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_14; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_656 = 7'hf == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_15; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_657 = 7'h10 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_16; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_658 = 7'h11 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_17; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_659 = 7'h12 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_18; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_660 = 7'h13 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_19; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_661 = 7'h14 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_20; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_662 = 7'h15 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_21; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_663 = 7'h16 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_22; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_664 = 7'h17 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_23; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_665 = 7'h18 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_24; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_666 = 7'h19 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_25; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_667 = 7'h1a == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_26; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_668 = 7'h1b == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_27; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_669 = 7'h1c == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_28; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_670 = 7'h1d == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_29; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_671 = 7'h1e == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_30; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_672 = 7'h1f == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_31; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_673 = 7'h20 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_32; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_674 = 7'h21 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_33; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_675 = 7'h22 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_34; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_676 = 7'h23 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_35; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_677 = 7'h24 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_36; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_678 = 7'h25 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_37; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_679 = 7'h26 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_38; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_680 = 7'h27 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_39; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_681 = 7'h28 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_40; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_682 = 7'h29 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_41; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_683 = 7'h2a == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_42; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_684 = 7'h2b == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_43; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_685 = 7'h2c == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_44; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_686 = 7'h2d == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_45; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_687 = 7'h2e == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_46; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_688 = 7'h2f == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_47; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_689 = 7'h30 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_48; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_690 = 7'h31 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_49; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_691 = 7'h32 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_50; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_692 = 7'h33 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_51; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_693 = 7'h34 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_52; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_694 = 7'h35 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_53; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_695 = 7'h36 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_54; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_696 = 7'h37 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_55; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_697 = 7'h38 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_56; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_698 = 7'h39 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_57; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_699 = 7'h3a == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_58; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_700 = 7'h3b == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_59; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_701 = 7'h3c == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_60; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_702 = 7'h3d == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_61; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_703 = 7'h3e == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_62; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_704 = 7'h3f == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_63; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_705 = 7'h40 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_64; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_706 = 7'h41 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_65; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_707 = 7'h42 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_66; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_708 = 7'h43 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_67; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_709 = 7'h44 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_68; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_710 = 7'h45 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_69; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_711 = 7'h46 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_70; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_712 = 7'h47 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_71; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_713 = 7'h48 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_72; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_714 = 7'h49 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_73; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_715 = 7'h4a == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_74; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_716 = 7'h4b == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_75; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_717 = 7'h4c == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_76; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_718 = 7'h4d == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_77; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_719 = 7'h4e == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_78; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_720 = 7'h4f == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_79; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_721 = 7'h50 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_80; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_722 = 7'h51 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_81; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_723 = 7'h52 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_82; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_724 = 7'h53 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_83; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_725 = 7'h54 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_84; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_726 = 7'h55 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_85; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_727 = 7'h56 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_86; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_728 = 7'h57 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_87; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_729 = 7'h58 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_88; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_730 = 7'h59 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_89; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_731 = 7'h5a == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_90; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_732 = 7'h5b == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_91; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_733 = 7'h5c == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_92; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_734 = 7'h5d == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_93; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_735 = 7'h5e == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_94; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_736 = 7'h5f == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_95; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_737 = 7'h60 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_96; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_738 = 7'h61 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_97; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_739 = 7'h62 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_98; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_740 = 7'h63 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_99; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_741 = 7'h64 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_100; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_742 = 7'h65 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_101; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_743 = 7'h66 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_102; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_744 = 7'h67 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_103; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_745 = 7'h68 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_104; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_746 = 7'h69 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_105; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_747 = 7'h6a == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_106; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_748 = 7'h6b == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_107; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_749 = 7'h6c == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_108; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_750 = 7'h6d == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_109; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_751 = 7'h6e == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_110; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_752 = 7'h6f == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_111; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_753 = 7'h70 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_112; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_754 = 7'h71 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_113; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_755 = 7'h72 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_114; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_756 = 7'h73 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_115; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_757 = 7'h74 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_116; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_758 = 7'h75 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_117; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_759 = 7'h76 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_118; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_760 = 7'h77 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_119; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_761 = 7'h78 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_120; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_762 = 7'h79 == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_121; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_763 = 7'h7a == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_122; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_764 = 7'h7b == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_123; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_765 = 7'h7c == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_124; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_766 = 7'h7d == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_125; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_767 = 7'h7e == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_126; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_768 = 7'h7f == rob_alloc_ids_0 ? _rob_n_flits_T_27 : rob_n_flits_127; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_769 = 7'h0 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_0; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_770 = 7'h1 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_1; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_771 = 7'h2 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_2; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_772 = 7'h3 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_3; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_773 = 7'h4 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_4; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_774 = 7'h5 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_5; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_775 = 7'h6 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_6; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_776 = 7'h7 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_7; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_777 = 7'h8 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_8; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_778 = 7'h9 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_9; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_779 = 7'ha == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_10; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_780 = 7'hb == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_11; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_781 = 7'hc == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_12; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_782 = 7'hd == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_13; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_783 = 7'he == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_14; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_784 = 7'hf == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_15; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_785 = 7'h10 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_16; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_786 = 7'h11 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_17; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_787 = 7'h12 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_18; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_788 = 7'h13 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_19; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_789 = 7'h14 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_20; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_790 = 7'h15 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_21; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_791 = 7'h16 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_22; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_792 = 7'h17 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_23; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_793 = 7'h18 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_24; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_794 = 7'h19 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_25; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_795 = 7'h1a == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_26; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_796 = 7'h1b == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_27; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_797 = 7'h1c == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_28; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_798 = 7'h1d == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_29; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_799 = 7'h1e == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_30; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_800 = 7'h1f == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_31; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_801 = 7'h20 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_32; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_802 = 7'h21 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_33; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_803 = 7'h22 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_34; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_804 = 7'h23 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_35; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_805 = 7'h24 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_36; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_806 = 7'h25 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_37; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_807 = 7'h26 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_38; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_808 = 7'h27 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_39; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_809 = 7'h28 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_40; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_810 = 7'h29 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_41; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_811 = 7'h2a == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_42; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_812 = 7'h2b == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_43; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_813 = 7'h2c == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_44; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_814 = 7'h2d == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_45; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_815 = 7'h2e == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_46; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_816 = 7'h2f == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_47; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_817 = 7'h30 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_48; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_818 = 7'h31 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_49; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_819 = 7'h32 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_50; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_820 = 7'h33 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_51; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_821 = 7'h34 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_52; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_822 = 7'h35 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_53; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_823 = 7'h36 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_54; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_824 = 7'h37 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_55; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_825 = 7'h38 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_56; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_826 = 7'h39 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_57; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_827 = 7'h3a == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_58; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_828 = 7'h3b == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_59; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_829 = 7'h3c == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_60; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_830 = 7'h3d == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_61; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_831 = 7'h3e == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_62; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_832 = 7'h3f == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_63; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_833 = 7'h40 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_64; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_834 = 7'h41 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_65; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_835 = 7'h42 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_66; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_836 = 7'h43 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_67; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_837 = 7'h44 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_68; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_838 = 7'h45 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_69; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_839 = 7'h46 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_70; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_840 = 7'h47 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_71; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_841 = 7'h48 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_72; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_842 = 7'h49 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_73; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_843 = 7'h4a == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_74; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_844 = 7'h4b == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_75; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_845 = 7'h4c == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_76; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_846 = 7'h4d == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_77; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_847 = 7'h4e == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_78; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_848 = 7'h4f == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_79; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_849 = 7'h50 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_80; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_850 = 7'h51 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_81; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_851 = 7'h52 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_82; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_852 = 7'h53 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_83; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_853 = 7'h54 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_84; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_854 = 7'h55 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_85; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_855 = 7'h56 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_86; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_856 = 7'h57 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_87; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_857 = 7'h58 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_88; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_858 = 7'h59 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_89; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_859 = 7'h5a == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_90; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_860 = 7'h5b == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_91; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_861 = 7'h5c == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_92; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_862 = 7'h5d == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_93; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_863 = 7'h5e == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_94; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_864 = 7'h5f == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_95; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_865 = 7'h60 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_96; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_866 = 7'h61 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_97; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_867 = 7'h62 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_98; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_868 = 7'h63 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_99; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_869 = 7'h64 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_100; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_870 = 7'h65 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_101; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_871 = 7'h66 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_102; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_872 = 7'h67 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_103; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_873 = 7'h68 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_104; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_874 = 7'h69 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_105; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_875 = 7'h6a == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_106; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_876 = 7'h6b == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_107; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_877 = 7'h6c == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_108; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_878 = 7'h6d == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_109; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_879 = 7'h6e == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_110; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_880 = 7'h6f == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_111; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_881 = 7'h70 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_112; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_882 = 7'h71 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_113; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_883 = 7'h72 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_114; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_884 = 7'h73 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_115; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_885 = 7'h74 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_116; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_886 = 7'h75 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_117; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_887 = 7'h76 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_118; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_888 = 7'h77 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_119; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_889 = 7'h78 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_120; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_890 = 7'h79 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_121; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_891 = 7'h7a == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_122; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_892 = 7'h7b == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_123; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_893 = 7'h7c == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_124; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_894 = 7'h7d == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_125; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_895 = 7'h7e == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_126; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_896 = 7'h7f == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_127; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [63:0] _rob_tscs_T_31 = {{32'd0}, tsc}; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_897 = 7'h0 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_0; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_898 = 7'h1 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_1; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_899 = 7'h2 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_2; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_900 = 7'h3 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_3; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_901 = 7'h4 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_4; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_902 = 7'h5 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_5; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_903 = 7'h6 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_6; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_904 = 7'h7 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_7; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_905 = 7'h8 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_8; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_906 = 7'h9 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_9; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_907 = 7'ha == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_10; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_908 = 7'hb == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_11; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_909 = 7'hc == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_12; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_910 = 7'hd == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_13; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_911 = 7'he == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_14; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_912 = 7'hf == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_15; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_913 = 7'h10 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_16; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_914 = 7'h11 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_17; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_915 = 7'h12 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_18; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_916 = 7'h13 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_19; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_917 = 7'h14 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_20; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_918 = 7'h15 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_21; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_919 = 7'h16 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_22; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_920 = 7'h17 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_23; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_921 = 7'h18 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_24; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_922 = 7'h19 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_25; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_923 = 7'h1a == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_26; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_924 = 7'h1b == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_27; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_925 = 7'h1c == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_28; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_926 = 7'h1d == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_29; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_927 = 7'h1e == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_30; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_928 = 7'h1f == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_31; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_929 = 7'h20 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_32; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_930 = 7'h21 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_33; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_931 = 7'h22 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_34; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_932 = 7'h23 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_35; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_933 = 7'h24 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_36; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_934 = 7'h25 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_37; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_935 = 7'h26 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_38; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_936 = 7'h27 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_39; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_937 = 7'h28 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_40; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_938 = 7'h29 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_41; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_939 = 7'h2a == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_42; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_940 = 7'h2b == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_43; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_941 = 7'h2c == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_44; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_942 = 7'h2d == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_45; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_943 = 7'h2e == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_46; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_944 = 7'h2f == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_47; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_945 = 7'h30 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_48; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_946 = 7'h31 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_49; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_947 = 7'h32 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_50; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_948 = 7'h33 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_51; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_949 = 7'h34 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_52; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_950 = 7'h35 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_53; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_951 = 7'h36 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_54; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_952 = 7'h37 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_55; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_953 = 7'h38 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_56; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_954 = 7'h39 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_57; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_955 = 7'h3a == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_58; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_956 = 7'h3b == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_59; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_957 = 7'h3c == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_60; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_958 = 7'h3d == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_61; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_959 = 7'h3e == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_62; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_960 = 7'h3f == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_63; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_961 = 7'h40 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_64; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_962 = 7'h41 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_65; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_963 = 7'h42 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_66; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_964 = 7'h43 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_67; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_965 = 7'h44 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_68; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_966 = 7'h45 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_69; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_967 = 7'h46 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_70; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_968 = 7'h47 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_71; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_969 = 7'h48 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_72; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_970 = 7'h49 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_73; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_971 = 7'h4a == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_74; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_972 = 7'h4b == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_75; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_973 = 7'h4c == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_76; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_974 = 7'h4d == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_77; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_975 = 7'h4e == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_78; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_976 = 7'h4f == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_79; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_977 = 7'h50 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_80; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_978 = 7'h51 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_81; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_979 = 7'h52 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_82; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_980 = 7'h53 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_83; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_981 = 7'h54 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_84; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_982 = 7'h55 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_85; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_983 = 7'h56 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_86; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_984 = 7'h57 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_87; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_985 = 7'h58 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_88; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_986 = 7'h59 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_89; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_987 = 7'h5a == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_90; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_988 = 7'h5b == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_91; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_989 = 7'h5c == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_92; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_990 = 7'h5d == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_93; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_991 = 7'h5e == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_94; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_992 = 7'h5f == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_95; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_993 = 7'h60 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_96; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_994 = 7'h61 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_97; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_995 = 7'h62 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_98; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_996 = 7'h63 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_99; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_997 = 7'h64 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_100; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_998 = 7'h65 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_101; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_999 = 7'h66 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_102; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1000 = 7'h67 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_103; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1001 = 7'h68 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_104; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1002 = 7'h69 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_105; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1003 = 7'h6a == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_106; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1004 = 7'h6b == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_107; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1005 = 7'h6c == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_108; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1006 = 7'h6d == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_109; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1007 = 7'h6e == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_110; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1008 = 7'h6f == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_111; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1009 = 7'h70 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_112; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1010 = 7'h71 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_113; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1011 = 7'h72 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_114; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1012 = 7'h73 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_115; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1013 = 7'h74 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_116; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1014 = 7'h75 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_117; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1015 = 7'h76 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_118; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1016 = 7'h77 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_119; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1017 = 7'h78 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_120; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1018 = 7'h79 == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_121; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1019 = 7'h7a == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_122; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1020 = 7'h7b == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_123; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1021 = 7'h7c == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_124; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1022 = 7'h7d == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_125; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1023 = 7'h7e == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_126; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1024 = 7'h7f == rob_alloc_ids_0 ? _rob_tscs_T_31 : rob_tscs_127; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [31:0] _GEN_1025 = igen_io_fire ? _GEN_1 : rob_payload_0_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1026 = igen_io_fire ? _GEN_2 : rob_payload_1_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1027 = igen_io_fire ? _GEN_3 : rob_payload_2_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1028 = igen_io_fire ? _GEN_4 : rob_payload_3_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1029 = igen_io_fire ? _GEN_5 : rob_payload_4_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1030 = igen_io_fire ? _GEN_6 : rob_payload_5_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1031 = igen_io_fire ? _GEN_7 : rob_payload_6_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1032 = igen_io_fire ? _GEN_8 : rob_payload_7_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1033 = igen_io_fire ? _GEN_9 : rob_payload_8_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1034 = igen_io_fire ? _GEN_10 : rob_payload_9_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1035 = igen_io_fire ? _GEN_11 : rob_payload_10_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1036 = igen_io_fire ? _GEN_12 : rob_payload_11_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1037 = igen_io_fire ? _GEN_13 : rob_payload_12_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1038 = igen_io_fire ? _GEN_14 : rob_payload_13_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1039 = igen_io_fire ? _GEN_15 : rob_payload_14_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1040 = igen_io_fire ? _GEN_16 : rob_payload_15_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1041 = igen_io_fire ? _GEN_17 : rob_payload_16_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1042 = igen_io_fire ? _GEN_18 : rob_payload_17_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1043 = igen_io_fire ? _GEN_19 : rob_payload_18_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1044 = igen_io_fire ? _GEN_20 : rob_payload_19_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1045 = igen_io_fire ? _GEN_21 : rob_payload_20_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1046 = igen_io_fire ? _GEN_22 : rob_payload_21_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1047 = igen_io_fire ? _GEN_23 : rob_payload_22_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1048 = igen_io_fire ? _GEN_24 : rob_payload_23_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1049 = igen_io_fire ? _GEN_25 : rob_payload_24_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1050 = igen_io_fire ? _GEN_26 : rob_payload_25_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1051 = igen_io_fire ? _GEN_27 : rob_payload_26_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1052 = igen_io_fire ? _GEN_28 : rob_payload_27_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1053 = igen_io_fire ? _GEN_29 : rob_payload_28_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1054 = igen_io_fire ? _GEN_30 : rob_payload_29_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1055 = igen_io_fire ? _GEN_31 : rob_payload_30_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1056 = igen_io_fire ? _GEN_32 : rob_payload_31_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1057 = igen_io_fire ? _GEN_33 : rob_payload_32_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1058 = igen_io_fire ? _GEN_34 : rob_payload_33_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1059 = igen_io_fire ? _GEN_35 : rob_payload_34_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1060 = igen_io_fire ? _GEN_36 : rob_payload_35_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1061 = igen_io_fire ? _GEN_37 : rob_payload_36_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1062 = igen_io_fire ? _GEN_38 : rob_payload_37_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1063 = igen_io_fire ? _GEN_39 : rob_payload_38_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1064 = igen_io_fire ? _GEN_40 : rob_payload_39_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1065 = igen_io_fire ? _GEN_41 : rob_payload_40_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1066 = igen_io_fire ? _GEN_42 : rob_payload_41_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1067 = igen_io_fire ? _GEN_43 : rob_payload_42_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1068 = igen_io_fire ? _GEN_44 : rob_payload_43_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1069 = igen_io_fire ? _GEN_45 : rob_payload_44_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1070 = igen_io_fire ? _GEN_46 : rob_payload_45_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1071 = igen_io_fire ? _GEN_47 : rob_payload_46_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1072 = igen_io_fire ? _GEN_48 : rob_payload_47_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1073 = igen_io_fire ? _GEN_49 : rob_payload_48_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1074 = igen_io_fire ? _GEN_50 : rob_payload_49_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1075 = igen_io_fire ? _GEN_51 : rob_payload_50_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1076 = igen_io_fire ? _GEN_52 : rob_payload_51_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1077 = igen_io_fire ? _GEN_53 : rob_payload_52_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1078 = igen_io_fire ? _GEN_54 : rob_payload_53_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1079 = igen_io_fire ? _GEN_55 : rob_payload_54_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1080 = igen_io_fire ? _GEN_56 : rob_payload_55_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1081 = igen_io_fire ? _GEN_57 : rob_payload_56_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1082 = igen_io_fire ? _GEN_58 : rob_payload_57_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1083 = igen_io_fire ? _GEN_59 : rob_payload_58_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1084 = igen_io_fire ? _GEN_60 : rob_payload_59_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1085 = igen_io_fire ? _GEN_61 : rob_payload_60_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1086 = igen_io_fire ? _GEN_62 : rob_payload_61_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1087 = igen_io_fire ? _GEN_63 : rob_payload_62_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1088 = igen_io_fire ? _GEN_64 : rob_payload_63_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1089 = igen_io_fire ? _GEN_65 : rob_payload_64_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1090 = igen_io_fire ? _GEN_66 : rob_payload_65_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1091 = igen_io_fire ? _GEN_67 : rob_payload_66_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1092 = igen_io_fire ? _GEN_68 : rob_payload_67_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1093 = igen_io_fire ? _GEN_69 : rob_payload_68_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1094 = igen_io_fire ? _GEN_70 : rob_payload_69_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1095 = igen_io_fire ? _GEN_71 : rob_payload_70_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1096 = igen_io_fire ? _GEN_72 : rob_payload_71_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1097 = igen_io_fire ? _GEN_73 : rob_payload_72_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1098 = igen_io_fire ? _GEN_74 : rob_payload_73_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1099 = igen_io_fire ? _GEN_75 : rob_payload_74_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1100 = igen_io_fire ? _GEN_76 : rob_payload_75_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1101 = igen_io_fire ? _GEN_77 : rob_payload_76_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1102 = igen_io_fire ? _GEN_78 : rob_payload_77_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1103 = igen_io_fire ? _GEN_79 : rob_payload_78_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1104 = igen_io_fire ? _GEN_80 : rob_payload_79_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1105 = igen_io_fire ? _GEN_81 : rob_payload_80_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1106 = igen_io_fire ? _GEN_82 : rob_payload_81_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1107 = igen_io_fire ? _GEN_83 : rob_payload_82_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1108 = igen_io_fire ? _GEN_84 : rob_payload_83_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1109 = igen_io_fire ? _GEN_85 : rob_payload_84_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1110 = igen_io_fire ? _GEN_86 : rob_payload_85_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1111 = igen_io_fire ? _GEN_87 : rob_payload_86_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1112 = igen_io_fire ? _GEN_88 : rob_payload_87_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1113 = igen_io_fire ? _GEN_89 : rob_payload_88_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1114 = igen_io_fire ? _GEN_90 : rob_payload_89_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1115 = igen_io_fire ? _GEN_91 : rob_payload_90_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1116 = igen_io_fire ? _GEN_92 : rob_payload_91_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1117 = igen_io_fire ? _GEN_93 : rob_payload_92_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1118 = igen_io_fire ? _GEN_94 : rob_payload_93_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1119 = igen_io_fire ? _GEN_95 : rob_payload_94_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1120 = igen_io_fire ? _GEN_96 : rob_payload_95_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1121 = igen_io_fire ? _GEN_97 : rob_payload_96_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1122 = igen_io_fire ? _GEN_98 : rob_payload_97_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1123 = igen_io_fire ? _GEN_99 : rob_payload_98_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1124 = igen_io_fire ? _GEN_100 : rob_payload_99_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1125 = igen_io_fire ? _GEN_101 : rob_payload_100_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1126 = igen_io_fire ? _GEN_102 : rob_payload_101_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1127 = igen_io_fire ? _GEN_103 : rob_payload_102_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1128 = igen_io_fire ? _GEN_104 : rob_payload_103_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1129 = igen_io_fire ? _GEN_105 : rob_payload_104_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1130 = igen_io_fire ? _GEN_106 : rob_payload_105_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1131 = igen_io_fire ? _GEN_107 : rob_payload_106_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1132 = igen_io_fire ? _GEN_108 : rob_payload_107_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1133 = igen_io_fire ? _GEN_109 : rob_payload_108_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1134 = igen_io_fire ? _GEN_110 : rob_payload_109_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1135 = igen_io_fire ? _GEN_111 : rob_payload_110_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1136 = igen_io_fire ? _GEN_112 : rob_payload_111_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1137 = igen_io_fire ? _GEN_113 : rob_payload_112_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1138 = igen_io_fire ? _GEN_114 : rob_payload_113_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1139 = igen_io_fire ? _GEN_115 : rob_payload_114_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1140 = igen_io_fire ? _GEN_116 : rob_payload_115_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1141 = igen_io_fire ? _GEN_117 : rob_payload_116_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1142 = igen_io_fire ? _GEN_118 : rob_payload_117_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1143 = igen_io_fire ? _GEN_119 : rob_payload_118_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1144 = igen_io_fire ? _GEN_120 : rob_payload_119_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1145 = igen_io_fire ? _GEN_121 : rob_payload_120_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1146 = igen_io_fire ? _GEN_122 : rob_payload_121_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1147 = igen_io_fire ? _GEN_123 : rob_payload_122_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1148 = igen_io_fire ? _GEN_124 : rob_payload_123_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1149 = igen_io_fire ? _GEN_125 : rob_payload_124_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1150 = igen_io_fire ? _GEN_126 : rob_payload_125_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1151 = igen_io_fire ? _GEN_127 : rob_payload_126_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1152 = igen_io_fire ? _GEN_128 : rob_payload_127_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1153 = igen_io_fire ? _GEN_129 : rob_payload_0_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1154 = igen_io_fire ? _GEN_130 : rob_payload_1_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1155 = igen_io_fire ? _GEN_131 : rob_payload_2_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1156 = igen_io_fire ? _GEN_132 : rob_payload_3_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1157 = igen_io_fire ? _GEN_133 : rob_payload_4_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1158 = igen_io_fire ? _GEN_134 : rob_payload_5_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1159 = igen_io_fire ? _GEN_135 : rob_payload_6_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1160 = igen_io_fire ? _GEN_136 : rob_payload_7_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1161 = igen_io_fire ? _GEN_137 : rob_payload_8_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1162 = igen_io_fire ? _GEN_138 : rob_payload_9_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1163 = igen_io_fire ? _GEN_139 : rob_payload_10_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1164 = igen_io_fire ? _GEN_140 : rob_payload_11_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1165 = igen_io_fire ? _GEN_141 : rob_payload_12_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1166 = igen_io_fire ? _GEN_142 : rob_payload_13_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1167 = igen_io_fire ? _GEN_143 : rob_payload_14_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1168 = igen_io_fire ? _GEN_144 : rob_payload_15_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1169 = igen_io_fire ? _GEN_145 : rob_payload_16_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1170 = igen_io_fire ? _GEN_146 : rob_payload_17_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1171 = igen_io_fire ? _GEN_147 : rob_payload_18_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1172 = igen_io_fire ? _GEN_148 : rob_payload_19_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1173 = igen_io_fire ? _GEN_149 : rob_payload_20_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1174 = igen_io_fire ? _GEN_150 : rob_payload_21_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1175 = igen_io_fire ? _GEN_151 : rob_payload_22_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1176 = igen_io_fire ? _GEN_152 : rob_payload_23_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1177 = igen_io_fire ? _GEN_153 : rob_payload_24_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1178 = igen_io_fire ? _GEN_154 : rob_payload_25_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1179 = igen_io_fire ? _GEN_155 : rob_payload_26_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1180 = igen_io_fire ? _GEN_156 : rob_payload_27_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1181 = igen_io_fire ? _GEN_157 : rob_payload_28_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1182 = igen_io_fire ? _GEN_158 : rob_payload_29_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1183 = igen_io_fire ? _GEN_159 : rob_payload_30_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1184 = igen_io_fire ? _GEN_160 : rob_payload_31_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1185 = igen_io_fire ? _GEN_161 : rob_payload_32_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1186 = igen_io_fire ? _GEN_162 : rob_payload_33_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1187 = igen_io_fire ? _GEN_163 : rob_payload_34_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1188 = igen_io_fire ? _GEN_164 : rob_payload_35_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1189 = igen_io_fire ? _GEN_165 : rob_payload_36_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1190 = igen_io_fire ? _GEN_166 : rob_payload_37_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1191 = igen_io_fire ? _GEN_167 : rob_payload_38_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1192 = igen_io_fire ? _GEN_168 : rob_payload_39_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1193 = igen_io_fire ? _GEN_169 : rob_payload_40_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1194 = igen_io_fire ? _GEN_170 : rob_payload_41_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1195 = igen_io_fire ? _GEN_171 : rob_payload_42_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1196 = igen_io_fire ? _GEN_172 : rob_payload_43_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1197 = igen_io_fire ? _GEN_173 : rob_payload_44_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1198 = igen_io_fire ? _GEN_174 : rob_payload_45_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1199 = igen_io_fire ? _GEN_175 : rob_payload_46_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1200 = igen_io_fire ? _GEN_176 : rob_payload_47_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1201 = igen_io_fire ? _GEN_177 : rob_payload_48_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1202 = igen_io_fire ? _GEN_178 : rob_payload_49_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1203 = igen_io_fire ? _GEN_179 : rob_payload_50_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1204 = igen_io_fire ? _GEN_180 : rob_payload_51_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1205 = igen_io_fire ? _GEN_181 : rob_payload_52_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1206 = igen_io_fire ? _GEN_182 : rob_payload_53_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1207 = igen_io_fire ? _GEN_183 : rob_payload_54_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1208 = igen_io_fire ? _GEN_184 : rob_payload_55_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1209 = igen_io_fire ? _GEN_185 : rob_payload_56_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1210 = igen_io_fire ? _GEN_186 : rob_payload_57_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1211 = igen_io_fire ? _GEN_187 : rob_payload_58_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1212 = igen_io_fire ? _GEN_188 : rob_payload_59_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1213 = igen_io_fire ? _GEN_189 : rob_payload_60_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1214 = igen_io_fire ? _GEN_190 : rob_payload_61_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1215 = igen_io_fire ? _GEN_191 : rob_payload_62_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1216 = igen_io_fire ? _GEN_192 : rob_payload_63_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1217 = igen_io_fire ? _GEN_193 : rob_payload_64_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1218 = igen_io_fire ? _GEN_194 : rob_payload_65_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1219 = igen_io_fire ? _GEN_195 : rob_payload_66_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1220 = igen_io_fire ? _GEN_196 : rob_payload_67_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1221 = igen_io_fire ? _GEN_197 : rob_payload_68_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1222 = igen_io_fire ? _GEN_198 : rob_payload_69_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1223 = igen_io_fire ? _GEN_199 : rob_payload_70_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1224 = igen_io_fire ? _GEN_200 : rob_payload_71_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1225 = igen_io_fire ? _GEN_201 : rob_payload_72_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1226 = igen_io_fire ? _GEN_202 : rob_payload_73_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1227 = igen_io_fire ? _GEN_203 : rob_payload_74_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1228 = igen_io_fire ? _GEN_204 : rob_payload_75_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1229 = igen_io_fire ? _GEN_205 : rob_payload_76_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1230 = igen_io_fire ? _GEN_206 : rob_payload_77_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1231 = igen_io_fire ? _GEN_207 : rob_payload_78_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1232 = igen_io_fire ? _GEN_208 : rob_payload_79_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1233 = igen_io_fire ? _GEN_209 : rob_payload_80_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1234 = igen_io_fire ? _GEN_210 : rob_payload_81_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1235 = igen_io_fire ? _GEN_211 : rob_payload_82_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1236 = igen_io_fire ? _GEN_212 : rob_payload_83_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1237 = igen_io_fire ? _GEN_213 : rob_payload_84_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1238 = igen_io_fire ? _GEN_214 : rob_payload_85_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1239 = igen_io_fire ? _GEN_215 : rob_payload_86_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1240 = igen_io_fire ? _GEN_216 : rob_payload_87_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1241 = igen_io_fire ? _GEN_217 : rob_payload_88_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1242 = igen_io_fire ? _GEN_218 : rob_payload_89_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1243 = igen_io_fire ? _GEN_219 : rob_payload_90_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1244 = igen_io_fire ? _GEN_220 : rob_payload_91_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1245 = igen_io_fire ? _GEN_221 : rob_payload_92_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1246 = igen_io_fire ? _GEN_222 : rob_payload_93_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1247 = igen_io_fire ? _GEN_223 : rob_payload_94_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1248 = igen_io_fire ? _GEN_224 : rob_payload_95_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1249 = igen_io_fire ? _GEN_225 : rob_payload_96_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1250 = igen_io_fire ? _GEN_226 : rob_payload_97_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1251 = igen_io_fire ? _GEN_227 : rob_payload_98_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1252 = igen_io_fire ? _GEN_228 : rob_payload_99_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1253 = igen_io_fire ? _GEN_229 : rob_payload_100_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1254 = igen_io_fire ? _GEN_230 : rob_payload_101_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1255 = igen_io_fire ? _GEN_231 : rob_payload_102_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1256 = igen_io_fire ? _GEN_232 : rob_payload_103_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1257 = igen_io_fire ? _GEN_233 : rob_payload_104_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1258 = igen_io_fire ? _GEN_234 : rob_payload_105_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1259 = igen_io_fire ? _GEN_235 : rob_payload_106_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1260 = igen_io_fire ? _GEN_236 : rob_payload_107_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1261 = igen_io_fire ? _GEN_237 : rob_payload_108_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1262 = igen_io_fire ? _GEN_238 : rob_payload_109_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1263 = igen_io_fire ? _GEN_239 : rob_payload_110_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1264 = igen_io_fire ? _GEN_240 : rob_payload_111_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1265 = igen_io_fire ? _GEN_241 : rob_payload_112_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1266 = igen_io_fire ? _GEN_242 : rob_payload_113_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1267 = igen_io_fire ? _GEN_243 : rob_payload_114_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1268 = igen_io_fire ? _GEN_244 : rob_payload_115_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1269 = igen_io_fire ? _GEN_245 : rob_payload_116_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1270 = igen_io_fire ? _GEN_246 : rob_payload_117_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1271 = igen_io_fire ? _GEN_247 : rob_payload_118_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1272 = igen_io_fire ? _GEN_248 : rob_payload_119_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1273 = igen_io_fire ? _GEN_249 : rob_payload_120_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1274 = igen_io_fire ? _GEN_250 : rob_payload_121_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1275 = igen_io_fire ? _GEN_251 : rob_payload_122_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1276 = igen_io_fire ? _GEN_252 : rob_payload_123_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1277 = igen_io_fire ? _GEN_253 : rob_payload_124_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1278 = igen_io_fire ? _GEN_254 : rob_payload_125_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1279 = igen_io_fire ? _GEN_255 : rob_payload_126_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1280 = igen_io_fire ? _GEN_256 : rob_payload_127_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1281 = igen_io_fire ? _GEN_257 : rob_payload_0_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1282 = igen_io_fire ? _GEN_258 : rob_payload_1_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1283 = igen_io_fire ? _GEN_259 : rob_payload_2_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1284 = igen_io_fire ? _GEN_260 : rob_payload_3_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1285 = igen_io_fire ? _GEN_261 : rob_payload_4_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1286 = igen_io_fire ? _GEN_262 : rob_payload_5_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1287 = igen_io_fire ? _GEN_263 : rob_payload_6_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1288 = igen_io_fire ? _GEN_264 : rob_payload_7_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1289 = igen_io_fire ? _GEN_265 : rob_payload_8_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1290 = igen_io_fire ? _GEN_266 : rob_payload_9_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1291 = igen_io_fire ? _GEN_267 : rob_payload_10_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1292 = igen_io_fire ? _GEN_268 : rob_payload_11_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1293 = igen_io_fire ? _GEN_269 : rob_payload_12_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1294 = igen_io_fire ? _GEN_270 : rob_payload_13_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1295 = igen_io_fire ? _GEN_271 : rob_payload_14_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1296 = igen_io_fire ? _GEN_272 : rob_payload_15_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1297 = igen_io_fire ? _GEN_273 : rob_payload_16_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1298 = igen_io_fire ? _GEN_274 : rob_payload_17_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1299 = igen_io_fire ? _GEN_275 : rob_payload_18_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1300 = igen_io_fire ? _GEN_276 : rob_payload_19_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1301 = igen_io_fire ? _GEN_277 : rob_payload_20_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1302 = igen_io_fire ? _GEN_278 : rob_payload_21_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1303 = igen_io_fire ? _GEN_279 : rob_payload_22_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1304 = igen_io_fire ? _GEN_280 : rob_payload_23_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1305 = igen_io_fire ? _GEN_281 : rob_payload_24_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1306 = igen_io_fire ? _GEN_282 : rob_payload_25_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1307 = igen_io_fire ? _GEN_283 : rob_payload_26_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1308 = igen_io_fire ? _GEN_284 : rob_payload_27_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1309 = igen_io_fire ? _GEN_285 : rob_payload_28_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1310 = igen_io_fire ? _GEN_286 : rob_payload_29_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1311 = igen_io_fire ? _GEN_287 : rob_payload_30_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1312 = igen_io_fire ? _GEN_288 : rob_payload_31_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1313 = igen_io_fire ? _GEN_289 : rob_payload_32_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1314 = igen_io_fire ? _GEN_290 : rob_payload_33_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1315 = igen_io_fire ? _GEN_291 : rob_payload_34_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1316 = igen_io_fire ? _GEN_292 : rob_payload_35_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1317 = igen_io_fire ? _GEN_293 : rob_payload_36_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1318 = igen_io_fire ? _GEN_294 : rob_payload_37_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1319 = igen_io_fire ? _GEN_295 : rob_payload_38_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1320 = igen_io_fire ? _GEN_296 : rob_payload_39_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1321 = igen_io_fire ? _GEN_297 : rob_payload_40_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1322 = igen_io_fire ? _GEN_298 : rob_payload_41_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1323 = igen_io_fire ? _GEN_299 : rob_payload_42_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1324 = igen_io_fire ? _GEN_300 : rob_payload_43_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1325 = igen_io_fire ? _GEN_301 : rob_payload_44_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1326 = igen_io_fire ? _GEN_302 : rob_payload_45_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1327 = igen_io_fire ? _GEN_303 : rob_payload_46_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1328 = igen_io_fire ? _GEN_304 : rob_payload_47_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1329 = igen_io_fire ? _GEN_305 : rob_payload_48_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1330 = igen_io_fire ? _GEN_306 : rob_payload_49_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1331 = igen_io_fire ? _GEN_307 : rob_payload_50_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1332 = igen_io_fire ? _GEN_308 : rob_payload_51_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1333 = igen_io_fire ? _GEN_309 : rob_payload_52_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1334 = igen_io_fire ? _GEN_310 : rob_payload_53_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1335 = igen_io_fire ? _GEN_311 : rob_payload_54_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1336 = igen_io_fire ? _GEN_312 : rob_payload_55_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1337 = igen_io_fire ? _GEN_313 : rob_payload_56_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1338 = igen_io_fire ? _GEN_314 : rob_payload_57_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1339 = igen_io_fire ? _GEN_315 : rob_payload_58_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1340 = igen_io_fire ? _GEN_316 : rob_payload_59_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1341 = igen_io_fire ? _GEN_317 : rob_payload_60_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1342 = igen_io_fire ? _GEN_318 : rob_payload_61_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1343 = igen_io_fire ? _GEN_319 : rob_payload_62_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1344 = igen_io_fire ? _GEN_320 : rob_payload_63_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1345 = igen_io_fire ? _GEN_321 : rob_payload_64_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1346 = igen_io_fire ? _GEN_322 : rob_payload_65_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1347 = igen_io_fire ? _GEN_323 : rob_payload_66_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1348 = igen_io_fire ? _GEN_324 : rob_payload_67_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1349 = igen_io_fire ? _GEN_325 : rob_payload_68_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1350 = igen_io_fire ? _GEN_326 : rob_payload_69_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1351 = igen_io_fire ? _GEN_327 : rob_payload_70_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1352 = igen_io_fire ? _GEN_328 : rob_payload_71_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1353 = igen_io_fire ? _GEN_329 : rob_payload_72_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1354 = igen_io_fire ? _GEN_330 : rob_payload_73_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1355 = igen_io_fire ? _GEN_331 : rob_payload_74_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1356 = igen_io_fire ? _GEN_332 : rob_payload_75_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1357 = igen_io_fire ? _GEN_333 : rob_payload_76_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1358 = igen_io_fire ? _GEN_334 : rob_payload_77_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1359 = igen_io_fire ? _GEN_335 : rob_payload_78_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1360 = igen_io_fire ? _GEN_336 : rob_payload_79_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1361 = igen_io_fire ? _GEN_337 : rob_payload_80_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1362 = igen_io_fire ? _GEN_338 : rob_payload_81_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1363 = igen_io_fire ? _GEN_339 : rob_payload_82_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1364 = igen_io_fire ? _GEN_340 : rob_payload_83_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1365 = igen_io_fire ? _GEN_341 : rob_payload_84_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1366 = igen_io_fire ? _GEN_342 : rob_payload_85_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1367 = igen_io_fire ? _GEN_343 : rob_payload_86_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1368 = igen_io_fire ? _GEN_344 : rob_payload_87_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1369 = igen_io_fire ? _GEN_345 : rob_payload_88_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1370 = igen_io_fire ? _GEN_346 : rob_payload_89_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1371 = igen_io_fire ? _GEN_347 : rob_payload_90_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1372 = igen_io_fire ? _GEN_348 : rob_payload_91_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1373 = igen_io_fire ? _GEN_349 : rob_payload_92_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1374 = igen_io_fire ? _GEN_350 : rob_payload_93_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1375 = igen_io_fire ? _GEN_351 : rob_payload_94_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1376 = igen_io_fire ? _GEN_352 : rob_payload_95_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1377 = igen_io_fire ? _GEN_353 : rob_payload_96_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1378 = igen_io_fire ? _GEN_354 : rob_payload_97_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1379 = igen_io_fire ? _GEN_355 : rob_payload_98_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1380 = igen_io_fire ? _GEN_356 : rob_payload_99_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1381 = igen_io_fire ? _GEN_357 : rob_payload_100_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1382 = igen_io_fire ? _GEN_358 : rob_payload_101_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1383 = igen_io_fire ? _GEN_359 : rob_payload_102_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1384 = igen_io_fire ? _GEN_360 : rob_payload_103_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1385 = igen_io_fire ? _GEN_361 : rob_payload_104_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1386 = igen_io_fire ? _GEN_362 : rob_payload_105_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1387 = igen_io_fire ? _GEN_363 : rob_payload_106_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1388 = igen_io_fire ? _GEN_364 : rob_payload_107_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1389 = igen_io_fire ? _GEN_365 : rob_payload_108_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1390 = igen_io_fire ? _GEN_366 : rob_payload_109_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1391 = igen_io_fire ? _GEN_367 : rob_payload_110_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1392 = igen_io_fire ? _GEN_368 : rob_payload_111_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1393 = igen_io_fire ? _GEN_369 : rob_payload_112_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1394 = igen_io_fire ? _GEN_370 : rob_payload_113_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1395 = igen_io_fire ? _GEN_371 : rob_payload_114_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1396 = igen_io_fire ? _GEN_372 : rob_payload_115_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1397 = igen_io_fire ? _GEN_373 : rob_payload_116_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1398 = igen_io_fire ? _GEN_374 : rob_payload_117_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1399 = igen_io_fire ? _GEN_375 : rob_payload_118_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1400 = igen_io_fire ? _GEN_376 : rob_payload_119_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1401 = igen_io_fire ? _GEN_377 : rob_payload_120_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1402 = igen_io_fire ? _GEN_378 : rob_payload_121_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1403 = igen_io_fire ? _GEN_379 : rob_payload_122_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1404 = igen_io_fire ? _GEN_380 : rob_payload_123_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1405 = igen_io_fire ? _GEN_381 : rob_payload_124_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1406 = igen_io_fire ? _GEN_382 : rob_payload_125_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1407 = igen_io_fire ? _GEN_383 : rob_payload_126_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1408 = igen_io_fire ? _GEN_384 : rob_payload_127_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [1:0] _GEN_1409 = igen_io_fire ? _GEN_385 : rob_egress_id_0; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1410 = igen_io_fire ? _GEN_386 : rob_egress_id_1; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1411 = igen_io_fire ? _GEN_387 : rob_egress_id_2; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1412 = igen_io_fire ? _GEN_388 : rob_egress_id_3; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1413 = igen_io_fire ? _GEN_389 : rob_egress_id_4; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1414 = igen_io_fire ? _GEN_390 : rob_egress_id_5; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1415 = igen_io_fire ? _GEN_391 : rob_egress_id_6; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1416 = igen_io_fire ? _GEN_392 : rob_egress_id_7; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1417 = igen_io_fire ? _GEN_393 : rob_egress_id_8; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1418 = igen_io_fire ? _GEN_394 : rob_egress_id_9; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1419 = igen_io_fire ? _GEN_395 : rob_egress_id_10; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1420 = igen_io_fire ? _GEN_396 : rob_egress_id_11; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1421 = igen_io_fire ? _GEN_397 : rob_egress_id_12; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1422 = igen_io_fire ? _GEN_398 : rob_egress_id_13; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1423 = igen_io_fire ? _GEN_399 : rob_egress_id_14; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1424 = igen_io_fire ? _GEN_400 : rob_egress_id_15; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1425 = igen_io_fire ? _GEN_401 : rob_egress_id_16; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1426 = igen_io_fire ? _GEN_402 : rob_egress_id_17; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1427 = igen_io_fire ? _GEN_403 : rob_egress_id_18; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1428 = igen_io_fire ? _GEN_404 : rob_egress_id_19; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1429 = igen_io_fire ? _GEN_405 : rob_egress_id_20; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1430 = igen_io_fire ? _GEN_406 : rob_egress_id_21; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1431 = igen_io_fire ? _GEN_407 : rob_egress_id_22; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1432 = igen_io_fire ? _GEN_408 : rob_egress_id_23; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1433 = igen_io_fire ? _GEN_409 : rob_egress_id_24; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1434 = igen_io_fire ? _GEN_410 : rob_egress_id_25; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1435 = igen_io_fire ? _GEN_411 : rob_egress_id_26; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1436 = igen_io_fire ? _GEN_412 : rob_egress_id_27; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1437 = igen_io_fire ? _GEN_413 : rob_egress_id_28; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1438 = igen_io_fire ? _GEN_414 : rob_egress_id_29; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1439 = igen_io_fire ? _GEN_415 : rob_egress_id_30; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1440 = igen_io_fire ? _GEN_416 : rob_egress_id_31; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1441 = igen_io_fire ? _GEN_417 : rob_egress_id_32; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1442 = igen_io_fire ? _GEN_418 : rob_egress_id_33; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1443 = igen_io_fire ? _GEN_419 : rob_egress_id_34; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1444 = igen_io_fire ? _GEN_420 : rob_egress_id_35; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1445 = igen_io_fire ? _GEN_421 : rob_egress_id_36; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1446 = igen_io_fire ? _GEN_422 : rob_egress_id_37; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1447 = igen_io_fire ? _GEN_423 : rob_egress_id_38; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1448 = igen_io_fire ? _GEN_424 : rob_egress_id_39; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1449 = igen_io_fire ? _GEN_425 : rob_egress_id_40; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1450 = igen_io_fire ? _GEN_426 : rob_egress_id_41; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1451 = igen_io_fire ? _GEN_427 : rob_egress_id_42; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1452 = igen_io_fire ? _GEN_428 : rob_egress_id_43; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1453 = igen_io_fire ? _GEN_429 : rob_egress_id_44; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1454 = igen_io_fire ? _GEN_430 : rob_egress_id_45; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1455 = igen_io_fire ? _GEN_431 : rob_egress_id_46; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1456 = igen_io_fire ? _GEN_432 : rob_egress_id_47; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1457 = igen_io_fire ? _GEN_433 : rob_egress_id_48; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1458 = igen_io_fire ? _GEN_434 : rob_egress_id_49; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1459 = igen_io_fire ? _GEN_435 : rob_egress_id_50; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1460 = igen_io_fire ? _GEN_436 : rob_egress_id_51; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1461 = igen_io_fire ? _GEN_437 : rob_egress_id_52; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1462 = igen_io_fire ? _GEN_438 : rob_egress_id_53; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1463 = igen_io_fire ? _GEN_439 : rob_egress_id_54; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1464 = igen_io_fire ? _GEN_440 : rob_egress_id_55; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1465 = igen_io_fire ? _GEN_441 : rob_egress_id_56; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1466 = igen_io_fire ? _GEN_442 : rob_egress_id_57; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1467 = igen_io_fire ? _GEN_443 : rob_egress_id_58; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1468 = igen_io_fire ? _GEN_444 : rob_egress_id_59; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1469 = igen_io_fire ? _GEN_445 : rob_egress_id_60; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1470 = igen_io_fire ? _GEN_446 : rob_egress_id_61; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1471 = igen_io_fire ? _GEN_447 : rob_egress_id_62; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1472 = igen_io_fire ? _GEN_448 : rob_egress_id_63; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1473 = igen_io_fire ? _GEN_449 : rob_egress_id_64; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1474 = igen_io_fire ? _GEN_450 : rob_egress_id_65; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1475 = igen_io_fire ? _GEN_451 : rob_egress_id_66; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1476 = igen_io_fire ? _GEN_452 : rob_egress_id_67; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1477 = igen_io_fire ? _GEN_453 : rob_egress_id_68; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1478 = igen_io_fire ? _GEN_454 : rob_egress_id_69; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1479 = igen_io_fire ? _GEN_455 : rob_egress_id_70; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1480 = igen_io_fire ? _GEN_456 : rob_egress_id_71; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1481 = igen_io_fire ? _GEN_457 : rob_egress_id_72; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1482 = igen_io_fire ? _GEN_458 : rob_egress_id_73; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1483 = igen_io_fire ? _GEN_459 : rob_egress_id_74; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1484 = igen_io_fire ? _GEN_460 : rob_egress_id_75; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1485 = igen_io_fire ? _GEN_461 : rob_egress_id_76; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1486 = igen_io_fire ? _GEN_462 : rob_egress_id_77; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1487 = igen_io_fire ? _GEN_463 : rob_egress_id_78; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1488 = igen_io_fire ? _GEN_464 : rob_egress_id_79; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1489 = igen_io_fire ? _GEN_465 : rob_egress_id_80; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1490 = igen_io_fire ? _GEN_466 : rob_egress_id_81; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1491 = igen_io_fire ? _GEN_467 : rob_egress_id_82; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1492 = igen_io_fire ? _GEN_468 : rob_egress_id_83; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1493 = igen_io_fire ? _GEN_469 : rob_egress_id_84; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1494 = igen_io_fire ? _GEN_470 : rob_egress_id_85; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1495 = igen_io_fire ? _GEN_471 : rob_egress_id_86; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1496 = igen_io_fire ? _GEN_472 : rob_egress_id_87; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1497 = igen_io_fire ? _GEN_473 : rob_egress_id_88; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1498 = igen_io_fire ? _GEN_474 : rob_egress_id_89; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1499 = igen_io_fire ? _GEN_475 : rob_egress_id_90; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1500 = igen_io_fire ? _GEN_476 : rob_egress_id_91; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1501 = igen_io_fire ? _GEN_477 : rob_egress_id_92; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1502 = igen_io_fire ? _GEN_478 : rob_egress_id_93; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1503 = igen_io_fire ? _GEN_479 : rob_egress_id_94; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1504 = igen_io_fire ? _GEN_480 : rob_egress_id_95; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1505 = igen_io_fire ? _GEN_481 : rob_egress_id_96; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1506 = igen_io_fire ? _GEN_482 : rob_egress_id_97; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1507 = igen_io_fire ? _GEN_483 : rob_egress_id_98; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1508 = igen_io_fire ? _GEN_484 : rob_egress_id_99; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1509 = igen_io_fire ? _GEN_485 : rob_egress_id_100; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1510 = igen_io_fire ? _GEN_486 : rob_egress_id_101; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1511 = igen_io_fire ? _GEN_487 : rob_egress_id_102; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1512 = igen_io_fire ? _GEN_488 : rob_egress_id_103; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1513 = igen_io_fire ? _GEN_489 : rob_egress_id_104; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1514 = igen_io_fire ? _GEN_490 : rob_egress_id_105; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1515 = igen_io_fire ? _GEN_491 : rob_egress_id_106; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1516 = igen_io_fire ? _GEN_492 : rob_egress_id_107; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1517 = igen_io_fire ? _GEN_493 : rob_egress_id_108; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1518 = igen_io_fire ? _GEN_494 : rob_egress_id_109; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1519 = igen_io_fire ? _GEN_495 : rob_egress_id_110; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1520 = igen_io_fire ? _GEN_496 : rob_egress_id_111; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1521 = igen_io_fire ? _GEN_497 : rob_egress_id_112; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1522 = igen_io_fire ? _GEN_498 : rob_egress_id_113; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1523 = igen_io_fire ? _GEN_499 : rob_egress_id_114; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1524 = igen_io_fire ? _GEN_500 : rob_egress_id_115; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1525 = igen_io_fire ? _GEN_501 : rob_egress_id_116; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1526 = igen_io_fire ? _GEN_502 : rob_egress_id_117; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1527 = igen_io_fire ? _GEN_503 : rob_egress_id_118; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1528 = igen_io_fire ? _GEN_504 : rob_egress_id_119; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1529 = igen_io_fire ? _GEN_505 : rob_egress_id_120; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1530 = igen_io_fire ? _GEN_506 : rob_egress_id_121; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1531 = igen_io_fire ? _GEN_507 : rob_egress_id_122; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1532 = igen_io_fire ? _GEN_508 : rob_egress_id_123; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1533 = igen_io_fire ? _GEN_509 : rob_egress_id_124; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1534 = igen_io_fire ? _GEN_510 : rob_egress_id_125; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1535 = igen_io_fire ? _GEN_511 : rob_egress_id_126; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1536 = igen_io_fire ? _GEN_512 : rob_egress_id_127; // @[TestHarness.scala 178:25 151:26]
  wire [1:0] _GEN_1537 = igen_io_fire ? _GEN_513 : rob_ingress_id_0; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1538 = igen_io_fire ? _GEN_514 : rob_ingress_id_1; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1539 = igen_io_fire ? _GEN_515 : rob_ingress_id_2; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1540 = igen_io_fire ? _GEN_516 : rob_ingress_id_3; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1541 = igen_io_fire ? _GEN_517 : rob_ingress_id_4; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1542 = igen_io_fire ? _GEN_518 : rob_ingress_id_5; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1543 = igen_io_fire ? _GEN_519 : rob_ingress_id_6; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1544 = igen_io_fire ? _GEN_520 : rob_ingress_id_7; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1545 = igen_io_fire ? _GEN_521 : rob_ingress_id_8; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1546 = igen_io_fire ? _GEN_522 : rob_ingress_id_9; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1547 = igen_io_fire ? _GEN_523 : rob_ingress_id_10; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1548 = igen_io_fire ? _GEN_524 : rob_ingress_id_11; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1549 = igen_io_fire ? _GEN_525 : rob_ingress_id_12; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1550 = igen_io_fire ? _GEN_526 : rob_ingress_id_13; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1551 = igen_io_fire ? _GEN_527 : rob_ingress_id_14; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1552 = igen_io_fire ? _GEN_528 : rob_ingress_id_15; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1553 = igen_io_fire ? _GEN_529 : rob_ingress_id_16; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1554 = igen_io_fire ? _GEN_530 : rob_ingress_id_17; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1555 = igen_io_fire ? _GEN_531 : rob_ingress_id_18; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1556 = igen_io_fire ? _GEN_532 : rob_ingress_id_19; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1557 = igen_io_fire ? _GEN_533 : rob_ingress_id_20; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1558 = igen_io_fire ? _GEN_534 : rob_ingress_id_21; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1559 = igen_io_fire ? _GEN_535 : rob_ingress_id_22; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1560 = igen_io_fire ? _GEN_536 : rob_ingress_id_23; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1561 = igen_io_fire ? _GEN_537 : rob_ingress_id_24; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1562 = igen_io_fire ? _GEN_538 : rob_ingress_id_25; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1563 = igen_io_fire ? _GEN_539 : rob_ingress_id_26; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1564 = igen_io_fire ? _GEN_540 : rob_ingress_id_27; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1565 = igen_io_fire ? _GEN_541 : rob_ingress_id_28; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1566 = igen_io_fire ? _GEN_542 : rob_ingress_id_29; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1567 = igen_io_fire ? _GEN_543 : rob_ingress_id_30; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1568 = igen_io_fire ? _GEN_544 : rob_ingress_id_31; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1569 = igen_io_fire ? _GEN_545 : rob_ingress_id_32; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1570 = igen_io_fire ? _GEN_546 : rob_ingress_id_33; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1571 = igen_io_fire ? _GEN_547 : rob_ingress_id_34; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1572 = igen_io_fire ? _GEN_548 : rob_ingress_id_35; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1573 = igen_io_fire ? _GEN_549 : rob_ingress_id_36; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1574 = igen_io_fire ? _GEN_550 : rob_ingress_id_37; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1575 = igen_io_fire ? _GEN_551 : rob_ingress_id_38; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1576 = igen_io_fire ? _GEN_552 : rob_ingress_id_39; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1577 = igen_io_fire ? _GEN_553 : rob_ingress_id_40; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1578 = igen_io_fire ? _GEN_554 : rob_ingress_id_41; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1579 = igen_io_fire ? _GEN_555 : rob_ingress_id_42; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1580 = igen_io_fire ? _GEN_556 : rob_ingress_id_43; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1581 = igen_io_fire ? _GEN_557 : rob_ingress_id_44; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1582 = igen_io_fire ? _GEN_558 : rob_ingress_id_45; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1583 = igen_io_fire ? _GEN_559 : rob_ingress_id_46; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1584 = igen_io_fire ? _GEN_560 : rob_ingress_id_47; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1585 = igen_io_fire ? _GEN_561 : rob_ingress_id_48; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1586 = igen_io_fire ? _GEN_562 : rob_ingress_id_49; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1587 = igen_io_fire ? _GEN_563 : rob_ingress_id_50; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1588 = igen_io_fire ? _GEN_564 : rob_ingress_id_51; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1589 = igen_io_fire ? _GEN_565 : rob_ingress_id_52; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1590 = igen_io_fire ? _GEN_566 : rob_ingress_id_53; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1591 = igen_io_fire ? _GEN_567 : rob_ingress_id_54; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1592 = igen_io_fire ? _GEN_568 : rob_ingress_id_55; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1593 = igen_io_fire ? _GEN_569 : rob_ingress_id_56; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1594 = igen_io_fire ? _GEN_570 : rob_ingress_id_57; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1595 = igen_io_fire ? _GEN_571 : rob_ingress_id_58; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1596 = igen_io_fire ? _GEN_572 : rob_ingress_id_59; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1597 = igen_io_fire ? _GEN_573 : rob_ingress_id_60; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1598 = igen_io_fire ? _GEN_574 : rob_ingress_id_61; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1599 = igen_io_fire ? _GEN_575 : rob_ingress_id_62; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1600 = igen_io_fire ? _GEN_576 : rob_ingress_id_63; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1601 = igen_io_fire ? _GEN_577 : rob_ingress_id_64; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1602 = igen_io_fire ? _GEN_578 : rob_ingress_id_65; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1603 = igen_io_fire ? _GEN_579 : rob_ingress_id_66; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1604 = igen_io_fire ? _GEN_580 : rob_ingress_id_67; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1605 = igen_io_fire ? _GEN_581 : rob_ingress_id_68; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1606 = igen_io_fire ? _GEN_582 : rob_ingress_id_69; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1607 = igen_io_fire ? _GEN_583 : rob_ingress_id_70; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1608 = igen_io_fire ? _GEN_584 : rob_ingress_id_71; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1609 = igen_io_fire ? _GEN_585 : rob_ingress_id_72; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1610 = igen_io_fire ? _GEN_586 : rob_ingress_id_73; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1611 = igen_io_fire ? _GEN_587 : rob_ingress_id_74; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1612 = igen_io_fire ? _GEN_588 : rob_ingress_id_75; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1613 = igen_io_fire ? _GEN_589 : rob_ingress_id_76; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1614 = igen_io_fire ? _GEN_590 : rob_ingress_id_77; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1615 = igen_io_fire ? _GEN_591 : rob_ingress_id_78; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1616 = igen_io_fire ? _GEN_592 : rob_ingress_id_79; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1617 = igen_io_fire ? _GEN_593 : rob_ingress_id_80; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1618 = igen_io_fire ? _GEN_594 : rob_ingress_id_81; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1619 = igen_io_fire ? _GEN_595 : rob_ingress_id_82; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1620 = igen_io_fire ? _GEN_596 : rob_ingress_id_83; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1621 = igen_io_fire ? _GEN_597 : rob_ingress_id_84; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1622 = igen_io_fire ? _GEN_598 : rob_ingress_id_85; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1623 = igen_io_fire ? _GEN_599 : rob_ingress_id_86; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1624 = igen_io_fire ? _GEN_600 : rob_ingress_id_87; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1625 = igen_io_fire ? _GEN_601 : rob_ingress_id_88; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1626 = igen_io_fire ? _GEN_602 : rob_ingress_id_89; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1627 = igen_io_fire ? _GEN_603 : rob_ingress_id_90; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1628 = igen_io_fire ? _GEN_604 : rob_ingress_id_91; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1629 = igen_io_fire ? _GEN_605 : rob_ingress_id_92; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1630 = igen_io_fire ? _GEN_606 : rob_ingress_id_93; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1631 = igen_io_fire ? _GEN_607 : rob_ingress_id_94; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1632 = igen_io_fire ? _GEN_608 : rob_ingress_id_95; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1633 = igen_io_fire ? _GEN_609 : rob_ingress_id_96; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1634 = igen_io_fire ? _GEN_610 : rob_ingress_id_97; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1635 = igen_io_fire ? _GEN_611 : rob_ingress_id_98; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1636 = igen_io_fire ? _GEN_612 : rob_ingress_id_99; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1637 = igen_io_fire ? _GEN_613 : rob_ingress_id_100; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1638 = igen_io_fire ? _GEN_614 : rob_ingress_id_101; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1639 = igen_io_fire ? _GEN_615 : rob_ingress_id_102; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1640 = igen_io_fire ? _GEN_616 : rob_ingress_id_103; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1641 = igen_io_fire ? _GEN_617 : rob_ingress_id_104; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1642 = igen_io_fire ? _GEN_618 : rob_ingress_id_105; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1643 = igen_io_fire ? _GEN_619 : rob_ingress_id_106; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1644 = igen_io_fire ? _GEN_620 : rob_ingress_id_107; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1645 = igen_io_fire ? _GEN_621 : rob_ingress_id_108; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1646 = igen_io_fire ? _GEN_622 : rob_ingress_id_109; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1647 = igen_io_fire ? _GEN_623 : rob_ingress_id_110; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1648 = igen_io_fire ? _GEN_624 : rob_ingress_id_111; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1649 = igen_io_fire ? _GEN_625 : rob_ingress_id_112; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1650 = igen_io_fire ? _GEN_626 : rob_ingress_id_113; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1651 = igen_io_fire ? _GEN_627 : rob_ingress_id_114; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1652 = igen_io_fire ? _GEN_628 : rob_ingress_id_115; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1653 = igen_io_fire ? _GEN_629 : rob_ingress_id_116; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1654 = igen_io_fire ? _GEN_630 : rob_ingress_id_117; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1655 = igen_io_fire ? _GEN_631 : rob_ingress_id_118; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1656 = igen_io_fire ? _GEN_632 : rob_ingress_id_119; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1657 = igen_io_fire ? _GEN_633 : rob_ingress_id_120; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1658 = igen_io_fire ? _GEN_634 : rob_ingress_id_121; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1659 = igen_io_fire ? _GEN_635 : rob_ingress_id_122; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1660 = igen_io_fire ? _GEN_636 : rob_ingress_id_123; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1661 = igen_io_fire ? _GEN_637 : rob_ingress_id_124; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1662 = igen_io_fire ? _GEN_638 : rob_ingress_id_125; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1663 = igen_io_fire ? _GEN_639 : rob_ingress_id_126; // @[TestHarness.scala 178:25 152:27]
  wire [1:0] _GEN_1664 = igen_io_fire ? _GEN_640 : rob_ingress_id_127; // @[TestHarness.scala 178:25 152:27]
  wire [3:0] _GEN_1665 = igen_io_fire ? _GEN_641 : rob_n_flits_0; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1666 = igen_io_fire ? _GEN_642 : rob_n_flits_1; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1667 = igen_io_fire ? _GEN_643 : rob_n_flits_2; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1668 = igen_io_fire ? _GEN_644 : rob_n_flits_3; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1669 = igen_io_fire ? _GEN_645 : rob_n_flits_4; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1670 = igen_io_fire ? _GEN_646 : rob_n_flits_5; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1671 = igen_io_fire ? _GEN_647 : rob_n_flits_6; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1672 = igen_io_fire ? _GEN_648 : rob_n_flits_7; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1673 = igen_io_fire ? _GEN_649 : rob_n_flits_8; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1674 = igen_io_fire ? _GEN_650 : rob_n_flits_9; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1675 = igen_io_fire ? _GEN_651 : rob_n_flits_10; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1676 = igen_io_fire ? _GEN_652 : rob_n_flits_11; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1677 = igen_io_fire ? _GEN_653 : rob_n_flits_12; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1678 = igen_io_fire ? _GEN_654 : rob_n_flits_13; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1679 = igen_io_fire ? _GEN_655 : rob_n_flits_14; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1680 = igen_io_fire ? _GEN_656 : rob_n_flits_15; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1681 = igen_io_fire ? _GEN_657 : rob_n_flits_16; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1682 = igen_io_fire ? _GEN_658 : rob_n_flits_17; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1683 = igen_io_fire ? _GEN_659 : rob_n_flits_18; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1684 = igen_io_fire ? _GEN_660 : rob_n_flits_19; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1685 = igen_io_fire ? _GEN_661 : rob_n_flits_20; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1686 = igen_io_fire ? _GEN_662 : rob_n_flits_21; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1687 = igen_io_fire ? _GEN_663 : rob_n_flits_22; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1688 = igen_io_fire ? _GEN_664 : rob_n_flits_23; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1689 = igen_io_fire ? _GEN_665 : rob_n_flits_24; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1690 = igen_io_fire ? _GEN_666 : rob_n_flits_25; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1691 = igen_io_fire ? _GEN_667 : rob_n_flits_26; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1692 = igen_io_fire ? _GEN_668 : rob_n_flits_27; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1693 = igen_io_fire ? _GEN_669 : rob_n_flits_28; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1694 = igen_io_fire ? _GEN_670 : rob_n_flits_29; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1695 = igen_io_fire ? _GEN_671 : rob_n_flits_30; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1696 = igen_io_fire ? _GEN_672 : rob_n_flits_31; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1697 = igen_io_fire ? _GEN_673 : rob_n_flits_32; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1698 = igen_io_fire ? _GEN_674 : rob_n_flits_33; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1699 = igen_io_fire ? _GEN_675 : rob_n_flits_34; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1700 = igen_io_fire ? _GEN_676 : rob_n_flits_35; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1701 = igen_io_fire ? _GEN_677 : rob_n_flits_36; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1702 = igen_io_fire ? _GEN_678 : rob_n_flits_37; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1703 = igen_io_fire ? _GEN_679 : rob_n_flits_38; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1704 = igen_io_fire ? _GEN_680 : rob_n_flits_39; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1705 = igen_io_fire ? _GEN_681 : rob_n_flits_40; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1706 = igen_io_fire ? _GEN_682 : rob_n_flits_41; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1707 = igen_io_fire ? _GEN_683 : rob_n_flits_42; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1708 = igen_io_fire ? _GEN_684 : rob_n_flits_43; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1709 = igen_io_fire ? _GEN_685 : rob_n_flits_44; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1710 = igen_io_fire ? _GEN_686 : rob_n_flits_45; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1711 = igen_io_fire ? _GEN_687 : rob_n_flits_46; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1712 = igen_io_fire ? _GEN_688 : rob_n_flits_47; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1713 = igen_io_fire ? _GEN_689 : rob_n_flits_48; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1714 = igen_io_fire ? _GEN_690 : rob_n_flits_49; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1715 = igen_io_fire ? _GEN_691 : rob_n_flits_50; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1716 = igen_io_fire ? _GEN_692 : rob_n_flits_51; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1717 = igen_io_fire ? _GEN_693 : rob_n_flits_52; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1718 = igen_io_fire ? _GEN_694 : rob_n_flits_53; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1719 = igen_io_fire ? _GEN_695 : rob_n_flits_54; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1720 = igen_io_fire ? _GEN_696 : rob_n_flits_55; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1721 = igen_io_fire ? _GEN_697 : rob_n_flits_56; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1722 = igen_io_fire ? _GEN_698 : rob_n_flits_57; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1723 = igen_io_fire ? _GEN_699 : rob_n_flits_58; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1724 = igen_io_fire ? _GEN_700 : rob_n_flits_59; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1725 = igen_io_fire ? _GEN_701 : rob_n_flits_60; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1726 = igen_io_fire ? _GEN_702 : rob_n_flits_61; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1727 = igen_io_fire ? _GEN_703 : rob_n_flits_62; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1728 = igen_io_fire ? _GEN_704 : rob_n_flits_63; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1729 = igen_io_fire ? _GEN_705 : rob_n_flits_64; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1730 = igen_io_fire ? _GEN_706 : rob_n_flits_65; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1731 = igen_io_fire ? _GEN_707 : rob_n_flits_66; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1732 = igen_io_fire ? _GEN_708 : rob_n_flits_67; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1733 = igen_io_fire ? _GEN_709 : rob_n_flits_68; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1734 = igen_io_fire ? _GEN_710 : rob_n_flits_69; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1735 = igen_io_fire ? _GEN_711 : rob_n_flits_70; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1736 = igen_io_fire ? _GEN_712 : rob_n_flits_71; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1737 = igen_io_fire ? _GEN_713 : rob_n_flits_72; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1738 = igen_io_fire ? _GEN_714 : rob_n_flits_73; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1739 = igen_io_fire ? _GEN_715 : rob_n_flits_74; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1740 = igen_io_fire ? _GEN_716 : rob_n_flits_75; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1741 = igen_io_fire ? _GEN_717 : rob_n_flits_76; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1742 = igen_io_fire ? _GEN_718 : rob_n_flits_77; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1743 = igen_io_fire ? _GEN_719 : rob_n_flits_78; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1744 = igen_io_fire ? _GEN_720 : rob_n_flits_79; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1745 = igen_io_fire ? _GEN_721 : rob_n_flits_80; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1746 = igen_io_fire ? _GEN_722 : rob_n_flits_81; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1747 = igen_io_fire ? _GEN_723 : rob_n_flits_82; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1748 = igen_io_fire ? _GEN_724 : rob_n_flits_83; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1749 = igen_io_fire ? _GEN_725 : rob_n_flits_84; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1750 = igen_io_fire ? _GEN_726 : rob_n_flits_85; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1751 = igen_io_fire ? _GEN_727 : rob_n_flits_86; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1752 = igen_io_fire ? _GEN_728 : rob_n_flits_87; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1753 = igen_io_fire ? _GEN_729 : rob_n_flits_88; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1754 = igen_io_fire ? _GEN_730 : rob_n_flits_89; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1755 = igen_io_fire ? _GEN_731 : rob_n_flits_90; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1756 = igen_io_fire ? _GEN_732 : rob_n_flits_91; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1757 = igen_io_fire ? _GEN_733 : rob_n_flits_92; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1758 = igen_io_fire ? _GEN_734 : rob_n_flits_93; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1759 = igen_io_fire ? _GEN_735 : rob_n_flits_94; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1760 = igen_io_fire ? _GEN_736 : rob_n_flits_95; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1761 = igen_io_fire ? _GEN_737 : rob_n_flits_96; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1762 = igen_io_fire ? _GEN_738 : rob_n_flits_97; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1763 = igen_io_fire ? _GEN_739 : rob_n_flits_98; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1764 = igen_io_fire ? _GEN_740 : rob_n_flits_99; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1765 = igen_io_fire ? _GEN_741 : rob_n_flits_100; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1766 = igen_io_fire ? _GEN_742 : rob_n_flits_101; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1767 = igen_io_fire ? _GEN_743 : rob_n_flits_102; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1768 = igen_io_fire ? _GEN_744 : rob_n_flits_103; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1769 = igen_io_fire ? _GEN_745 : rob_n_flits_104; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1770 = igen_io_fire ? _GEN_746 : rob_n_flits_105; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1771 = igen_io_fire ? _GEN_747 : rob_n_flits_106; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1772 = igen_io_fire ? _GEN_748 : rob_n_flits_107; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1773 = igen_io_fire ? _GEN_749 : rob_n_flits_108; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1774 = igen_io_fire ? _GEN_750 : rob_n_flits_109; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1775 = igen_io_fire ? _GEN_751 : rob_n_flits_110; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1776 = igen_io_fire ? _GEN_752 : rob_n_flits_111; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1777 = igen_io_fire ? _GEN_753 : rob_n_flits_112; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1778 = igen_io_fire ? _GEN_754 : rob_n_flits_113; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1779 = igen_io_fire ? _GEN_755 : rob_n_flits_114; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1780 = igen_io_fire ? _GEN_756 : rob_n_flits_115; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1781 = igen_io_fire ? _GEN_757 : rob_n_flits_116; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1782 = igen_io_fire ? _GEN_758 : rob_n_flits_117; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1783 = igen_io_fire ? _GEN_759 : rob_n_flits_118; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1784 = igen_io_fire ? _GEN_760 : rob_n_flits_119; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1785 = igen_io_fire ? _GEN_761 : rob_n_flits_120; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1786 = igen_io_fire ? _GEN_762 : rob_n_flits_121; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1787 = igen_io_fire ? _GEN_763 : rob_n_flits_122; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1788 = igen_io_fire ? _GEN_764 : rob_n_flits_123; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1789 = igen_io_fire ? _GEN_765 : rob_n_flits_124; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1790 = igen_io_fire ? _GEN_766 : rob_n_flits_125; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1791 = igen_io_fire ? _GEN_767 : rob_n_flits_126; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1792 = igen_io_fire ? _GEN_768 : rob_n_flits_127; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1793 = igen_io_fire ? _GEN_769 : rob_flits_returned_0; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1794 = igen_io_fire ? _GEN_770 : rob_flits_returned_1; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1795 = igen_io_fire ? _GEN_771 : rob_flits_returned_2; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1796 = igen_io_fire ? _GEN_772 : rob_flits_returned_3; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1797 = igen_io_fire ? _GEN_773 : rob_flits_returned_4; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1798 = igen_io_fire ? _GEN_774 : rob_flits_returned_5; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1799 = igen_io_fire ? _GEN_775 : rob_flits_returned_6; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1800 = igen_io_fire ? _GEN_776 : rob_flits_returned_7; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1801 = igen_io_fire ? _GEN_777 : rob_flits_returned_8; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1802 = igen_io_fire ? _GEN_778 : rob_flits_returned_9; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1803 = igen_io_fire ? _GEN_779 : rob_flits_returned_10; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1804 = igen_io_fire ? _GEN_780 : rob_flits_returned_11; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1805 = igen_io_fire ? _GEN_781 : rob_flits_returned_12; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1806 = igen_io_fire ? _GEN_782 : rob_flits_returned_13; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1807 = igen_io_fire ? _GEN_783 : rob_flits_returned_14; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1808 = igen_io_fire ? _GEN_784 : rob_flits_returned_15; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1809 = igen_io_fire ? _GEN_785 : rob_flits_returned_16; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1810 = igen_io_fire ? _GEN_786 : rob_flits_returned_17; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1811 = igen_io_fire ? _GEN_787 : rob_flits_returned_18; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1812 = igen_io_fire ? _GEN_788 : rob_flits_returned_19; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1813 = igen_io_fire ? _GEN_789 : rob_flits_returned_20; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1814 = igen_io_fire ? _GEN_790 : rob_flits_returned_21; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1815 = igen_io_fire ? _GEN_791 : rob_flits_returned_22; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1816 = igen_io_fire ? _GEN_792 : rob_flits_returned_23; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1817 = igen_io_fire ? _GEN_793 : rob_flits_returned_24; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1818 = igen_io_fire ? _GEN_794 : rob_flits_returned_25; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1819 = igen_io_fire ? _GEN_795 : rob_flits_returned_26; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1820 = igen_io_fire ? _GEN_796 : rob_flits_returned_27; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1821 = igen_io_fire ? _GEN_797 : rob_flits_returned_28; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1822 = igen_io_fire ? _GEN_798 : rob_flits_returned_29; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1823 = igen_io_fire ? _GEN_799 : rob_flits_returned_30; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1824 = igen_io_fire ? _GEN_800 : rob_flits_returned_31; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1825 = igen_io_fire ? _GEN_801 : rob_flits_returned_32; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1826 = igen_io_fire ? _GEN_802 : rob_flits_returned_33; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1827 = igen_io_fire ? _GEN_803 : rob_flits_returned_34; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1828 = igen_io_fire ? _GEN_804 : rob_flits_returned_35; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1829 = igen_io_fire ? _GEN_805 : rob_flits_returned_36; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1830 = igen_io_fire ? _GEN_806 : rob_flits_returned_37; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1831 = igen_io_fire ? _GEN_807 : rob_flits_returned_38; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1832 = igen_io_fire ? _GEN_808 : rob_flits_returned_39; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1833 = igen_io_fire ? _GEN_809 : rob_flits_returned_40; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1834 = igen_io_fire ? _GEN_810 : rob_flits_returned_41; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1835 = igen_io_fire ? _GEN_811 : rob_flits_returned_42; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1836 = igen_io_fire ? _GEN_812 : rob_flits_returned_43; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1837 = igen_io_fire ? _GEN_813 : rob_flits_returned_44; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1838 = igen_io_fire ? _GEN_814 : rob_flits_returned_45; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1839 = igen_io_fire ? _GEN_815 : rob_flits_returned_46; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1840 = igen_io_fire ? _GEN_816 : rob_flits_returned_47; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1841 = igen_io_fire ? _GEN_817 : rob_flits_returned_48; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1842 = igen_io_fire ? _GEN_818 : rob_flits_returned_49; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1843 = igen_io_fire ? _GEN_819 : rob_flits_returned_50; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1844 = igen_io_fire ? _GEN_820 : rob_flits_returned_51; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1845 = igen_io_fire ? _GEN_821 : rob_flits_returned_52; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1846 = igen_io_fire ? _GEN_822 : rob_flits_returned_53; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1847 = igen_io_fire ? _GEN_823 : rob_flits_returned_54; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1848 = igen_io_fire ? _GEN_824 : rob_flits_returned_55; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1849 = igen_io_fire ? _GEN_825 : rob_flits_returned_56; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1850 = igen_io_fire ? _GEN_826 : rob_flits_returned_57; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1851 = igen_io_fire ? _GEN_827 : rob_flits_returned_58; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1852 = igen_io_fire ? _GEN_828 : rob_flits_returned_59; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1853 = igen_io_fire ? _GEN_829 : rob_flits_returned_60; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1854 = igen_io_fire ? _GEN_830 : rob_flits_returned_61; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1855 = igen_io_fire ? _GEN_831 : rob_flits_returned_62; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1856 = igen_io_fire ? _GEN_832 : rob_flits_returned_63; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1857 = igen_io_fire ? _GEN_833 : rob_flits_returned_64; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1858 = igen_io_fire ? _GEN_834 : rob_flits_returned_65; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1859 = igen_io_fire ? _GEN_835 : rob_flits_returned_66; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1860 = igen_io_fire ? _GEN_836 : rob_flits_returned_67; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1861 = igen_io_fire ? _GEN_837 : rob_flits_returned_68; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1862 = igen_io_fire ? _GEN_838 : rob_flits_returned_69; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1863 = igen_io_fire ? _GEN_839 : rob_flits_returned_70; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1864 = igen_io_fire ? _GEN_840 : rob_flits_returned_71; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1865 = igen_io_fire ? _GEN_841 : rob_flits_returned_72; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1866 = igen_io_fire ? _GEN_842 : rob_flits_returned_73; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1867 = igen_io_fire ? _GEN_843 : rob_flits_returned_74; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1868 = igen_io_fire ? _GEN_844 : rob_flits_returned_75; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1869 = igen_io_fire ? _GEN_845 : rob_flits_returned_76; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1870 = igen_io_fire ? _GEN_846 : rob_flits_returned_77; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1871 = igen_io_fire ? _GEN_847 : rob_flits_returned_78; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1872 = igen_io_fire ? _GEN_848 : rob_flits_returned_79; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1873 = igen_io_fire ? _GEN_849 : rob_flits_returned_80; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1874 = igen_io_fire ? _GEN_850 : rob_flits_returned_81; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1875 = igen_io_fire ? _GEN_851 : rob_flits_returned_82; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1876 = igen_io_fire ? _GEN_852 : rob_flits_returned_83; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1877 = igen_io_fire ? _GEN_853 : rob_flits_returned_84; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1878 = igen_io_fire ? _GEN_854 : rob_flits_returned_85; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1879 = igen_io_fire ? _GEN_855 : rob_flits_returned_86; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1880 = igen_io_fire ? _GEN_856 : rob_flits_returned_87; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1881 = igen_io_fire ? _GEN_857 : rob_flits_returned_88; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1882 = igen_io_fire ? _GEN_858 : rob_flits_returned_89; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1883 = igen_io_fire ? _GEN_859 : rob_flits_returned_90; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1884 = igen_io_fire ? _GEN_860 : rob_flits_returned_91; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1885 = igen_io_fire ? _GEN_861 : rob_flits_returned_92; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1886 = igen_io_fire ? _GEN_862 : rob_flits_returned_93; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1887 = igen_io_fire ? _GEN_863 : rob_flits_returned_94; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1888 = igen_io_fire ? _GEN_864 : rob_flits_returned_95; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1889 = igen_io_fire ? _GEN_865 : rob_flits_returned_96; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1890 = igen_io_fire ? _GEN_866 : rob_flits_returned_97; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1891 = igen_io_fire ? _GEN_867 : rob_flits_returned_98; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1892 = igen_io_fire ? _GEN_868 : rob_flits_returned_99; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1893 = igen_io_fire ? _GEN_869 : rob_flits_returned_100; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1894 = igen_io_fire ? _GEN_870 : rob_flits_returned_101; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1895 = igen_io_fire ? _GEN_871 : rob_flits_returned_102; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1896 = igen_io_fire ? _GEN_872 : rob_flits_returned_103; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1897 = igen_io_fire ? _GEN_873 : rob_flits_returned_104; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1898 = igen_io_fire ? _GEN_874 : rob_flits_returned_105; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1899 = igen_io_fire ? _GEN_875 : rob_flits_returned_106; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1900 = igen_io_fire ? _GEN_876 : rob_flits_returned_107; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1901 = igen_io_fire ? _GEN_877 : rob_flits_returned_108; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1902 = igen_io_fire ? _GEN_878 : rob_flits_returned_109; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1903 = igen_io_fire ? _GEN_879 : rob_flits_returned_110; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1904 = igen_io_fire ? _GEN_880 : rob_flits_returned_111; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1905 = igen_io_fire ? _GEN_881 : rob_flits_returned_112; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1906 = igen_io_fire ? _GEN_882 : rob_flits_returned_113; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1907 = igen_io_fire ? _GEN_883 : rob_flits_returned_114; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1908 = igen_io_fire ? _GEN_884 : rob_flits_returned_115; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1909 = igen_io_fire ? _GEN_885 : rob_flits_returned_116; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1910 = igen_io_fire ? _GEN_886 : rob_flits_returned_117; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1911 = igen_io_fire ? _GEN_887 : rob_flits_returned_118; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1912 = igen_io_fire ? _GEN_888 : rob_flits_returned_119; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1913 = igen_io_fire ? _GEN_889 : rob_flits_returned_120; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1914 = igen_io_fire ? _GEN_890 : rob_flits_returned_121; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1915 = igen_io_fire ? _GEN_891 : rob_flits_returned_122; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1916 = igen_io_fire ? _GEN_892 : rob_flits_returned_123; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1917 = igen_io_fire ? _GEN_893 : rob_flits_returned_124; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1918 = igen_io_fire ? _GEN_894 : rob_flits_returned_125; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1919 = igen_io_fire ? _GEN_895 : rob_flits_returned_126; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1920 = igen_io_fire ? _GEN_896 : rob_flits_returned_127; // @[TestHarness.scala 178:25 154:31]
  wire [63:0] _GEN_1921 = igen_io_fire ? _GEN_897 : rob_tscs_0; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1922 = igen_io_fire ? _GEN_898 : rob_tscs_1; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1923 = igen_io_fire ? _GEN_899 : rob_tscs_2; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1924 = igen_io_fire ? _GEN_900 : rob_tscs_3; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1925 = igen_io_fire ? _GEN_901 : rob_tscs_4; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1926 = igen_io_fire ? _GEN_902 : rob_tscs_5; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1927 = igen_io_fire ? _GEN_903 : rob_tscs_6; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1928 = igen_io_fire ? _GEN_904 : rob_tscs_7; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1929 = igen_io_fire ? _GEN_905 : rob_tscs_8; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1930 = igen_io_fire ? _GEN_906 : rob_tscs_9; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1931 = igen_io_fire ? _GEN_907 : rob_tscs_10; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1932 = igen_io_fire ? _GEN_908 : rob_tscs_11; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1933 = igen_io_fire ? _GEN_909 : rob_tscs_12; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1934 = igen_io_fire ? _GEN_910 : rob_tscs_13; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1935 = igen_io_fire ? _GEN_911 : rob_tscs_14; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1936 = igen_io_fire ? _GEN_912 : rob_tscs_15; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1937 = igen_io_fire ? _GEN_913 : rob_tscs_16; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1938 = igen_io_fire ? _GEN_914 : rob_tscs_17; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1939 = igen_io_fire ? _GEN_915 : rob_tscs_18; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1940 = igen_io_fire ? _GEN_916 : rob_tscs_19; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1941 = igen_io_fire ? _GEN_917 : rob_tscs_20; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1942 = igen_io_fire ? _GEN_918 : rob_tscs_21; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1943 = igen_io_fire ? _GEN_919 : rob_tscs_22; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1944 = igen_io_fire ? _GEN_920 : rob_tscs_23; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1945 = igen_io_fire ? _GEN_921 : rob_tscs_24; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1946 = igen_io_fire ? _GEN_922 : rob_tscs_25; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1947 = igen_io_fire ? _GEN_923 : rob_tscs_26; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1948 = igen_io_fire ? _GEN_924 : rob_tscs_27; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1949 = igen_io_fire ? _GEN_925 : rob_tscs_28; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1950 = igen_io_fire ? _GEN_926 : rob_tscs_29; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1951 = igen_io_fire ? _GEN_927 : rob_tscs_30; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1952 = igen_io_fire ? _GEN_928 : rob_tscs_31; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1953 = igen_io_fire ? _GEN_929 : rob_tscs_32; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1954 = igen_io_fire ? _GEN_930 : rob_tscs_33; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1955 = igen_io_fire ? _GEN_931 : rob_tscs_34; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1956 = igen_io_fire ? _GEN_932 : rob_tscs_35; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1957 = igen_io_fire ? _GEN_933 : rob_tscs_36; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1958 = igen_io_fire ? _GEN_934 : rob_tscs_37; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1959 = igen_io_fire ? _GEN_935 : rob_tscs_38; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1960 = igen_io_fire ? _GEN_936 : rob_tscs_39; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1961 = igen_io_fire ? _GEN_937 : rob_tscs_40; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1962 = igen_io_fire ? _GEN_938 : rob_tscs_41; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1963 = igen_io_fire ? _GEN_939 : rob_tscs_42; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1964 = igen_io_fire ? _GEN_940 : rob_tscs_43; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1965 = igen_io_fire ? _GEN_941 : rob_tscs_44; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1966 = igen_io_fire ? _GEN_942 : rob_tscs_45; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1967 = igen_io_fire ? _GEN_943 : rob_tscs_46; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1968 = igen_io_fire ? _GEN_944 : rob_tscs_47; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1969 = igen_io_fire ? _GEN_945 : rob_tscs_48; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1970 = igen_io_fire ? _GEN_946 : rob_tscs_49; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1971 = igen_io_fire ? _GEN_947 : rob_tscs_50; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1972 = igen_io_fire ? _GEN_948 : rob_tscs_51; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1973 = igen_io_fire ? _GEN_949 : rob_tscs_52; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1974 = igen_io_fire ? _GEN_950 : rob_tscs_53; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1975 = igen_io_fire ? _GEN_951 : rob_tscs_54; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1976 = igen_io_fire ? _GEN_952 : rob_tscs_55; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1977 = igen_io_fire ? _GEN_953 : rob_tscs_56; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1978 = igen_io_fire ? _GEN_954 : rob_tscs_57; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1979 = igen_io_fire ? _GEN_955 : rob_tscs_58; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1980 = igen_io_fire ? _GEN_956 : rob_tscs_59; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1981 = igen_io_fire ? _GEN_957 : rob_tscs_60; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1982 = igen_io_fire ? _GEN_958 : rob_tscs_61; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1983 = igen_io_fire ? _GEN_959 : rob_tscs_62; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1984 = igen_io_fire ? _GEN_960 : rob_tscs_63; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1985 = igen_io_fire ? _GEN_961 : rob_tscs_64; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1986 = igen_io_fire ? _GEN_962 : rob_tscs_65; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1987 = igen_io_fire ? _GEN_963 : rob_tscs_66; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1988 = igen_io_fire ? _GEN_964 : rob_tscs_67; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1989 = igen_io_fire ? _GEN_965 : rob_tscs_68; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1990 = igen_io_fire ? _GEN_966 : rob_tscs_69; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1991 = igen_io_fire ? _GEN_967 : rob_tscs_70; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1992 = igen_io_fire ? _GEN_968 : rob_tscs_71; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1993 = igen_io_fire ? _GEN_969 : rob_tscs_72; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1994 = igen_io_fire ? _GEN_970 : rob_tscs_73; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1995 = igen_io_fire ? _GEN_971 : rob_tscs_74; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1996 = igen_io_fire ? _GEN_972 : rob_tscs_75; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1997 = igen_io_fire ? _GEN_973 : rob_tscs_76; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1998 = igen_io_fire ? _GEN_974 : rob_tscs_77; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1999 = igen_io_fire ? _GEN_975 : rob_tscs_78; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2000 = igen_io_fire ? _GEN_976 : rob_tscs_79; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2001 = igen_io_fire ? _GEN_977 : rob_tscs_80; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2002 = igen_io_fire ? _GEN_978 : rob_tscs_81; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2003 = igen_io_fire ? _GEN_979 : rob_tscs_82; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2004 = igen_io_fire ? _GEN_980 : rob_tscs_83; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2005 = igen_io_fire ? _GEN_981 : rob_tscs_84; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2006 = igen_io_fire ? _GEN_982 : rob_tscs_85; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2007 = igen_io_fire ? _GEN_983 : rob_tscs_86; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2008 = igen_io_fire ? _GEN_984 : rob_tscs_87; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2009 = igen_io_fire ? _GEN_985 : rob_tscs_88; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2010 = igen_io_fire ? _GEN_986 : rob_tscs_89; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2011 = igen_io_fire ? _GEN_987 : rob_tscs_90; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2012 = igen_io_fire ? _GEN_988 : rob_tscs_91; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2013 = igen_io_fire ? _GEN_989 : rob_tscs_92; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2014 = igen_io_fire ? _GEN_990 : rob_tscs_93; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2015 = igen_io_fire ? _GEN_991 : rob_tscs_94; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2016 = igen_io_fire ? _GEN_992 : rob_tscs_95; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2017 = igen_io_fire ? _GEN_993 : rob_tscs_96; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2018 = igen_io_fire ? _GEN_994 : rob_tscs_97; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2019 = igen_io_fire ? _GEN_995 : rob_tscs_98; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2020 = igen_io_fire ? _GEN_996 : rob_tscs_99; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2021 = igen_io_fire ? _GEN_997 : rob_tscs_100; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2022 = igen_io_fire ? _GEN_998 : rob_tscs_101; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2023 = igen_io_fire ? _GEN_999 : rob_tscs_102; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2024 = igen_io_fire ? _GEN_1000 : rob_tscs_103; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2025 = igen_io_fire ? _GEN_1001 : rob_tscs_104; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2026 = igen_io_fire ? _GEN_1002 : rob_tscs_105; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2027 = igen_io_fire ? _GEN_1003 : rob_tscs_106; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2028 = igen_io_fire ? _GEN_1004 : rob_tscs_107; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2029 = igen_io_fire ? _GEN_1005 : rob_tscs_108; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2030 = igen_io_fire ? _GEN_1006 : rob_tscs_109; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2031 = igen_io_fire ? _GEN_1007 : rob_tscs_110; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2032 = igen_io_fire ? _GEN_1008 : rob_tscs_111; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2033 = igen_io_fire ? _GEN_1009 : rob_tscs_112; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2034 = igen_io_fire ? _GEN_1010 : rob_tscs_113; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2035 = igen_io_fire ? _GEN_1011 : rob_tscs_114; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2036 = igen_io_fire ? _GEN_1012 : rob_tscs_115; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2037 = igen_io_fire ? _GEN_1013 : rob_tscs_116; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2038 = igen_io_fire ? _GEN_1014 : rob_tscs_117; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2039 = igen_io_fire ? _GEN_1015 : rob_tscs_118; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2040 = igen_io_fire ? _GEN_1016 : rob_tscs_119; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2041 = igen_io_fire ? _GEN_1017 : rob_tscs_120; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2042 = igen_io_fire ? _GEN_1018 : rob_tscs_121; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2043 = igen_io_fire ? _GEN_1019 : rob_tscs_122; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2044 = igen_io_fire ? _GEN_1020 : rob_tscs_123; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2045 = igen_io_fire ? _GEN_1021 : rob_tscs_124; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2046 = igen_io_fire ? _GEN_1022 : rob_tscs_125; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2047 = igen_io_fire ? _GEN_1023 : rob_tscs_126; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2048 = igen_io_fire ? _GEN_1024 : rob_tscs_127; // @[TestHarness.scala 155:21 178:25]
  wire  _igen_io_rob_ready_T_7 = rob_alloc_avail_1 & rob_alloc_fires_1 & _igen_io_rob_ready_T_1; // @[TestHarness.scala 174:72]
  wire [63:0] _rob_payload_WIRE_3 = igen_1_io_out_bits_payload; // @[TestHarness.scala 179:{72,72}]
  wire [31:0] _GEN_2049 = 7'h0 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1025; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2050 = 7'h1 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1026; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2051 = 7'h2 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1027; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2052 = 7'h3 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1028; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2053 = 7'h4 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1029; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2054 = 7'h5 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1030; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2055 = 7'h6 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1031; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2056 = 7'h7 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1032; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2057 = 7'h8 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1033; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2058 = 7'h9 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1034; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2059 = 7'ha == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1035; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2060 = 7'hb == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1036; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2061 = 7'hc == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1037; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2062 = 7'hd == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1038; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2063 = 7'he == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1039; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2064 = 7'hf == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1040; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2065 = 7'h10 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1041; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2066 = 7'h11 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1042; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2067 = 7'h12 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1043; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2068 = 7'h13 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1044; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2069 = 7'h14 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1045; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2070 = 7'h15 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1046; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2071 = 7'h16 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1047; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2072 = 7'h17 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1048; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2073 = 7'h18 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1049; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2074 = 7'h19 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1050; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2075 = 7'h1a == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1051; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2076 = 7'h1b == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1052; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2077 = 7'h1c == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1053; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2078 = 7'h1d == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1054; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2079 = 7'h1e == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1055; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2080 = 7'h1f == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1056; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2081 = 7'h20 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1057; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2082 = 7'h21 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1058; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2083 = 7'h22 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1059; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2084 = 7'h23 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1060; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2085 = 7'h24 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1061; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2086 = 7'h25 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1062; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2087 = 7'h26 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1063; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2088 = 7'h27 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1064; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2089 = 7'h28 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1065; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2090 = 7'h29 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1066; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2091 = 7'h2a == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1067; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2092 = 7'h2b == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1068; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2093 = 7'h2c == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1069; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2094 = 7'h2d == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1070; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2095 = 7'h2e == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1071; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2096 = 7'h2f == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1072; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2097 = 7'h30 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1073; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2098 = 7'h31 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1074; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2099 = 7'h32 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1075; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2100 = 7'h33 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1076; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2101 = 7'h34 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1077; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2102 = 7'h35 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1078; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2103 = 7'h36 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1079; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2104 = 7'h37 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1080; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2105 = 7'h38 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1081; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2106 = 7'h39 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1082; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2107 = 7'h3a == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1083; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2108 = 7'h3b == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1084; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2109 = 7'h3c == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1085; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2110 = 7'h3d == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1086; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2111 = 7'h3e == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1087; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2112 = 7'h3f == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1088; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2113 = 7'h40 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1089; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2114 = 7'h41 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1090; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2115 = 7'h42 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1091; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2116 = 7'h43 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1092; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2117 = 7'h44 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1093; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2118 = 7'h45 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1094; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2119 = 7'h46 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1095; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2120 = 7'h47 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1096; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2121 = 7'h48 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1097; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2122 = 7'h49 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1098; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2123 = 7'h4a == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1099; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2124 = 7'h4b == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1100; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2125 = 7'h4c == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1101; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2126 = 7'h4d == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1102; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2127 = 7'h4e == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1103; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2128 = 7'h4f == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1104; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2129 = 7'h50 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1105; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2130 = 7'h51 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1106; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2131 = 7'h52 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1107; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2132 = 7'h53 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1108; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2133 = 7'h54 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1109; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2134 = 7'h55 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1110; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2135 = 7'h56 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1111; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2136 = 7'h57 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1112; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2137 = 7'h58 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1113; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2138 = 7'h59 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1114; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2139 = 7'h5a == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1115; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2140 = 7'h5b == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1116; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2141 = 7'h5c == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1117; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2142 = 7'h5d == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1118; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2143 = 7'h5e == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1119; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2144 = 7'h5f == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1120; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2145 = 7'h60 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1121; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2146 = 7'h61 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1122; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2147 = 7'h62 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1123; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2148 = 7'h63 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1124; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2149 = 7'h64 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1125; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2150 = 7'h65 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1126; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2151 = 7'h66 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1127; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2152 = 7'h67 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1128; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2153 = 7'h68 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1129; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2154 = 7'h69 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1130; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2155 = 7'h6a == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1131; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2156 = 7'h6b == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1132; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2157 = 7'h6c == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1133; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2158 = 7'h6d == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1134; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2159 = 7'h6e == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1135; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2160 = 7'h6f == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1136; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2161 = 7'h70 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1137; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2162 = 7'h71 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1138; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2163 = 7'h72 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1139; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2164 = 7'h73 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1140; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2165 = 7'h74 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1141; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2166 = 7'h75 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1142; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2167 = 7'h76 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1143; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2168 = 7'h77 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1144; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2169 = 7'h78 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1145; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2170 = 7'h79 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1146; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2171 = 7'h7a == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1147; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2172 = 7'h7b == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1148; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2173 = 7'h7c == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1149; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2174 = 7'h7d == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1150; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2175 = 7'h7e == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1151; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_2176 = 7'h7f == rob_alloc_ids_1 ? _rob_payload_WIRE_3[63:32] : _GEN_1152; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2177 = 7'h0 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1153; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2178 = 7'h1 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1154; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2179 = 7'h2 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1155; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2180 = 7'h3 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1156; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2181 = 7'h4 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1157; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2182 = 7'h5 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1158; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2183 = 7'h6 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1159; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2184 = 7'h7 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1160; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2185 = 7'h8 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1161; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2186 = 7'h9 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1162; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2187 = 7'ha == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1163; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2188 = 7'hb == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1164; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2189 = 7'hc == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1165; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2190 = 7'hd == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1166; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2191 = 7'he == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1167; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2192 = 7'hf == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1168; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2193 = 7'h10 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1169; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2194 = 7'h11 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1170; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2195 = 7'h12 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1171; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2196 = 7'h13 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1172; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2197 = 7'h14 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1173; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2198 = 7'h15 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1174; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2199 = 7'h16 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1175; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2200 = 7'h17 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1176; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2201 = 7'h18 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1177; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2202 = 7'h19 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1178; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2203 = 7'h1a == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1179; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2204 = 7'h1b == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1180; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2205 = 7'h1c == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1181; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2206 = 7'h1d == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1182; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2207 = 7'h1e == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1183; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2208 = 7'h1f == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1184; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2209 = 7'h20 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1185; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2210 = 7'h21 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1186; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2211 = 7'h22 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1187; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2212 = 7'h23 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1188; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2213 = 7'h24 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1189; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2214 = 7'h25 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1190; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2215 = 7'h26 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1191; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2216 = 7'h27 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1192; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2217 = 7'h28 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1193; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2218 = 7'h29 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1194; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2219 = 7'h2a == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1195; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2220 = 7'h2b == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1196; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2221 = 7'h2c == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1197; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2222 = 7'h2d == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1198; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2223 = 7'h2e == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1199; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2224 = 7'h2f == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1200; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2225 = 7'h30 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1201; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2226 = 7'h31 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1202; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2227 = 7'h32 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1203; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2228 = 7'h33 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1204; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2229 = 7'h34 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1205; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2230 = 7'h35 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1206; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2231 = 7'h36 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1207; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2232 = 7'h37 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1208; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2233 = 7'h38 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1209; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2234 = 7'h39 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1210; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2235 = 7'h3a == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1211; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2236 = 7'h3b == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1212; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2237 = 7'h3c == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1213; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2238 = 7'h3d == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1214; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2239 = 7'h3e == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1215; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2240 = 7'h3f == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1216; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2241 = 7'h40 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1217; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2242 = 7'h41 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1218; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2243 = 7'h42 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1219; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2244 = 7'h43 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1220; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2245 = 7'h44 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1221; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2246 = 7'h45 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1222; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2247 = 7'h46 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1223; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2248 = 7'h47 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1224; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2249 = 7'h48 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1225; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2250 = 7'h49 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1226; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2251 = 7'h4a == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1227; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2252 = 7'h4b == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1228; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2253 = 7'h4c == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1229; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2254 = 7'h4d == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1230; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2255 = 7'h4e == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1231; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2256 = 7'h4f == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1232; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2257 = 7'h50 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1233; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2258 = 7'h51 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1234; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2259 = 7'h52 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1235; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2260 = 7'h53 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1236; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2261 = 7'h54 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1237; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2262 = 7'h55 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1238; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2263 = 7'h56 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1239; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2264 = 7'h57 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1240; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2265 = 7'h58 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1241; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2266 = 7'h59 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1242; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2267 = 7'h5a == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1243; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2268 = 7'h5b == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1244; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2269 = 7'h5c == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1245; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2270 = 7'h5d == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1246; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2271 = 7'h5e == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1247; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2272 = 7'h5f == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1248; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2273 = 7'h60 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1249; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2274 = 7'h61 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1250; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2275 = 7'h62 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1251; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2276 = 7'h63 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1252; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2277 = 7'h64 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1253; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2278 = 7'h65 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1254; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2279 = 7'h66 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1255; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2280 = 7'h67 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1256; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2281 = 7'h68 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1257; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2282 = 7'h69 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1258; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2283 = 7'h6a == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1259; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2284 = 7'h6b == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1260; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2285 = 7'h6c == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1261; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2286 = 7'h6d == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1262; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2287 = 7'h6e == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1263; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2288 = 7'h6f == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1264; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2289 = 7'h70 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1265; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2290 = 7'h71 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1266; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2291 = 7'h72 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1267; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2292 = 7'h73 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1268; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2293 = 7'h74 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1269; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2294 = 7'h75 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1270; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2295 = 7'h76 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1271; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2296 = 7'h77 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1272; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2297 = 7'h78 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1273; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2298 = 7'h79 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1274; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2299 = 7'h7a == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1275; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2300 = 7'h7b == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1276; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2301 = 7'h7c == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1277; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2302 = 7'h7d == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1278; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2303 = 7'h7e == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1279; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2304 = 7'h7f == rob_alloc_ids_1 ? _rob_payload_WIRE_3[31:16] : _GEN_1280; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2305 = 7'h0 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1281; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2306 = 7'h1 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1282; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2307 = 7'h2 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1283; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2308 = 7'h3 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1284; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2309 = 7'h4 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1285; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2310 = 7'h5 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1286; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2311 = 7'h6 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1287; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2312 = 7'h7 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1288; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2313 = 7'h8 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1289; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2314 = 7'h9 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1290; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2315 = 7'ha == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1291; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2316 = 7'hb == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1292; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2317 = 7'hc == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1293; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2318 = 7'hd == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1294; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2319 = 7'he == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1295; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2320 = 7'hf == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1296; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2321 = 7'h10 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1297; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2322 = 7'h11 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1298; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2323 = 7'h12 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1299; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2324 = 7'h13 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1300; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2325 = 7'h14 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1301; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2326 = 7'h15 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1302; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2327 = 7'h16 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1303; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2328 = 7'h17 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1304; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2329 = 7'h18 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1305; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2330 = 7'h19 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1306; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2331 = 7'h1a == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1307; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2332 = 7'h1b == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1308; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2333 = 7'h1c == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1309; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2334 = 7'h1d == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1310; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2335 = 7'h1e == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1311; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2336 = 7'h1f == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1312; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2337 = 7'h20 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1313; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2338 = 7'h21 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1314; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2339 = 7'h22 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1315; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2340 = 7'h23 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1316; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2341 = 7'h24 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1317; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2342 = 7'h25 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1318; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2343 = 7'h26 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1319; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2344 = 7'h27 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1320; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2345 = 7'h28 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1321; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2346 = 7'h29 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1322; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2347 = 7'h2a == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1323; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2348 = 7'h2b == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1324; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2349 = 7'h2c == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1325; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2350 = 7'h2d == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1326; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2351 = 7'h2e == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1327; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2352 = 7'h2f == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1328; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2353 = 7'h30 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1329; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2354 = 7'h31 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1330; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2355 = 7'h32 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1331; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2356 = 7'h33 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1332; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2357 = 7'h34 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1333; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2358 = 7'h35 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1334; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2359 = 7'h36 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1335; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2360 = 7'h37 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1336; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2361 = 7'h38 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1337; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2362 = 7'h39 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1338; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2363 = 7'h3a == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1339; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2364 = 7'h3b == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1340; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2365 = 7'h3c == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1341; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2366 = 7'h3d == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1342; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2367 = 7'h3e == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1343; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2368 = 7'h3f == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1344; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2369 = 7'h40 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1345; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2370 = 7'h41 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1346; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2371 = 7'h42 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1347; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2372 = 7'h43 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1348; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2373 = 7'h44 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1349; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2374 = 7'h45 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1350; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2375 = 7'h46 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1351; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2376 = 7'h47 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1352; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2377 = 7'h48 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1353; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2378 = 7'h49 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1354; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2379 = 7'h4a == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1355; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2380 = 7'h4b == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1356; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2381 = 7'h4c == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1357; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2382 = 7'h4d == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1358; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2383 = 7'h4e == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1359; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2384 = 7'h4f == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1360; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2385 = 7'h50 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1361; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2386 = 7'h51 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1362; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2387 = 7'h52 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1363; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2388 = 7'h53 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1364; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2389 = 7'h54 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1365; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2390 = 7'h55 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1366; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2391 = 7'h56 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1367; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2392 = 7'h57 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1368; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2393 = 7'h58 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1369; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2394 = 7'h59 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1370; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2395 = 7'h5a == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1371; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2396 = 7'h5b == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1372; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2397 = 7'h5c == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1373; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2398 = 7'h5d == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1374; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2399 = 7'h5e == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1375; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2400 = 7'h5f == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1376; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2401 = 7'h60 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1377; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2402 = 7'h61 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1378; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2403 = 7'h62 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1379; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2404 = 7'h63 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1380; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2405 = 7'h64 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1381; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2406 = 7'h65 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1382; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2407 = 7'h66 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1383; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2408 = 7'h67 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1384; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2409 = 7'h68 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1385; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2410 = 7'h69 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1386; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2411 = 7'h6a == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1387; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2412 = 7'h6b == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1388; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2413 = 7'h6c == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1389; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2414 = 7'h6d == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1390; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2415 = 7'h6e == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1391; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2416 = 7'h6f == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1392; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2417 = 7'h70 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1393; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2418 = 7'h71 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1394; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2419 = 7'h72 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1395; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2420 = 7'h73 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1396; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2421 = 7'h74 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1397; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2422 = 7'h75 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1398; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2423 = 7'h76 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1399; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2424 = 7'h77 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1400; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2425 = 7'h78 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1401; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2426 = 7'h79 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1402; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2427 = 7'h7a == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1403; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2428 = 7'h7b == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1404; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2429 = 7'h7c == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1405; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2430 = 7'h7d == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1406; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2431 = 7'h7e == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1407; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2432 = 7'h7f == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1408; // @[TestHarness.scala 179:{36,36}]
  wire [1:0] _rob_egress_id_T_37 = igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2433 = 7'h0 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1409; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2434 = 7'h1 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1410; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2435 = 7'h2 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1411; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2436 = 7'h3 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1412; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2437 = 7'h4 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1413; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2438 = 7'h5 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1414; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2439 = 7'h6 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1415; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2440 = 7'h7 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1416; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2441 = 7'h8 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1417; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2442 = 7'h9 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1418; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2443 = 7'ha == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1419; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2444 = 7'hb == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1420; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2445 = 7'hc == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1421; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2446 = 7'hd == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1422; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2447 = 7'he == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1423; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2448 = 7'hf == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1424; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2449 = 7'h10 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1425; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2450 = 7'h11 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1426; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2451 = 7'h12 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1427; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2452 = 7'h13 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1428; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2453 = 7'h14 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1429; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2454 = 7'h15 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1430; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2455 = 7'h16 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1431; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2456 = 7'h17 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1432; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2457 = 7'h18 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1433; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2458 = 7'h19 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1434; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2459 = 7'h1a == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1435; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2460 = 7'h1b == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1436; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2461 = 7'h1c == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1437; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2462 = 7'h1d == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1438; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2463 = 7'h1e == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1439; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2464 = 7'h1f == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1440; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2465 = 7'h20 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1441; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2466 = 7'h21 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1442; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2467 = 7'h22 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1443; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2468 = 7'h23 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1444; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2469 = 7'h24 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1445; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2470 = 7'h25 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1446; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2471 = 7'h26 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1447; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2472 = 7'h27 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1448; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2473 = 7'h28 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1449; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2474 = 7'h29 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1450; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2475 = 7'h2a == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1451; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2476 = 7'h2b == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1452; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2477 = 7'h2c == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1453; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2478 = 7'h2d == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1454; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2479 = 7'h2e == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1455; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2480 = 7'h2f == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1456; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2481 = 7'h30 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1457; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2482 = 7'h31 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1458; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2483 = 7'h32 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1459; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2484 = 7'h33 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1460; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2485 = 7'h34 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1461; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2486 = 7'h35 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1462; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2487 = 7'h36 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1463; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2488 = 7'h37 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1464; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2489 = 7'h38 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1465; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2490 = 7'h39 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1466; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2491 = 7'h3a == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1467; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2492 = 7'h3b == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1468; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2493 = 7'h3c == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1469; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2494 = 7'h3d == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1470; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2495 = 7'h3e == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1471; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2496 = 7'h3f == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1472; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2497 = 7'h40 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1473; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2498 = 7'h41 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1474; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2499 = 7'h42 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1475; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2500 = 7'h43 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1476; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2501 = 7'h44 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1477; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2502 = 7'h45 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1478; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2503 = 7'h46 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1479; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2504 = 7'h47 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1480; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2505 = 7'h48 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1481; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2506 = 7'h49 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1482; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2507 = 7'h4a == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1483; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2508 = 7'h4b == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1484; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2509 = 7'h4c == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1485; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2510 = 7'h4d == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1486; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2511 = 7'h4e == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1487; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2512 = 7'h4f == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1488; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2513 = 7'h50 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1489; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2514 = 7'h51 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1490; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2515 = 7'h52 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1491; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2516 = 7'h53 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1492; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2517 = 7'h54 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1493; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2518 = 7'h55 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1494; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2519 = 7'h56 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1495; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2520 = 7'h57 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1496; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2521 = 7'h58 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1497; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2522 = 7'h59 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1498; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2523 = 7'h5a == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1499; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2524 = 7'h5b == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1500; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2525 = 7'h5c == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1501; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2526 = 7'h5d == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1502; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2527 = 7'h5e == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1503; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2528 = 7'h5f == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1504; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2529 = 7'h60 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1505; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2530 = 7'h61 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1506; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2531 = 7'h62 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1507; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2532 = 7'h63 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1508; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2533 = 7'h64 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1509; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2534 = 7'h65 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1510; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2535 = 7'h66 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1511; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2536 = 7'h67 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1512; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2537 = 7'h68 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1513; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2538 = 7'h69 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1514; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2539 = 7'h6a == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1515; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2540 = 7'h6b == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1516; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2541 = 7'h6c == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1517; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2542 = 7'h6d == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1518; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2543 = 7'h6e == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1519; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2544 = 7'h6f == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1520; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2545 = 7'h70 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1521; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2546 = 7'h71 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1522; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2547 = 7'h72 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1523; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2548 = 7'h73 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1524; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2549 = 7'h74 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1525; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2550 = 7'h75 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1526; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2551 = 7'h76 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1527; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2552 = 7'h77 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1528; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2553 = 7'h78 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1529; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2554 = 7'h79 == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1530; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2555 = 7'h7a == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1531; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2556 = 7'h7b == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1532; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2557 = 7'h7c == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1533; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2558 = 7'h7d == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1534; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2559 = 7'h7e == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1535; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2560 = 7'h7f == rob_alloc_ids_1 ? _rob_egress_id_T_37 : _GEN_1536; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_2561 = 7'h0 == rob_alloc_ids_1 ? 2'h1 : _GEN_1537; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2562 = 7'h1 == rob_alloc_ids_1 ? 2'h1 : _GEN_1538; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2563 = 7'h2 == rob_alloc_ids_1 ? 2'h1 : _GEN_1539; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2564 = 7'h3 == rob_alloc_ids_1 ? 2'h1 : _GEN_1540; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2565 = 7'h4 == rob_alloc_ids_1 ? 2'h1 : _GEN_1541; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2566 = 7'h5 == rob_alloc_ids_1 ? 2'h1 : _GEN_1542; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2567 = 7'h6 == rob_alloc_ids_1 ? 2'h1 : _GEN_1543; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2568 = 7'h7 == rob_alloc_ids_1 ? 2'h1 : _GEN_1544; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2569 = 7'h8 == rob_alloc_ids_1 ? 2'h1 : _GEN_1545; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2570 = 7'h9 == rob_alloc_ids_1 ? 2'h1 : _GEN_1546; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2571 = 7'ha == rob_alloc_ids_1 ? 2'h1 : _GEN_1547; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2572 = 7'hb == rob_alloc_ids_1 ? 2'h1 : _GEN_1548; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2573 = 7'hc == rob_alloc_ids_1 ? 2'h1 : _GEN_1549; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2574 = 7'hd == rob_alloc_ids_1 ? 2'h1 : _GEN_1550; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2575 = 7'he == rob_alloc_ids_1 ? 2'h1 : _GEN_1551; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2576 = 7'hf == rob_alloc_ids_1 ? 2'h1 : _GEN_1552; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2577 = 7'h10 == rob_alloc_ids_1 ? 2'h1 : _GEN_1553; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2578 = 7'h11 == rob_alloc_ids_1 ? 2'h1 : _GEN_1554; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2579 = 7'h12 == rob_alloc_ids_1 ? 2'h1 : _GEN_1555; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2580 = 7'h13 == rob_alloc_ids_1 ? 2'h1 : _GEN_1556; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2581 = 7'h14 == rob_alloc_ids_1 ? 2'h1 : _GEN_1557; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2582 = 7'h15 == rob_alloc_ids_1 ? 2'h1 : _GEN_1558; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2583 = 7'h16 == rob_alloc_ids_1 ? 2'h1 : _GEN_1559; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2584 = 7'h17 == rob_alloc_ids_1 ? 2'h1 : _GEN_1560; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2585 = 7'h18 == rob_alloc_ids_1 ? 2'h1 : _GEN_1561; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2586 = 7'h19 == rob_alloc_ids_1 ? 2'h1 : _GEN_1562; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2587 = 7'h1a == rob_alloc_ids_1 ? 2'h1 : _GEN_1563; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2588 = 7'h1b == rob_alloc_ids_1 ? 2'h1 : _GEN_1564; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2589 = 7'h1c == rob_alloc_ids_1 ? 2'h1 : _GEN_1565; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2590 = 7'h1d == rob_alloc_ids_1 ? 2'h1 : _GEN_1566; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2591 = 7'h1e == rob_alloc_ids_1 ? 2'h1 : _GEN_1567; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2592 = 7'h1f == rob_alloc_ids_1 ? 2'h1 : _GEN_1568; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2593 = 7'h20 == rob_alloc_ids_1 ? 2'h1 : _GEN_1569; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2594 = 7'h21 == rob_alloc_ids_1 ? 2'h1 : _GEN_1570; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2595 = 7'h22 == rob_alloc_ids_1 ? 2'h1 : _GEN_1571; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2596 = 7'h23 == rob_alloc_ids_1 ? 2'h1 : _GEN_1572; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2597 = 7'h24 == rob_alloc_ids_1 ? 2'h1 : _GEN_1573; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2598 = 7'h25 == rob_alloc_ids_1 ? 2'h1 : _GEN_1574; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2599 = 7'h26 == rob_alloc_ids_1 ? 2'h1 : _GEN_1575; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2600 = 7'h27 == rob_alloc_ids_1 ? 2'h1 : _GEN_1576; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2601 = 7'h28 == rob_alloc_ids_1 ? 2'h1 : _GEN_1577; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2602 = 7'h29 == rob_alloc_ids_1 ? 2'h1 : _GEN_1578; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2603 = 7'h2a == rob_alloc_ids_1 ? 2'h1 : _GEN_1579; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2604 = 7'h2b == rob_alloc_ids_1 ? 2'h1 : _GEN_1580; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2605 = 7'h2c == rob_alloc_ids_1 ? 2'h1 : _GEN_1581; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2606 = 7'h2d == rob_alloc_ids_1 ? 2'h1 : _GEN_1582; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2607 = 7'h2e == rob_alloc_ids_1 ? 2'h1 : _GEN_1583; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2608 = 7'h2f == rob_alloc_ids_1 ? 2'h1 : _GEN_1584; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2609 = 7'h30 == rob_alloc_ids_1 ? 2'h1 : _GEN_1585; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2610 = 7'h31 == rob_alloc_ids_1 ? 2'h1 : _GEN_1586; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2611 = 7'h32 == rob_alloc_ids_1 ? 2'h1 : _GEN_1587; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2612 = 7'h33 == rob_alloc_ids_1 ? 2'h1 : _GEN_1588; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2613 = 7'h34 == rob_alloc_ids_1 ? 2'h1 : _GEN_1589; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2614 = 7'h35 == rob_alloc_ids_1 ? 2'h1 : _GEN_1590; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2615 = 7'h36 == rob_alloc_ids_1 ? 2'h1 : _GEN_1591; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2616 = 7'h37 == rob_alloc_ids_1 ? 2'h1 : _GEN_1592; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2617 = 7'h38 == rob_alloc_ids_1 ? 2'h1 : _GEN_1593; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2618 = 7'h39 == rob_alloc_ids_1 ? 2'h1 : _GEN_1594; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2619 = 7'h3a == rob_alloc_ids_1 ? 2'h1 : _GEN_1595; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2620 = 7'h3b == rob_alloc_ids_1 ? 2'h1 : _GEN_1596; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2621 = 7'h3c == rob_alloc_ids_1 ? 2'h1 : _GEN_1597; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2622 = 7'h3d == rob_alloc_ids_1 ? 2'h1 : _GEN_1598; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2623 = 7'h3e == rob_alloc_ids_1 ? 2'h1 : _GEN_1599; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2624 = 7'h3f == rob_alloc_ids_1 ? 2'h1 : _GEN_1600; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2625 = 7'h40 == rob_alloc_ids_1 ? 2'h1 : _GEN_1601; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2626 = 7'h41 == rob_alloc_ids_1 ? 2'h1 : _GEN_1602; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2627 = 7'h42 == rob_alloc_ids_1 ? 2'h1 : _GEN_1603; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2628 = 7'h43 == rob_alloc_ids_1 ? 2'h1 : _GEN_1604; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2629 = 7'h44 == rob_alloc_ids_1 ? 2'h1 : _GEN_1605; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2630 = 7'h45 == rob_alloc_ids_1 ? 2'h1 : _GEN_1606; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2631 = 7'h46 == rob_alloc_ids_1 ? 2'h1 : _GEN_1607; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2632 = 7'h47 == rob_alloc_ids_1 ? 2'h1 : _GEN_1608; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2633 = 7'h48 == rob_alloc_ids_1 ? 2'h1 : _GEN_1609; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2634 = 7'h49 == rob_alloc_ids_1 ? 2'h1 : _GEN_1610; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2635 = 7'h4a == rob_alloc_ids_1 ? 2'h1 : _GEN_1611; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2636 = 7'h4b == rob_alloc_ids_1 ? 2'h1 : _GEN_1612; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2637 = 7'h4c == rob_alloc_ids_1 ? 2'h1 : _GEN_1613; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2638 = 7'h4d == rob_alloc_ids_1 ? 2'h1 : _GEN_1614; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2639 = 7'h4e == rob_alloc_ids_1 ? 2'h1 : _GEN_1615; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2640 = 7'h4f == rob_alloc_ids_1 ? 2'h1 : _GEN_1616; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2641 = 7'h50 == rob_alloc_ids_1 ? 2'h1 : _GEN_1617; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2642 = 7'h51 == rob_alloc_ids_1 ? 2'h1 : _GEN_1618; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2643 = 7'h52 == rob_alloc_ids_1 ? 2'h1 : _GEN_1619; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2644 = 7'h53 == rob_alloc_ids_1 ? 2'h1 : _GEN_1620; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2645 = 7'h54 == rob_alloc_ids_1 ? 2'h1 : _GEN_1621; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2646 = 7'h55 == rob_alloc_ids_1 ? 2'h1 : _GEN_1622; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2647 = 7'h56 == rob_alloc_ids_1 ? 2'h1 : _GEN_1623; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2648 = 7'h57 == rob_alloc_ids_1 ? 2'h1 : _GEN_1624; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2649 = 7'h58 == rob_alloc_ids_1 ? 2'h1 : _GEN_1625; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2650 = 7'h59 == rob_alloc_ids_1 ? 2'h1 : _GEN_1626; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2651 = 7'h5a == rob_alloc_ids_1 ? 2'h1 : _GEN_1627; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2652 = 7'h5b == rob_alloc_ids_1 ? 2'h1 : _GEN_1628; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2653 = 7'h5c == rob_alloc_ids_1 ? 2'h1 : _GEN_1629; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2654 = 7'h5d == rob_alloc_ids_1 ? 2'h1 : _GEN_1630; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2655 = 7'h5e == rob_alloc_ids_1 ? 2'h1 : _GEN_1631; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2656 = 7'h5f == rob_alloc_ids_1 ? 2'h1 : _GEN_1632; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2657 = 7'h60 == rob_alloc_ids_1 ? 2'h1 : _GEN_1633; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2658 = 7'h61 == rob_alloc_ids_1 ? 2'h1 : _GEN_1634; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2659 = 7'h62 == rob_alloc_ids_1 ? 2'h1 : _GEN_1635; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2660 = 7'h63 == rob_alloc_ids_1 ? 2'h1 : _GEN_1636; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2661 = 7'h64 == rob_alloc_ids_1 ? 2'h1 : _GEN_1637; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2662 = 7'h65 == rob_alloc_ids_1 ? 2'h1 : _GEN_1638; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2663 = 7'h66 == rob_alloc_ids_1 ? 2'h1 : _GEN_1639; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2664 = 7'h67 == rob_alloc_ids_1 ? 2'h1 : _GEN_1640; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2665 = 7'h68 == rob_alloc_ids_1 ? 2'h1 : _GEN_1641; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2666 = 7'h69 == rob_alloc_ids_1 ? 2'h1 : _GEN_1642; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2667 = 7'h6a == rob_alloc_ids_1 ? 2'h1 : _GEN_1643; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2668 = 7'h6b == rob_alloc_ids_1 ? 2'h1 : _GEN_1644; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2669 = 7'h6c == rob_alloc_ids_1 ? 2'h1 : _GEN_1645; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2670 = 7'h6d == rob_alloc_ids_1 ? 2'h1 : _GEN_1646; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2671 = 7'h6e == rob_alloc_ids_1 ? 2'h1 : _GEN_1647; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2672 = 7'h6f == rob_alloc_ids_1 ? 2'h1 : _GEN_1648; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2673 = 7'h70 == rob_alloc_ids_1 ? 2'h1 : _GEN_1649; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2674 = 7'h71 == rob_alloc_ids_1 ? 2'h1 : _GEN_1650; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2675 = 7'h72 == rob_alloc_ids_1 ? 2'h1 : _GEN_1651; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2676 = 7'h73 == rob_alloc_ids_1 ? 2'h1 : _GEN_1652; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2677 = 7'h74 == rob_alloc_ids_1 ? 2'h1 : _GEN_1653; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2678 = 7'h75 == rob_alloc_ids_1 ? 2'h1 : _GEN_1654; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2679 = 7'h76 == rob_alloc_ids_1 ? 2'h1 : _GEN_1655; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2680 = 7'h77 == rob_alloc_ids_1 ? 2'h1 : _GEN_1656; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2681 = 7'h78 == rob_alloc_ids_1 ? 2'h1 : _GEN_1657; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2682 = 7'h79 == rob_alloc_ids_1 ? 2'h1 : _GEN_1658; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2683 = 7'h7a == rob_alloc_ids_1 ? 2'h1 : _GEN_1659; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2684 = 7'h7b == rob_alloc_ids_1 ? 2'h1 : _GEN_1660; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2685 = 7'h7c == rob_alloc_ids_1 ? 2'h1 : _GEN_1661; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2686 = 7'h7d == rob_alloc_ids_1 ? 2'h1 : _GEN_1662; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2687 = 7'h7e == rob_alloc_ids_1 ? 2'h1 : _GEN_1663; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_2688 = 7'h7f == rob_alloc_ids_1 ? 2'h1 : _GEN_1664; // @[TestHarness.scala 181:{36,36}]
  wire [3:0] _rob_n_flits_T_41 = igen_1_io_n_flits; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2689 = 7'h0 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1665; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2690 = 7'h1 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1666; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2691 = 7'h2 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1667; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2692 = 7'h3 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1668; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2693 = 7'h4 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1669; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2694 = 7'h5 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1670; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2695 = 7'h6 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1671; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2696 = 7'h7 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1672; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2697 = 7'h8 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1673; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2698 = 7'h9 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1674; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2699 = 7'ha == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1675; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2700 = 7'hb == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1676; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2701 = 7'hc == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1677; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2702 = 7'hd == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1678; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2703 = 7'he == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1679; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2704 = 7'hf == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1680; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2705 = 7'h10 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1681; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2706 = 7'h11 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1682; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2707 = 7'h12 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1683; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2708 = 7'h13 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1684; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2709 = 7'h14 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1685; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2710 = 7'h15 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1686; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2711 = 7'h16 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1687; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2712 = 7'h17 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1688; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2713 = 7'h18 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1689; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2714 = 7'h19 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1690; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2715 = 7'h1a == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1691; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2716 = 7'h1b == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1692; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2717 = 7'h1c == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1693; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2718 = 7'h1d == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1694; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2719 = 7'h1e == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1695; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2720 = 7'h1f == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1696; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2721 = 7'h20 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1697; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2722 = 7'h21 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1698; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2723 = 7'h22 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1699; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2724 = 7'h23 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1700; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2725 = 7'h24 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1701; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2726 = 7'h25 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1702; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2727 = 7'h26 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1703; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2728 = 7'h27 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1704; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2729 = 7'h28 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1705; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2730 = 7'h29 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1706; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2731 = 7'h2a == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1707; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2732 = 7'h2b == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1708; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2733 = 7'h2c == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1709; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2734 = 7'h2d == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1710; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2735 = 7'h2e == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1711; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2736 = 7'h2f == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1712; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2737 = 7'h30 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1713; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2738 = 7'h31 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1714; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2739 = 7'h32 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1715; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2740 = 7'h33 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1716; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2741 = 7'h34 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1717; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2742 = 7'h35 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1718; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2743 = 7'h36 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1719; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2744 = 7'h37 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1720; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2745 = 7'h38 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1721; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2746 = 7'h39 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1722; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2747 = 7'h3a == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1723; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2748 = 7'h3b == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1724; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2749 = 7'h3c == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1725; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2750 = 7'h3d == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1726; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2751 = 7'h3e == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1727; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2752 = 7'h3f == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1728; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2753 = 7'h40 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1729; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2754 = 7'h41 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1730; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2755 = 7'h42 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1731; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2756 = 7'h43 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1732; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2757 = 7'h44 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1733; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2758 = 7'h45 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1734; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2759 = 7'h46 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1735; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2760 = 7'h47 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1736; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2761 = 7'h48 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1737; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2762 = 7'h49 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1738; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2763 = 7'h4a == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1739; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2764 = 7'h4b == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1740; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2765 = 7'h4c == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1741; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2766 = 7'h4d == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1742; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2767 = 7'h4e == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1743; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2768 = 7'h4f == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1744; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2769 = 7'h50 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1745; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2770 = 7'h51 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1746; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2771 = 7'h52 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1747; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2772 = 7'h53 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1748; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2773 = 7'h54 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1749; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2774 = 7'h55 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1750; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2775 = 7'h56 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1751; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2776 = 7'h57 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1752; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2777 = 7'h58 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1753; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2778 = 7'h59 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1754; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2779 = 7'h5a == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1755; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2780 = 7'h5b == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1756; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2781 = 7'h5c == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1757; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2782 = 7'h5d == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1758; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2783 = 7'h5e == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1759; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2784 = 7'h5f == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1760; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2785 = 7'h60 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1761; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2786 = 7'h61 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1762; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2787 = 7'h62 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1763; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2788 = 7'h63 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1764; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2789 = 7'h64 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1765; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2790 = 7'h65 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1766; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2791 = 7'h66 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1767; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2792 = 7'h67 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1768; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2793 = 7'h68 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1769; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2794 = 7'h69 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1770; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2795 = 7'h6a == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1771; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2796 = 7'h6b == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1772; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2797 = 7'h6c == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1773; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2798 = 7'h6d == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1774; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2799 = 7'h6e == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1775; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2800 = 7'h6f == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1776; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2801 = 7'h70 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1777; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2802 = 7'h71 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1778; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2803 = 7'h72 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1779; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2804 = 7'h73 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1780; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2805 = 7'h74 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1781; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2806 = 7'h75 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1782; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2807 = 7'h76 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1783; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2808 = 7'h77 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1784; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2809 = 7'h78 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1785; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2810 = 7'h79 == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1786; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2811 = 7'h7a == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1787; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2812 = 7'h7b == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1788; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2813 = 7'h7c == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1789; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2814 = 7'h7d == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1790; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2815 = 7'h7e == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1791; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2816 = 7'h7f == rob_alloc_ids_1 ? _rob_n_flits_T_41 : _GEN_1792; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2817 = 7'h0 == rob_alloc_ids_1 ? 4'h0 : _GEN_1793; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2818 = 7'h1 == rob_alloc_ids_1 ? 4'h0 : _GEN_1794; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2819 = 7'h2 == rob_alloc_ids_1 ? 4'h0 : _GEN_1795; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2820 = 7'h3 == rob_alloc_ids_1 ? 4'h0 : _GEN_1796; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2821 = 7'h4 == rob_alloc_ids_1 ? 4'h0 : _GEN_1797; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2822 = 7'h5 == rob_alloc_ids_1 ? 4'h0 : _GEN_1798; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2823 = 7'h6 == rob_alloc_ids_1 ? 4'h0 : _GEN_1799; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2824 = 7'h7 == rob_alloc_ids_1 ? 4'h0 : _GEN_1800; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2825 = 7'h8 == rob_alloc_ids_1 ? 4'h0 : _GEN_1801; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2826 = 7'h9 == rob_alloc_ids_1 ? 4'h0 : _GEN_1802; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2827 = 7'ha == rob_alloc_ids_1 ? 4'h0 : _GEN_1803; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2828 = 7'hb == rob_alloc_ids_1 ? 4'h0 : _GEN_1804; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2829 = 7'hc == rob_alloc_ids_1 ? 4'h0 : _GEN_1805; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2830 = 7'hd == rob_alloc_ids_1 ? 4'h0 : _GEN_1806; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2831 = 7'he == rob_alloc_ids_1 ? 4'h0 : _GEN_1807; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2832 = 7'hf == rob_alloc_ids_1 ? 4'h0 : _GEN_1808; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2833 = 7'h10 == rob_alloc_ids_1 ? 4'h0 : _GEN_1809; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2834 = 7'h11 == rob_alloc_ids_1 ? 4'h0 : _GEN_1810; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2835 = 7'h12 == rob_alloc_ids_1 ? 4'h0 : _GEN_1811; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2836 = 7'h13 == rob_alloc_ids_1 ? 4'h0 : _GEN_1812; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2837 = 7'h14 == rob_alloc_ids_1 ? 4'h0 : _GEN_1813; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2838 = 7'h15 == rob_alloc_ids_1 ? 4'h0 : _GEN_1814; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2839 = 7'h16 == rob_alloc_ids_1 ? 4'h0 : _GEN_1815; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2840 = 7'h17 == rob_alloc_ids_1 ? 4'h0 : _GEN_1816; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2841 = 7'h18 == rob_alloc_ids_1 ? 4'h0 : _GEN_1817; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2842 = 7'h19 == rob_alloc_ids_1 ? 4'h0 : _GEN_1818; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2843 = 7'h1a == rob_alloc_ids_1 ? 4'h0 : _GEN_1819; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2844 = 7'h1b == rob_alloc_ids_1 ? 4'h0 : _GEN_1820; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2845 = 7'h1c == rob_alloc_ids_1 ? 4'h0 : _GEN_1821; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2846 = 7'h1d == rob_alloc_ids_1 ? 4'h0 : _GEN_1822; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2847 = 7'h1e == rob_alloc_ids_1 ? 4'h0 : _GEN_1823; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2848 = 7'h1f == rob_alloc_ids_1 ? 4'h0 : _GEN_1824; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2849 = 7'h20 == rob_alloc_ids_1 ? 4'h0 : _GEN_1825; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2850 = 7'h21 == rob_alloc_ids_1 ? 4'h0 : _GEN_1826; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2851 = 7'h22 == rob_alloc_ids_1 ? 4'h0 : _GEN_1827; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2852 = 7'h23 == rob_alloc_ids_1 ? 4'h0 : _GEN_1828; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2853 = 7'h24 == rob_alloc_ids_1 ? 4'h0 : _GEN_1829; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2854 = 7'h25 == rob_alloc_ids_1 ? 4'h0 : _GEN_1830; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2855 = 7'h26 == rob_alloc_ids_1 ? 4'h0 : _GEN_1831; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2856 = 7'h27 == rob_alloc_ids_1 ? 4'h0 : _GEN_1832; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2857 = 7'h28 == rob_alloc_ids_1 ? 4'h0 : _GEN_1833; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2858 = 7'h29 == rob_alloc_ids_1 ? 4'h0 : _GEN_1834; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2859 = 7'h2a == rob_alloc_ids_1 ? 4'h0 : _GEN_1835; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2860 = 7'h2b == rob_alloc_ids_1 ? 4'h0 : _GEN_1836; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2861 = 7'h2c == rob_alloc_ids_1 ? 4'h0 : _GEN_1837; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2862 = 7'h2d == rob_alloc_ids_1 ? 4'h0 : _GEN_1838; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2863 = 7'h2e == rob_alloc_ids_1 ? 4'h0 : _GEN_1839; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2864 = 7'h2f == rob_alloc_ids_1 ? 4'h0 : _GEN_1840; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2865 = 7'h30 == rob_alloc_ids_1 ? 4'h0 : _GEN_1841; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2866 = 7'h31 == rob_alloc_ids_1 ? 4'h0 : _GEN_1842; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2867 = 7'h32 == rob_alloc_ids_1 ? 4'h0 : _GEN_1843; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2868 = 7'h33 == rob_alloc_ids_1 ? 4'h0 : _GEN_1844; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2869 = 7'h34 == rob_alloc_ids_1 ? 4'h0 : _GEN_1845; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2870 = 7'h35 == rob_alloc_ids_1 ? 4'h0 : _GEN_1846; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2871 = 7'h36 == rob_alloc_ids_1 ? 4'h0 : _GEN_1847; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2872 = 7'h37 == rob_alloc_ids_1 ? 4'h0 : _GEN_1848; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2873 = 7'h38 == rob_alloc_ids_1 ? 4'h0 : _GEN_1849; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2874 = 7'h39 == rob_alloc_ids_1 ? 4'h0 : _GEN_1850; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2875 = 7'h3a == rob_alloc_ids_1 ? 4'h0 : _GEN_1851; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2876 = 7'h3b == rob_alloc_ids_1 ? 4'h0 : _GEN_1852; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2877 = 7'h3c == rob_alloc_ids_1 ? 4'h0 : _GEN_1853; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2878 = 7'h3d == rob_alloc_ids_1 ? 4'h0 : _GEN_1854; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2879 = 7'h3e == rob_alloc_ids_1 ? 4'h0 : _GEN_1855; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2880 = 7'h3f == rob_alloc_ids_1 ? 4'h0 : _GEN_1856; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2881 = 7'h40 == rob_alloc_ids_1 ? 4'h0 : _GEN_1857; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2882 = 7'h41 == rob_alloc_ids_1 ? 4'h0 : _GEN_1858; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2883 = 7'h42 == rob_alloc_ids_1 ? 4'h0 : _GEN_1859; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2884 = 7'h43 == rob_alloc_ids_1 ? 4'h0 : _GEN_1860; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2885 = 7'h44 == rob_alloc_ids_1 ? 4'h0 : _GEN_1861; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2886 = 7'h45 == rob_alloc_ids_1 ? 4'h0 : _GEN_1862; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2887 = 7'h46 == rob_alloc_ids_1 ? 4'h0 : _GEN_1863; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2888 = 7'h47 == rob_alloc_ids_1 ? 4'h0 : _GEN_1864; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2889 = 7'h48 == rob_alloc_ids_1 ? 4'h0 : _GEN_1865; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2890 = 7'h49 == rob_alloc_ids_1 ? 4'h0 : _GEN_1866; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2891 = 7'h4a == rob_alloc_ids_1 ? 4'h0 : _GEN_1867; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2892 = 7'h4b == rob_alloc_ids_1 ? 4'h0 : _GEN_1868; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2893 = 7'h4c == rob_alloc_ids_1 ? 4'h0 : _GEN_1869; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2894 = 7'h4d == rob_alloc_ids_1 ? 4'h0 : _GEN_1870; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2895 = 7'h4e == rob_alloc_ids_1 ? 4'h0 : _GEN_1871; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2896 = 7'h4f == rob_alloc_ids_1 ? 4'h0 : _GEN_1872; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2897 = 7'h50 == rob_alloc_ids_1 ? 4'h0 : _GEN_1873; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2898 = 7'h51 == rob_alloc_ids_1 ? 4'h0 : _GEN_1874; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2899 = 7'h52 == rob_alloc_ids_1 ? 4'h0 : _GEN_1875; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2900 = 7'h53 == rob_alloc_ids_1 ? 4'h0 : _GEN_1876; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2901 = 7'h54 == rob_alloc_ids_1 ? 4'h0 : _GEN_1877; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2902 = 7'h55 == rob_alloc_ids_1 ? 4'h0 : _GEN_1878; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2903 = 7'h56 == rob_alloc_ids_1 ? 4'h0 : _GEN_1879; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2904 = 7'h57 == rob_alloc_ids_1 ? 4'h0 : _GEN_1880; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2905 = 7'h58 == rob_alloc_ids_1 ? 4'h0 : _GEN_1881; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2906 = 7'h59 == rob_alloc_ids_1 ? 4'h0 : _GEN_1882; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2907 = 7'h5a == rob_alloc_ids_1 ? 4'h0 : _GEN_1883; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2908 = 7'h5b == rob_alloc_ids_1 ? 4'h0 : _GEN_1884; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2909 = 7'h5c == rob_alloc_ids_1 ? 4'h0 : _GEN_1885; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2910 = 7'h5d == rob_alloc_ids_1 ? 4'h0 : _GEN_1886; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2911 = 7'h5e == rob_alloc_ids_1 ? 4'h0 : _GEN_1887; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2912 = 7'h5f == rob_alloc_ids_1 ? 4'h0 : _GEN_1888; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2913 = 7'h60 == rob_alloc_ids_1 ? 4'h0 : _GEN_1889; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2914 = 7'h61 == rob_alloc_ids_1 ? 4'h0 : _GEN_1890; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2915 = 7'h62 == rob_alloc_ids_1 ? 4'h0 : _GEN_1891; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2916 = 7'h63 == rob_alloc_ids_1 ? 4'h0 : _GEN_1892; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2917 = 7'h64 == rob_alloc_ids_1 ? 4'h0 : _GEN_1893; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2918 = 7'h65 == rob_alloc_ids_1 ? 4'h0 : _GEN_1894; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2919 = 7'h66 == rob_alloc_ids_1 ? 4'h0 : _GEN_1895; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2920 = 7'h67 == rob_alloc_ids_1 ? 4'h0 : _GEN_1896; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2921 = 7'h68 == rob_alloc_ids_1 ? 4'h0 : _GEN_1897; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2922 = 7'h69 == rob_alloc_ids_1 ? 4'h0 : _GEN_1898; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2923 = 7'h6a == rob_alloc_ids_1 ? 4'h0 : _GEN_1899; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2924 = 7'h6b == rob_alloc_ids_1 ? 4'h0 : _GEN_1900; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2925 = 7'h6c == rob_alloc_ids_1 ? 4'h0 : _GEN_1901; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2926 = 7'h6d == rob_alloc_ids_1 ? 4'h0 : _GEN_1902; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2927 = 7'h6e == rob_alloc_ids_1 ? 4'h0 : _GEN_1903; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2928 = 7'h6f == rob_alloc_ids_1 ? 4'h0 : _GEN_1904; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2929 = 7'h70 == rob_alloc_ids_1 ? 4'h0 : _GEN_1905; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2930 = 7'h71 == rob_alloc_ids_1 ? 4'h0 : _GEN_1906; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2931 = 7'h72 == rob_alloc_ids_1 ? 4'h0 : _GEN_1907; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2932 = 7'h73 == rob_alloc_ids_1 ? 4'h0 : _GEN_1908; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2933 = 7'h74 == rob_alloc_ids_1 ? 4'h0 : _GEN_1909; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2934 = 7'h75 == rob_alloc_ids_1 ? 4'h0 : _GEN_1910; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2935 = 7'h76 == rob_alloc_ids_1 ? 4'h0 : _GEN_1911; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2936 = 7'h77 == rob_alloc_ids_1 ? 4'h0 : _GEN_1912; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2937 = 7'h78 == rob_alloc_ids_1 ? 4'h0 : _GEN_1913; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2938 = 7'h79 == rob_alloc_ids_1 ? 4'h0 : _GEN_1914; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2939 = 7'h7a == rob_alloc_ids_1 ? 4'h0 : _GEN_1915; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2940 = 7'h7b == rob_alloc_ids_1 ? 4'h0 : _GEN_1916; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2941 = 7'h7c == rob_alloc_ids_1 ? 4'h0 : _GEN_1917; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2942 = 7'h7d == rob_alloc_ids_1 ? 4'h0 : _GEN_1918; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2943 = 7'h7e == rob_alloc_ids_1 ? 4'h0 : _GEN_1919; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2944 = 7'h7f == rob_alloc_ids_1 ? 4'h0 : _GEN_1920; // @[TestHarness.scala 183:{36,36}]
  wire [63:0] _GEN_2945 = 7'h0 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1921; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2946 = 7'h1 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1922; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2947 = 7'h2 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1923; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2948 = 7'h3 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1924; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2949 = 7'h4 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1925; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2950 = 7'h5 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1926; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2951 = 7'h6 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1927; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2952 = 7'h7 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1928; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2953 = 7'h8 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1929; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2954 = 7'h9 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1930; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2955 = 7'ha == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1931; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2956 = 7'hb == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1932; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2957 = 7'hc == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1933; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2958 = 7'hd == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1934; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2959 = 7'he == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1935; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2960 = 7'hf == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1936; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2961 = 7'h10 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1937; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2962 = 7'h11 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1938; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2963 = 7'h12 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1939; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2964 = 7'h13 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1940; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2965 = 7'h14 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1941; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2966 = 7'h15 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1942; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2967 = 7'h16 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1943; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2968 = 7'h17 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1944; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2969 = 7'h18 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1945; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2970 = 7'h19 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1946; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2971 = 7'h1a == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1947; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2972 = 7'h1b == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1948; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2973 = 7'h1c == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1949; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2974 = 7'h1d == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1950; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2975 = 7'h1e == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1951; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2976 = 7'h1f == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1952; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2977 = 7'h20 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1953; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2978 = 7'h21 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1954; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2979 = 7'h22 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1955; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2980 = 7'h23 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1956; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2981 = 7'h24 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1957; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2982 = 7'h25 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1958; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2983 = 7'h26 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1959; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2984 = 7'h27 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1960; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2985 = 7'h28 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1961; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2986 = 7'h29 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1962; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2987 = 7'h2a == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1963; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2988 = 7'h2b == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1964; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2989 = 7'h2c == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1965; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2990 = 7'h2d == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1966; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2991 = 7'h2e == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1967; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2992 = 7'h2f == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1968; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2993 = 7'h30 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1969; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2994 = 7'h31 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1970; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2995 = 7'h32 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1971; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2996 = 7'h33 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1972; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2997 = 7'h34 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1973; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2998 = 7'h35 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1974; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_2999 = 7'h36 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1975; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3000 = 7'h37 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1976; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3001 = 7'h38 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1977; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3002 = 7'h39 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1978; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3003 = 7'h3a == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1979; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3004 = 7'h3b == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1980; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3005 = 7'h3c == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1981; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3006 = 7'h3d == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1982; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3007 = 7'h3e == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1983; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3008 = 7'h3f == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1984; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3009 = 7'h40 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1985; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3010 = 7'h41 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1986; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3011 = 7'h42 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1987; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3012 = 7'h43 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1988; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3013 = 7'h44 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1989; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3014 = 7'h45 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1990; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3015 = 7'h46 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1991; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3016 = 7'h47 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1992; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3017 = 7'h48 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1993; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3018 = 7'h49 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1994; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3019 = 7'h4a == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1995; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3020 = 7'h4b == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1996; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3021 = 7'h4c == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1997; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3022 = 7'h4d == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1998; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3023 = 7'h4e == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_1999; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3024 = 7'h4f == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2000; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3025 = 7'h50 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2001; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3026 = 7'h51 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2002; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3027 = 7'h52 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2003; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3028 = 7'h53 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2004; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3029 = 7'h54 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2005; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3030 = 7'h55 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2006; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3031 = 7'h56 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2007; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3032 = 7'h57 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2008; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3033 = 7'h58 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2009; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3034 = 7'h59 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2010; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3035 = 7'h5a == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2011; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3036 = 7'h5b == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2012; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3037 = 7'h5c == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2013; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3038 = 7'h5d == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2014; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3039 = 7'h5e == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2015; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3040 = 7'h5f == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2016; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3041 = 7'h60 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2017; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3042 = 7'h61 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2018; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3043 = 7'h62 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2019; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3044 = 7'h63 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2020; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3045 = 7'h64 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2021; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3046 = 7'h65 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2022; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3047 = 7'h66 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2023; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3048 = 7'h67 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2024; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3049 = 7'h68 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2025; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3050 = 7'h69 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2026; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3051 = 7'h6a == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2027; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3052 = 7'h6b == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2028; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3053 = 7'h6c == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2029; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3054 = 7'h6d == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2030; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3055 = 7'h6e == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2031; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3056 = 7'h6f == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2032; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3057 = 7'h70 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2033; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3058 = 7'h71 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2034; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3059 = 7'h72 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2035; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3060 = 7'h73 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2036; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3061 = 7'h74 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2037; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3062 = 7'h75 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2038; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3063 = 7'h76 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2039; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3064 = 7'h77 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2040; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3065 = 7'h78 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2041; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3066 = 7'h79 == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2042; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3067 = 7'h7a == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2043; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3068 = 7'h7b == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2044; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3069 = 7'h7c == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2045; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3070 = 7'h7d == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2046; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3071 = 7'h7e == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2047; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_3072 = 7'h7f == rob_alloc_ids_1 ? _rob_tscs_T_31 : _GEN_2048; // @[TestHarness.scala 184:{36,36}]
  wire [31:0] _GEN_3073 = igen_1_io_fire ? _GEN_2049 : _GEN_1025; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3074 = igen_1_io_fire ? _GEN_2050 : _GEN_1026; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3075 = igen_1_io_fire ? _GEN_2051 : _GEN_1027; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3076 = igen_1_io_fire ? _GEN_2052 : _GEN_1028; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3077 = igen_1_io_fire ? _GEN_2053 : _GEN_1029; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3078 = igen_1_io_fire ? _GEN_2054 : _GEN_1030; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3079 = igen_1_io_fire ? _GEN_2055 : _GEN_1031; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3080 = igen_1_io_fire ? _GEN_2056 : _GEN_1032; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3081 = igen_1_io_fire ? _GEN_2057 : _GEN_1033; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3082 = igen_1_io_fire ? _GEN_2058 : _GEN_1034; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3083 = igen_1_io_fire ? _GEN_2059 : _GEN_1035; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3084 = igen_1_io_fire ? _GEN_2060 : _GEN_1036; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3085 = igen_1_io_fire ? _GEN_2061 : _GEN_1037; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3086 = igen_1_io_fire ? _GEN_2062 : _GEN_1038; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3087 = igen_1_io_fire ? _GEN_2063 : _GEN_1039; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3088 = igen_1_io_fire ? _GEN_2064 : _GEN_1040; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3089 = igen_1_io_fire ? _GEN_2065 : _GEN_1041; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3090 = igen_1_io_fire ? _GEN_2066 : _GEN_1042; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3091 = igen_1_io_fire ? _GEN_2067 : _GEN_1043; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3092 = igen_1_io_fire ? _GEN_2068 : _GEN_1044; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3093 = igen_1_io_fire ? _GEN_2069 : _GEN_1045; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3094 = igen_1_io_fire ? _GEN_2070 : _GEN_1046; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3095 = igen_1_io_fire ? _GEN_2071 : _GEN_1047; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3096 = igen_1_io_fire ? _GEN_2072 : _GEN_1048; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3097 = igen_1_io_fire ? _GEN_2073 : _GEN_1049; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3098 = igen_1_io_fire ? _GEN_2074 : _GEN_1050; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3099 = igen_1_io_fire ? _GEN_2075 : _GEN_1051; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3100 = igen_1_io_fire ? _GEN_2076 : _GEN_1052; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3101 = igen_1_io_fire ? _GEN_2077 : _GEN_1053; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3102 = igen_1_io_fire ? _GEN_2078 : _GEN_1054; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3103 = igen_1_io_fire ? _GEN_2079 : _GEN_1055; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3104 = igen_1_io_fire ? _GEN_2080 : _GEN_1056; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3105 = igen_1_io_fire ? _GEN_2081 : _GEN_1057; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3106 = igen_1_io_fire ? _GEN_2082 : _GEN_1058; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3107 = igen_1_io_fire ? _GEN_2083 : _GEN_1059; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3108 = igen_1_io_fire ? _GEN_2084 : _GEN_1060; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3109 = igen_1_io_fire ? _GEN_2085 : _GEN_1061; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3110 = igen_1_io_fire ? _GEN_2086 : _GEN_1062; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3111 = igen_1_io_fire ? _GEN_2087 : _GEN_1063; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3112 = igen_1_io_fire ? _GEN_2088 : _GEN_1064; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3113 = igen_1_io_fire ? _GEN_2089 : _GEN_1065; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3114 = igen_1_io_fire ? _GEN_2090 : _GEN_1066; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3115 = igen_1_io_fire ? _GEN_2091 : _GEN_1067; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3116 = igen_1_io_fire ? _GEN_2092 : _GEN_1068; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3117 = igen_1_io_fire ? _GEN_2093 : _GEN_1069; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3118 = igen_1_io_fire ? _GEN_2094 : _GEN_1070; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3119 = igen_1_io_fire ? _GEN_2095 : _GEN_1071; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3120 = igen_1_io_fire ? _GEN_2096 : _GEN_1072; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3121 = igen_1_io_fire ? _GEN_2097 : _GEN_1073; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3122 = igen_1_io_fire ? _GEN_2098 : _GEN_1074; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3123 = igen_1_io_fire ? _GEN_2099 : _GEN_1075; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3124 = igen_1_io_fire ? _GEN_2100 : _GEN_1076; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3125 = igen_1_io_fire ? _GEN_2101 : _GEN_1077; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3126 = igen_1_io_fire ? _GEN_2102 : _GEN_1078; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3127 = igen_1_io_fire ? _GEN_2103 : _GEN_1079; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3128 = igen_1_io_fire ? _GEN_2104 : _GEN_1080; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3129 = igen_1_io_fire ? _GEN_2105 : _GEN_1081; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3130 = igen_1_io_fire ? _GEN_2106 : _GEN_1082; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3131 = igen_1_io_fire ? _GEN_2107 : _GEN_1083; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3132 = igen_1_io_fire ? _GEN_2108 : _GEN_1084; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3133 = igen_1_io_fire ? _GEN_2109 : _GEN_1085; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3134 = igen_1_io_fire ? _GEN_2110 : _GEN_1086; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3135 = igen_1_io_fire ? _GEN_2111 : _GEN_1087; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3136 = igen_1_io_fire ? _GEN_2112 : _GEN_1088; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3137 = igen_1_io_fire ? _GEN_2113 : _GEN_1089; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3138 = igen_1_io_fire ? _GEN_2114 : _GEN_1090; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3139 = igen_1_io_fire ? _GEN_2115 : _GEN_1091; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3140 = igen_1_io_fire ? _GEN_2116 : _GEN_1092; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3141 = igen_1_io_fire ? _GEN_2117 : _GEN_1093; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3142 = igen_1_io_fire ? _GEN_2118 : _GEN_1094; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3143 = igen_1_io_fire ? _GEN_2119 : _GEN_1095; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3144 = igen_1_io_fire ? _GEN_2120 : _GEN_1096; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3145 = igen_1_io_fire ? _GEN_2121 : _GEN_1097; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3146 = igen_1_io_fire ? _GEN_2122 : _GEN_1098; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3147 = igen_1_io_fire ? _GEN_2123 : _GEN_1099; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3148 = igen_1_io_fire ? _GEN_2124 : _GEN_1100; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3149 = igen_1_io_fire ? _GEN_2125 : _GEN_1101; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3150 = igen_1_io_fire ? _GEN_2126 : _GEN_1102; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3151 = igen_1_io_fire ? _GEN_2127 : _GEN_1103; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3152 = igen_1_io_fire ? _GEN_2128 : _GEN_1104; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3153 = igen_1_io_fire ? _GEN_2129 : _GEN_1105; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3154 = igen_1_io_fire ? _GEN_2130 : _GEN_1106; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3155 = igen_1_io_fire ? _GEN_2131 : _GEN_1107; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3156 = igen_1_io_fire ? _GEN_2132 : _GEN_1108; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3157 = igen_1_io_fire ? _GEN_2133 : _GEN_1109; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3158 = igen_1_io_fire ? _GEN_2134 : _GEN_1110; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3159 = igen_1_io_fire ? _GEN_2135 : _GEN_1111; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3160 = igen_1_io_fire ? _GEN_2136 : _GEN_1112; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3161 = igen_1_io_fire ? _GEN_2137 : _GEN_1113; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3162 = igen_1_io_fire ? _GEN_2138 : _GEN_1114; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3163 = igen_1_io_fire ? _GEN_2139 : _GEN_1115; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3164 = igen_1_io_fire ? _GEN_2140 : _GEN_1116; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3165 = igen_1_io_fire ? _GEN_2141 : _GEN_1117; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3166 = igen_1_io_fire ? _GEN_2142 : _GEN_1118; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3167 = igen_1_io_fire ? _GEN_2143 : _GEN_1119; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3168 = igen_1_io_fire ? _GEN_2144 : _GEN_1120; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3169 = igen_1_io_fire ? _GEN_2145 : _GEN_1121; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3170 = igen_1_io_fire ? _GEN_2146 : _GEN_1122; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3171 = igen_1_io_fire ? _GEN_2147 : _GEN_1123; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3172 = igen_1_io_fire ? _GEN_2148 : _GEN_1124; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3173 = igen_1_io_fire ? _GEN_2149 : _GEN_1125; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3174 = igen_1_io_fire ? _GEN_2150 : _GEN_1126; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3175 = igen_1_io_fire ? _GEN_2151 : _GEN_1127; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3176 = igen_1_io_fire ? _GEN_2152 : _GEN_1128; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3177 = igen_1_io_fire ? _GEN_2153 : _GEN_1129; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3178 = igen_1_io_fire ? _GEN_2154 : _GEN_1130; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3179 = igen_1_io_fire ? _GEN_2155 : _GEN_1131; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3180 = igen_1_io_fire ? _GEN_2156 : _GEN_1132; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3181 = igen_1_io_fire ? _GEN_2157 : _GEN_1133; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3182 = igen_1_io_fire ? _GEN_2158 : _GEN_1134; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3183 = igen_1_io_fire ? _GEN_2159 : _GEN_1135; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3184 = igen_1_io_fire ? _GEN_2160 : _GEN_1136; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3185 = igen_1_io_fire ? _GEN_2161 : _GEN_1137; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3186 = igen_1_io_fire ? _GEN_2162 : _GEN_1138; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3187 = igen_1_io_fire ? _GEN_2163 : _GEN_1139; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3188 = igen_1_io_fire ? _GEN_2164 : _GEN_1140; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3189 = igen_1_io_fire ? _GEN_2165 : _GEN_1141; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3190 = igen_1_io_fire ? _GEN_2166 : _GEN_1142; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3191 = igen_1_io_fire ? _GEN_2167 : _GEN_1143; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3192 = igen_1_io_fire ? _GEN_2168 : _GEN_1144; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3193 = igen_1_io_fire ? _GEN_2169 : _GEN_1145; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3194 = igen_1_io_fire ? _GEN_2170 : _GEN_1146; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3195 = igen_1_io_fire ? _GEN_2171 : _GEN_1147; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3196 = igen_1_io_fire ? _GEN_2172 : _GEN_1148; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3197 = igen_1_io_fire ? _GEN_2173 : _GEN_1149; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3198 = igen_1_io_fire ? _GEN_2174 : _GEN_1150; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3199 = igen_1_io_fire ? _GEN_2175 : _GEN_1151; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_3200 = igen_1_io_fire ? _GEN_2176 : _GEN_1152; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3201 = igen_1_io_fire ? _GEN_2177 : _GEN_1153; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3202 = igen_1_io_fire ? _GEN_2178 : _GEN_1154; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3203 = igen_1_io_fire ? _GEN_2179 : _GEN_1155; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3204 = igen_1_io_fire ? _GEN_2180 : _GEN_1156; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3205 = igen_1_io_fire ? _GEN_2181 : _GEN_1157; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3206 = igen_1_io_fire ? _GEN_2182 : _GEN_1158; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3207 = igen_1_io_fire ? _GEN_2183 : _GEN_1159; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3208 = igen_1_io_fire ? _GEN_2184 : _GEN_1160; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3209 = igen_1_io_fire ? _GEN_2185 : _GEN_1161; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3210 = igen_1_io_fire ? _GEN_2186 : _GEN_1162; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3211 = igen_1_io_fire ? _GEN_2187 : _GEN_1163; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3212 = igen_1_io_fire ? _GEN_2188 : _GEN_1164; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3213 = igen_1_io_fire ? _GEN_2189 : _GEN_1165; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3214 = igen_1_io_fire ? _GEN_2190 : _GEN_1166; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3215 = igen_1_io_fire ? _GEN_2191 : _GEN_1167; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3216 = igen_1_io_fire ? _GEN_2192 : _GEN_1168; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3217 = igen_1_io_fire ? _GEN_2193 : _GEN_1169; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3218 = igen_1_io_fire ? _GEN_2194 : _GEN_1170; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3219 = igen_1_io_fire ? _GEN_2195 : _GEN_1171; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3220 = igen_1_io_fire ? _GEN_2196 : _GEN_1172; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3221 = igen_1_io_fire ? _GEN_2197 : _GEN_1173; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3222 = igen_1_io_fire ? _GEN_2198 : _GEN_1174; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3223 = igen_1_io_fire ? _GEN_2199 : _GEN_1175; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3224 = igen_1_io_fire ? _GEN_2200 : _GEN_1176; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3225 = igen_1_io_fire ? _GEN_2201 : _GEN_1177; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3226 = igen_1_io_fire ? _GEN_2202 : _GEN_1178; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3227 = igen_1_io_fire ? _GEN_2203 : _GEN_1179; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3228 = igen_1_io_fire ? _GEN_2204 : _GEN_1180; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3229 = igen_1_io_fire ? _GEN_2205 : _GEN_1181; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3230 = igen_1_io_fire ? _GEN_2206 : _GEN_1182; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3231 = igen_1_io_fire ? _GEN_2207 : _GEN_1183; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3232 = igen_1_io_fire ? _GEN_2208 : _GEN_1184; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3233 = igen_1_io_fire ? _GEN_2209 : _GEN_1185; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3234 = igen_1_io_fire ? _GEN_2210 : _GEN_1186; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3235 = igen_1_io_fire ? _GEN_2211 : _GEN_1187; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3236 = igen_1_io_fire ? _GEN_2212 : _GEN_1188; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3237 = igen_1_io_fire ? _GEN_2213 : _GEN_1189; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3238 = igen_1_io_fire ? _GEN_2214 : _GEN_1190; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3239 = igen_1_io_fire ? _GEN_2215 : _GEN_1191; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3240 = igen_1_io_fire ? _GEN_2216 : _GEN_1192; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3241 = igen_1_io_fire ? _GEN_2217 : _GEN_1193; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3242 = igen_1_io_fire ? _GEN_2218 : _GEN_1194; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3243 = igen_1_io_fire ? _GEN_2219 : _GEN_1195; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3244 = igen_1_io_fire ? _GEN_2220 : _GEN_1196; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3245 = igen_1_io_fire ? _GEN_2221 : _GEN_1197; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3246 = igen_1_io_fire ? _GEN_2222 : _GEN_1198; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3247 = igen_1_io_fire ? _GEN_2223 : _GEN_1199; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3248 = igen_1_io_fire ? _GEN_2224 : _GEN_1200; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3249 = igen_1_io_fire ? _GEN_2225 : _GEN_1201; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3250 = igen_1_io_fire ? _GEN_2226 : _GEN_1202; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3251 = igen_1_io_fire ? _GEN_2227 : _GEN_1203; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3252 = igen_1_io_fire ? _GEN_2228 : _GEN_1204; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3253 = igen_1_io_fire ? _GEN_2229 : _GEN_1205; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3254 = igen_1_io_fire ? _GEN_2230 : _GEN_1206; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3255 = igen_1_io_fire ? _GEN_2231 : _GEN_1207; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3256 = igen_1_io_fire ? _GEN_2232 : _GEN_1208; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3257 = igen_1_io_fire ? _GEN_2233 : _GEN_1209; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3258 = igen_1_io_fire ? _GEN_2234 : _GEN_1210; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3259 = igen_1_io_fire ? _GEN_2235 : _GEN_1211; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3260 = igen_1_io_fire ? _GEN_2236 : _GEN_1212; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3261 = igen_1_io_fire ? _GEN_2237 : _GEN_1213; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3262 = igen_1_io_fire ? _GEN_2238 : _GEN_1214; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3263 = igen_1_io_fire ? _GEN_2239 : _GEN_1215; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3264 = igen_1_io_fire ? _GEN_2240 : _GEN_1216; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3265 = igen_1_io_fire ? _GEN_2241 : _GEN_1217; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3266 = igen_1_io_fire ? _GEN_2242 : _GEN_1218; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3267 = igen_1_io_fire ? _GEN_2243 : _GEN_1219; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3268 = igen_1_io_fire ? _GEN_2244 : _GEN_1220; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3269 = igen_1_io_fire ? _GEN_2245 : _GEN_1221; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3270 = igen_1_io_fire ? _GEN_2246 : _GEN_1222; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3271 = igen_1_io_fire ? _GEN_2247 : _GEN_1223; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3272 = igen_1_io_fire ? _GEN_2248 : _GEN_1224; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3273 = igen_1_io_fire ? _GEN_2249 : _GEN_1225; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3274 = igen_1_io_fire ? _GEN_2250 : _GEN_1226; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3275 = igen_1_io_fire ? _GEN_2251 : _GEN_1227; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3276 = igen_1_io_fire ? _GEN_2252 : _GEN_1228; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3277 = igen_1_io_fire ? _GEN_2253 : _GEN_1229; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3278 = igen_1_io_fire ? _GEN_2254 : _GEN_1230; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3279 = igen_1_io_fire ? _GEN_2255 : _GEN_1231; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3280 = igen_1_io_fire ? _GEN_2256 : _GEN_1232; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3281 = igen_1_io_fire ? _GEN_2257 : _GEN_1233; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3282 = igen_1_io_fire ? _GEN_2258 : _GEN_1234; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3283 = igen_1_io_fire ? _GEN_2259 : _GEN_1235; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3284 = igen_1_io_fire ? _GEN_2260 : _GEN_1236; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3285 = igen_1_io_fire ? _GEN_2261 : _GEN_1237; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3286 = igen_1_io_fire ? _GEN_2262 : _GEN_1238; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3287 = igen_1_io_fire ? _GEN_2263 : _GEN_1239; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3288 = igen_1_io_fire ? _GEN_2264 : _GEN_1240; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3289 = igen_1_io_fire ? _GEN_2265 : _GEN_1241; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3290 = igen_1_io_fire ? _GEN_2266 : _GEN_1242; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3291 = igen_1_io_fire ? _GEN_2267 : _GEN_1243; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3292 = igen_1_io_fire ? _GEN_2268 : _GEN_1244; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3293 = igen_1_io_fire ? _GEN_2269 : _GEN_1245; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3294 = igen_1_io_fire ? _GEN_2270 : _GEN_1246; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3295 = igen_1_io_fire ? _GEN_2271 : _GEN_1247; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3296 = igen_1_io_fire ? _GEN_2272 : _GEN_1248; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3297 = igen_1_io_fire ? _GEN_2273 : _GEN_1249; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3298 = igen_1_io_fire ? _GEN_2274 : _GEN_1250; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3299 = igen_1_io_fire ? _GEN_2275 : _GEN_1251; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3300 = igen_1_io_fire ? _GEN_2276 : _GEN_1252; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3301 = igen_1_io_fire ? _GEN_2277 : _GEN_1253; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3302 = igen_1_io_fire ? _GEN_2278 : _GEN_1254; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3303 = igen_1_io_fire ? _GEN_2279 : _GEN_1255; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3304 = igen_1_io_fire ? _GEN_2280 : _GEN_1256; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3305 = igen_1_io_fire ? _GEN_2281 : _GEN_1257; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3306 = igen_1_io_fire ? _GEN_2282 : _GEN_1258; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3307 = igen_1_io_fire ? _GEN_2283 : _GEN_1259; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3308 = igen_1_io_fire ? _GEN_2284 : _GEN_1260; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3309 = igen_1_io_fire ? _GEN_2285 : _GEN_1261; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3310 = igen_1_io_fire ? _GEN_2286 : _GEN_1262; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3311 = igen_1_io_fire ? _GEN_2287 : _GEN_1263; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3312 = igen_1_io_fire ? _GEN_2288 : _GEN_1264; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3313 = igen_1_io_fire ? _GEN_2289 : _GEN_1265; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3314 = igen_1_io_fire ? _GEN_2290 : _GEN_1266; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3315 = igen_1_io_fire ? _GEN_2291 : _GEN_1267; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3316 = igen_1_io_fire ? _GEN_2292 : _GEN_1268; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3317 = igen_1_io_fire ? _GEN_2293 : _GEN_1269; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3318 = igen_1_io_fire ? _GEN_2294 : _GEN_1270; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3319 = igen_1_io_fire ? _GEN_2295 : _GEN_1271; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3320 = igen_1_io_fire ? _GEN_2296 : _GEN_1272; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3321 = igen_1_io_fire ? _GEN_2297 : _GEN_1273; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3322 = igen_1_io_fire ? _GEN_2298 : _GEN_1274; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3323 = igen_1_io_fire ? _GEN_2299 : _GEN_1275; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3324 = igen_1_io_fire ? _GEN_2300 : _GEN_1276; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3325 = igen_1_io_fire ? _GEN_2301 : _GEN_1277; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3326 = igen_1_io_fire ? _GEN_2302 : _GEN_1278; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3327 = igen_1_io_fire ? _GEN_2303 : _GEN_1279; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3328 = igen_1_io_fire ? _GEN_2304 : _GEN_1280; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3329 = igen_1_io_fire ? _GEN_2305 : _GEN_1281; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3330 = igen_1_io_fire ? _GEN_2306 : _GEN_1282; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3331 = igen_1_io_fire ? _GEN_2307 : _GEN_1283; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3332 = igen_1_io_fire ? _GEN_2308 : _GEN_1284; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3333 = igen_1_io_fire ? _GEN_2309 : _GEN_1285; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3334 = igen_1_io_fire ? _GEN_2310 : _GEN_1286; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3335 = igen_1_io_fire ? _GEN_2311 : _GEN_1287; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3336 = igen_1_io_fire ? _GEN_2312 : _GEN_1288; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3337 = igen_1_io_fire ? _GEN_2313 : _GEN_1289; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3338 = igen_1_io_fire ? _GEN_2314 : _GEN_1290; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3339 = igen_1_io_fire ? _GEN_2315 : _GEN_1291; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3340 = igen_1_io_fire ? _GEN_2316 : _GEN_1292; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3341 = igen_1_io_fire ? _GEN_2317 : _GEN_1293; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3342 = igen_1_io_fire ? _GEN_2318 : _GEN_1294; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3343 = igen_1_io_fire ? _GEN_2319 : _GEN_1295; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3344 = igen_1_io_fire ? _GEN_2320 : _GEN_1296; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3345 = igen_1_io_fire ? _GEN_2321 : _GEN_1297; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3346 = igen_1_io_fire ? _GEN_2322 : _GEN_1298; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3347 = igen_1_io_fire ? _GEN_2323 : _GEN_1299; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3348 = igen_1_io_fire ? _GEN_2324 : _GEN_1300; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3349 = igen_1_io_fire ? _GEN_2325 : _GEN_1301; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3350 = igen_1_io_fire ? _GEN_2326 : _GEN_1302; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3351 = igen_1_io_fire ? _GEN_2327 : _GEN_1303; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3352 = igen_1_io_fire ? _GEN_2328 : _GEN_1304; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3353 = igen_1_io_fire ? _GEN_2329 : _GEN_1305; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3354 = igen_1_io_fire ? _GEN_2330 : _GEN_1306; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3355 = igen_1_io_fire ? _GEN_2331 : _GEN_1307; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3356 = igen_1_io_fire ? _GEN_2332 : _GEN_1308; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3357 = igen_1_io_fire ? _GEN_2333 : _GEN_1309; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3358 = igen_1_io_fire ? _GEN_2334 : _GEN_1310; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3359 = igen_1_io_fire ? _GEN_2335 : _GEN_1311; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3360 = igen_1_io_fire ? _GEN_2336 : _GEN_1312; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3361 = igen_1_io_fire ? _GEN_2337 : _GEN_1313; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3362 = igen_1_io_fire ? _GEN_2338 : _GEN_1314; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3363 = igen_1_io_fire ? _GEN_2339 : _GEN_1315; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3364 = igen_1_io_fire ? _GEN_2340 : _GEN_1316; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3365 = igen_1_io_fire ? _GEN_2341 : _GEN_1317; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3366 = igen_1_io_fire ? _GEN_2342 : _GEN_1318; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3367 = igen_1_io_fire ? _GEN_2343 : _GEN_1319; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3368 = igen_1_io_fire ? _GEN_2344 : _GEN_1320; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3369 = igen_1_io_fire ? _GEN_2345 : _GEN_1321; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3370 = igen_1_io_fire ? _GEN_2346 : _GEN_1322; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3371 = igen_1_io_fire ? _GEN_2347 : _GEN_1323; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3372 = igen_1_io_fire ? _GEN_2348 : _GEN_1324; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3373 = igen_1_io_fire ? _GEN_2349 : _GEN_1325; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3374 = igen_1_io_fire ? _GEN_2350 : _GEN_1326; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3375 = igen_1_io_fire ? _GEN_2351 : _GEN_1327; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3376 = igen_1_io_fire ? _GEN_2352 : _GEN_1328; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3377 = igen_1_io_fire ? _GEN_2353 : _GEN_1329; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3378 = igen_1_io_fire ? _GEN_2354 : _GEN_1330; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3379 = igen_1_io_fire ? _GEN_2355 : _GEN_1331; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3380 = igen_1_io_fire ? _GEN_2356 : _GEN_1332; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3381 = igen_1_io_fire ? _GEN_2357 : _GEN_1333; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3382 = igen_1_io_fire ? _GEN_2358 : _GEN_1334; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3383 = igen_1_io_fire ? _GEN_2359 : _GEN_1335; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3384 = igen_1_io_fire ? _GEN_2360 : _GEN_1336; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3385 = igen_1_io_fire ? _GEN_2361 : _GEN_1337; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3386 = igen_1_io_fire ? _GEN_2362 : _GEN_1338; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3387 = igen_1_io_fire ? _GEN_2363 : _GEN_1339; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3388 = igen_1_io_fire ? _GEN_2364 : _GEN_1340; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3389 = igen_1_io_fire ? _GEN_2365 : _GEN_1341; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3390 = igen_1_io_fire ? _GEN_2366 : _GEN_1342; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3391 = igen_1_io_fire ? _GEN_2367 : _GEN_1343; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3392 = igen_1_io_fire ? _GEN_2368 : _GEN_1344; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3393 = igen_1_io_fire ? _GEN_2369 : _GEN_1345; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3394 = igen_1_io_fire ? _GEN_2370 : _GEN_1346; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3395 = igen_1_io_fire ? _GEN_2371 : _GEN_1347; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3396 = igen_1_io_fire ? _GEN_2372 : _GEN_1348; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3397 = igen_1_io_fire ? _GEN_2373 : _GEN_1349; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3398 = igen_1_io_fire ? _GEN_2374 : _GEN_1350; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3399 = igen_1_io_fire ? _GEN_2375 : _GEN_1351; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3400 = igen_1_io_fire ? _GEN_2376 : _GEN_1352; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3401 = igen_1_io_fire ? _GEN_2377 : _GEN_1353; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3402 = igen_1_io_fire ? _GEN_2378 : _GEN_1354; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3403 = igen_1_io_fire ? _GEN_2379 : _GEN_1355; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3404 = igen_1_io_fire ? _GEN_2380 : _GEN_1356; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3405 = igen_1_io_fire ? _GEN_2381 : _GEN_1357; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3406 = igen_1_io_fire ? _GEN_2382 : _GEN_1358; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3407 = igen_1_io_fire ? _GEN_2383 : _GEN_1359; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3408 = igen_1_io_fire ? _GEN_2384 : _GEN_1360; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3409 = igen_1_io_fire ? _GEN_2385 : _GEN_1361; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3410 = igen_1_io_fire ? _GEN_2386 : _GEN_1362; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3411 = igen_1_io_fire ? _GEN_2387 : _GEN_1363; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3412 = igen_1_io_fire ? _GEN_2388 : _GEN_1364; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3413 = igen_1_io_fire ? _GEN_2389 : _GEN_1365; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3414 = igen_1_io_fire ? _GEN_2390 : _GEN_1366; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3415 = igen_1_io_fire ? _GEN_2391 : _GEN_1367; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3416 = igen_1_io_fire ? _GEN_2392 : _GEN_1368; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3417 = igen_1_io_fire ? _GEN_2393 : _GEN_1369; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3418 = igen_1_io_fire ? _GEN_2394 : _GEN_1370; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3419 = igen_1_io_fire ? _GEN_2395 : _GEN_1371; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3420 = igen_1_io_fire ? _GEN_2396 : _GEN_1372; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3421 = igen_1_io_fire ? _GEN_2397 : _GEN_1373; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3422 = igen_1_io_fire ? _GEN_2398 : _GEN_1374; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3423 = igen_1_io_fire ? _GEN_2399 : _GEN_1375; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3424 = igen_1_io_fire ? _GEN_2400 : _GEN_1376; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3425 = igen_1_io_fire ? _GEN_2401 : _GEN_1377; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3426 = igen_1_io_fire ? _GEN_2402 : _GEN_1378; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3427 = igen_1_io_fire ? _GEN_2403 : _GEN_1379; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3428 = igen_1_io_fire ? _GEN_2404 : _GEN_1380; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3429 = igen_1_io_fire ? _GEN_2405 : _GEN_1381; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3430 = igen_1_io_fire ? _GEN_2406 : _GEN_1382; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3431 = igen_1_io_fire ? _GEN_2407 : _GEN_1383; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3432 = igen_1_io_fire ? _GEN_2408 : _GEN_1384; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3433 = igen_1_io_fire ? _GEN_2409 : _GEN_1385; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3434 = igen_1_io_fire ? _GEN_2410 : _GEN_1386; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3435 = igen_1_io_fire ? _GEN_2411 : _GEN_1387; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3436 = igen_1_io_fire ? _GEN_2412 : _GEN_1388; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3437 = igen_1_io_fire ? _GEN_2413 : _GEN_1389; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3438 = igen_1_io_fire ? _GEN_2414 : _GEN_1390; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3439 = igen_1_io_fire ? _GEN_2415 : _GEN_1391; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3440 = igen_1_io_fire ? _GEN_2416 : _GEN_1392; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3441 = igen_1_io_fire ? _GEN_2417 : _GEN_1393; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3442 = igen_1_io_fire ? _GEN_2418 : _GEN_1394; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3443 = igen_1_io_fire ? _GEN_2419 : _GEN_1395; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3444 = igen_1_io_fire ? _GEN_2420 : _GEN_1396; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3445 = igen_1_io_fire ? _GEN_2421 : _GEN_1397; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3446 = igen_1_io_fire ? _GEN_2422 : _GEN_1398; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3447 = igen_1_io_fire ? _GEN_2423 : _GEN_1399; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3448 = igen_1_io_fire ? _GEN_2424 : _GEN_1400; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3449 = igen_1_io_fire ? _GEN_2425 : _GEN_1401; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3450 = igen_1_io_fire ? _GEN_2426 : _GEN_1402; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3451 = igen_1_io_fire ? _GEN_2427 : _GEN_1403; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3452 = igen_1_io_fire ? _GEN_2428 : _GEN_1404; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3453 = igen_1_io_fire ? _GEN_2429 : _GEN_1405; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3454 = igen_1_io_fire ? _GEN_2430 : _GEN_1406; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3455 = igen_1_io_fire ? _GEN_2431 : _GEN_1407; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3456 = igen_1_io_fire ? _GEN_2432 : _GEN_1408; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3457 = igen_1_io_fire ? _GEN_2433 : _GEN_1409; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3458 = igen_1_io_fire ? _GEN_2434 : _GEN_1410; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3459 = igen_1_io_fire ? _GEN_2435 : _GEN_1411; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3460 = igen_1_io_fire ? _GEN_2436 : _GEN_1412; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3461 = igen_1_io_fire ? _GEN_2437 : _GEN_1413; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3462 = igen_1_io_fire ? _GEN_2438 : _GEN_1414; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3463 = igen_1_io_fire ? _GEN_2439 : _GEN_1415; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3464 = igen_1_io_fire ? _GEN_2440 : _GEN_1416; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3465 = igen_1_io_fire ? _GEN_2441 : _GEN_1417; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3466 = igen_1_io_fire ? _GEN_2442 : _GEN_1418; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3467 = igen_1_io_fire ? _GEN_2443 : _GEN_1419; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3468 = igen_1_io_fire ? _GEN_2444 : _GEN_1420; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3469 = igen_1_io_fire ? _GEN_2445 : _GEN_1421; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3470 = igen_1_io_fire ? _GEN_2446 : _GEN_1422; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3471 = igen_1_io_fire ? _GEN_2447 : _GEN_1423; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3472 = igen_1_io_fire ? _GEN_2448 : _GEN_1424; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3473 = igen_1_io_fire ? _GEN_2449 : _GEN_1425; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3474 = igen_1_io_fire ? _GEN_2450 : _GEN_1426; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3475 = igen_1_io_fire ? _GEN_2451 : _GEN_1427; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3476 = igen_1_io_fire ? _GEN_2452 : _GEN_1428; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3477 = igen_1_io_fire ? _GEN_2453 : _GEN_1429; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3478 = igen_1_io_fire ? _GEN_2454 : _GEN_1430; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3479 = igen_1_io_fire ? _GEN_2455 : _GEN_1431; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3480 = igen_1_io_fire ? _GEN_2456 : _GEN_1432; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3481 = igen_1_io_fire ? _GEN_2457 : _GEN_1433; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3482 = igen_1_io_fire ? _GEN_2458 : _GEN_1434; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3483 = igen_1_io_fire ? _GEN_2459 : _GEN_1435; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3484 = igen_1_io_fire ? _GEN_2460 : _GEN_1436; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3485 = igen_1_io_fire ? _GEN_2461 : _GEN_1437; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3486 = igen_1_io_fire ? _GEN_2462 : _GEN_1438; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3487 = igen_1_io_fire ? _GEN_2463 : _GEN_1439; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3488 = igen_1_io_fire ? _GEN_2464 : _GEN_1440; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3489 = igen_1_io_fire ? _GEN_2465 : _GEN_1441; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3490 = igen_1_io_fire ? _GEN_2466 : _GEN_1442; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3491 = igen_1_io_fire ? _GEN_2467 : _GEN_1443; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3492 = igen_1_io_fire ? _GEN_2468 : _GEN_1444; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3493 = igen_1_io_fire ? _GEN_2469 : _GEN_1445; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3494 = igen_1_io_fire ? _GEN_2470 : _GEN_1446; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3495 = igen_1_io_fire ? _GEN_2471 : _GEN_1447; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3496 = igen_1_io_fire ? _GEN_2472 : _GEN_1448; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3497 = igen_1_io_fire ? _GEN_2473 : _GEN_1449; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3498 = igen_1_io_fire ? _GEN_2474 : _GEN_1450; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3499 = igen_1_io_fire ? _GEN_2475 : _GEN_1451; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3500 = igen_1_io_fire ? _GEN_2476 : _GEN_1452; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3501 = igen_1_io_fire ? _GEN_2477 : _GEN_1453; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3502 = igen_1_io_fire ? _GEN_2478 : _GEN_1454; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3503 = igen_1_io_fire ? _GEN_2479 : _GEN_1455; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3504 = igen_1_io_fire ? _GEN_2480 : _GEN_1456; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3505 = igen_1_io_fire ? _GEN_2481 : _GEN_1457; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3506 = igen_1_io_fire ? _GEN_2482 : _GEN_1458; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3507 = igen_1_io_fire ? _GEN_2483 : _GEN_1459; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3508 = igen_1_io_fire ? _GEN_2484 : _GEN_1460; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3509 = igen_1_io_fire ? _GEN_2485 : _GEN_1461; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3510 = igen_1_io_fire ? _GEN_2486 : _GEN_1462; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3511 = igen_1_io_fire ? _GEN_2487 : _GEN_1463; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3512 = igen_1_io_fire ? _GEN_2488 : _GEN_1464; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3513 = igen_1_io_fire ? _GEN_2489 : _GEN_1465; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3514 = igen_1_io_fire ? _GEN_2490 : _GEN_1466; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3515 = igen_1_io_fire ? _GEN_2491 : _GEN_1467; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3516 = igen_1_io_fire ? _GEN_2492 : _GEN_1468; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3517 = igen_1_io_fire ? _GEN_2493 : _GEN_1469; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3518 = igen_1_io_fire ? _GEN_2494 : _GEN_1470; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3519 = igen_1_io_fire ? _GEN_2495 : _GEN_1471; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3520 = igen_1_io_fire ? _GEN_2496 : _GEN_1472; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3521 = igen_1_io_fire ? _GEN_2497 : _GEN_1473; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3522 = igen_1_io_fire ? _GEN_2498 : _GEN_1474; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3523 = igen_1_io_fire ? _GEN_2499 : _GEN_1475; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3524 = igen_1_io_fire ? _GEN_2500 : _GEN_1476; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3525 = igen_1_io_fire ? _GEN_2501 : _GEN_1477; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3526 = igen_1_io_fire ? _GEN_2502 : _GEN_1478; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3527 = igen_1_io_fire ? _GEN_2503 : _GEN_1479; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3528 = igen_1_io_fire ? _GEN_2504 : _GEN_1480; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3529 = igen_1_io_fire ? _GEN_2505 : _GEN_1481; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3530 = igen_1_io_fire ? _GEN_2506 : _GEN_1482; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3531 = igen_1_io_fire ? _GEN_2507 : _GEN_1483; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3532 = igen_1_io_fire ? _GEN_2508 : _GEN_1484; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3533 = igen_1_io_fire ? _GEN_2509 : _GEN_1485; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3534 = igen_1_io_fire ? _GEN_2510 : _GEN_1486; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3535 = igen_1_io_fire ? _GEN_2511 : _GEN_1487; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3536 = igen_1_io_fire ? _GEN_2512 : _GEN_1488; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3537 = igen_1_io_fire ? _GEN_2513 : _GEN_1489; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3538 = igen_1_io_fire ? _GEN_2514 : _GEN_1490; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3539 = igen_1_io_fire ? _GEN_2515 : _GEN_1491; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3540 = igen_1_io_fire ? _GEN_2516 : _GEN_1492; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3541 = igen_1_io_fire ? _GEN_2517 : _GEN_1493; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3542 = igen_1_io_fire ? _GEN_2518 : _GEN_1494; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3543 = igen_1_io_fire ? _GEN_2519 : _GEN_1495; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3544 = igen_1_io_fire ? _GEN_2520 : _GEN_1496; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3545 = igen_1_io_fire ? _GEN_2521 : _GEN_1497; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3546 = igen_1_io_fire ? _GEN_2522 : _GEN_1498; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3547 = igen_1_io_fire ? _GEN_2523 : _GEN_1499; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3548 = igen_1_io_fire ? _GEN_2524 : _GEN_1500; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3549 = igen_1_io_fire ? _GEN_2525 : _GEN_1501; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3550 = igen_1_io_fire ? _GEN_2526 : _GEN_1502; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3551 = igen_1_io_fire ? _GEN_2527 : _GEN_1503; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3552 = igen_1_io_fire ? _GEN_2528 : _GEN_1504; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3553 = igen_1_io_fire ? _GEN_2529 : _GEN_1505; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3554 = igen_1_io_fire ? _GEN_2530 : _GEN_1506; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3555 = igen_1_io_fire ? _GEN_2531 : _GEN_1507; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3556 = igen_1_io_fire ? _GEN_2532 : _GEN_1508; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3557 = igen_1_io_fire ? _GEN_2533 : _GEN_1509; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3558 = igen_1_io_fire ? _GEN_2534 : _GEN_1510; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3559 = igen_1_io_fire ? _GEN_2535 : _GEN_1511; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3560 = igen_1_io_fire ? _GEN_2536 : _GEN_1512; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3561 = igen_1_io_fire ? _GEN_2537 : _GEN_1513; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3562 = igen_1_io_fire ? _GEN_2538 : _GEN_1514; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3563 = igen_1_io_fire ? _GEN_2539 : _GEN_1515; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3564 = igen_1_io_fire ? _GEN_2540 : _GEN_1516; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3565 = igen_1_io_fire ? _GEN_2541 : _GEN_1517; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3566 = igen_1_io_fire ? _GEN_2542 : _GEN_1518; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3567 = igen_1_io_fire ? _GEN_2543 : _GEN_1519; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3568 = igen_1_io_fire ? _GEN_2544 : _GEN_1520; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3569 = igen_1_io_fire ? _GEN_2545 : _GEN_1521; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3570 = igen_1_io_fire ? _GEN_2546 : _GEN_1522; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3571 = igen_1_io_fire ? _GEN_2547 : _GEN_1523; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3572 = igen_1_io_fire ? _GEN_2548 : _GEN_1524; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3573 = igen_1_io_fire ? _GEN_2549 : _GEN_1525; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3574 = igen_1_io_fire ? _GEN_2550 : _GEN_1526; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3575 = igen_1_io_fire ? _GEN_2551 : _GEN_1527; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3576 = igen_1_io_fire ? _GEN_2552 : _GEN_1528; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3577 = igen_1_io_fire ? _GEN_2553 : _GEN_1529; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3578 = igen_1_io_fire ? _GEN_2554 : _GEN_1530; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3579 = igen_1_io_fire ? _GEN_2555 : _GEN_1531; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3580 = igen_1_io_fire ? _GEN_2556 : _GEN_1532; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3581 = igen_1_io_fire ? _GEN_2557 : _GEN_1533; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3582 = igen_1_io_fire ? _GEN_2558 : _GEN_1534; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3583 = igen_1_io_fire ? _GEN_2559 : _GEN_1535; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3584 = igen_1_io_fire ? _GEN_2560 : _GEN_1536; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3585 = igen_1_io_fire ? _GEN_2561 : _GEN_1537; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3586 = igen_1_io_fire ? _GEN_2562 : _GEN_1538; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3587 = igen_1_io_fire ? _GEN_2563 : _GEN_1539; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3588 = igen_1_io_fire ? _GEN_2564 : _GEN_1540; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3589 = igen_1_io_fire ? _GEN_2565 : _GEN_1541; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3590 = igen_1_io_fire ? _GEN_2566 : _GEN_1542; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3591 = igen_1_io_fire ? _GEN_2567 : _GEN_1543; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3592 = igen_1_io_fire ? _GEN_2568 : _GEN_1544; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3593 = igen_1_io_fire ? _GEN_2569 : _GEN_1545; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3594 = igen_1_io_fire ? _GEN_2570 : _GEN_1546; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3595 = igen_1_io_fire ? _GEN_2571 : _GEN_1547; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3596 = igen_1_io_fire ? _GEN_2572 : _GEN_1548; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3597 = igen_1_io_fire ? _GEN_2573 : _GEN_1549; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3598 = igen_1_io_fire ? _GEN_2574 : _GEN_1550; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3599 = igen_1_io_fire ? _GEN_2575 : _GEN_1551; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3600 = igen_1_io_fire ? _GEN_2576 : _GEN_1552; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3601 = igen_1_io_fire ? _GEN_2577 : _GEN_1553; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3602 = igen_1_io_fire ? _GEN_2578 : _GEN_1554; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3603 = igen_1_io_fire ? _GEN_2579 : _GEN_1555; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3604 = igen_1_io_fire ? _GEN_2580 : _GEN_1556; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3605 = igen_1_io_fire ? _GEN_2581 : _GEN_1557; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3606 = igen_1_io_fire ? _GEN_2582 : _GEN_1558; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3607 = igen_1_io_fire ? _GEN_2583 : _GEN_1559; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3608 = igen_1_io_fire ? _GEN_2584 : _GEN_1560; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3609 = igen_1_io_fire ? _GEN_2585 : _GEN_1561; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3610 = igen_1_io_fire ? _GEN_2586 : _GEN_1562; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3611 = igen_1_io_fire ? _GEN_2587 : _GEN_1563; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3612 = igen_1_io_fire ? _GEN_2588 : _GEN_1564; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3613 = igen_1_io_fire ? _GEN_2589 : _GEN_1565; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3614 = igen_1_io_fire ? _GEN_2590 : _GEN_1566; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3615 = igen_1_io_fire ? _GEN_2591 : _GEN_1567; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3616 = igen_1_io_fire ? _GEN_2592 : _GEN_1568; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3617 = igen_1_io_fire ? _GEN_2593 : _GEN_1569; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3618 = igen_1_io_fire ? _GEN_2594 : _GEN_1570; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3619 = igen_1_io_fire ? _GEN_2595 : _GEN_1571; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3620 = igen_1_io_fire ? _GEN_2596 : _GEN_1572; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3621 = igen_1_io_fire ? _GEN_2597 : _GEN_1573; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3622 = igen_1_io_fire ? _GEN_2598 : _GEN_1574; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3623 = igen_1_io_fire ? _GEN_2599 : _GEN_1575; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3624 = igen_1_io_fire ? _GEN_2600 : _GEN_1576; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3625 = igen_1_io_fire ? _GEN_2601 : _GEN_1577; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3626 = igen_1_io_fire ? _GEN_2602 : _GEN_1578; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3627 = igen_1_io_fire ? _GEN_2603 : _GEN_1579; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3628 = igen_1_io_fire ? _GEN_2604 : _GEN_1580; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3629 = igen_1_io_fire ? _GEN_2605 : _GEN_1581; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3630 = igen_1_io_fire ? _GEN_2606 : _GEN_1582; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3631 = igen_1_io_fire ? _GEN_2607 : _GEN_1583; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3632 = igen_1_io_fire ? _GEN_2608 : _GEN_1584; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3633 = igen_1_io_fire ? _GEN_2609 : _GEN_1585; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3634 = igen_1_io_fire ? _GEN_2610 : _GEN_1586; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3635 = igen_1_io_fire ? _GEN_2611 : _GEN_1587; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3636 = igen_1_io_fire ? _GEN_2612 : _GEN_1588; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3637 = igen_1_io_fire ? _GEN_2613 : _GEN_1589; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3638 = igen_1_io_fire ? _GEN_2614 : _GEN_1590; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3639 = igen_1_io_fire ? _GEN_2615 : _GEN_1591; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3640 = igen_1_io_fire ? _GEN_2616 : _GEN_1592; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3641 = igen_1_io_fire ? _GEN_2617 : _GEN_1593; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3642 = igen_1_io_fire ? _GEN_2618 : _GEN_1594; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3643 = igen_1_io_fire ? _GEN_2619 : _GEN_1595; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3644 = igen_1_io_fire ? _GEN_2620 : _GEN_1596; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3645 = igen_1_io_fire ? _GEN_2621 : _GEN_1597; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3646 = igen_1_io_fire ? _GEN_2622 : _GEN_1598; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3647 = igen_1_io_fire ? _GEN_2623 : _GEN_1599; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3648 = igen_1_io_fire ? _GEN_2624 : _GEN_1600; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3649 = igen_1_io_fire ? _GEN_2625 : _GEN_1601; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3650 = igen_1_io_fire ? _GEN_2626 : _GEN_1602; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3651 = igen_1_io_fire ? _GEN_2627 : _GEN_1603; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3652 = igen_1_io_fire ? _GEN_2628 : _GEN_1604; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3653 = igen_1_io_fire ? _GEN_2629 : _GEN_1605; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3654 = igen_1_io_fire ? _GEN_2630 : _GEN_1606; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3655 = igen_1_io_fire ? _GEN_2631 : _GEN_1607; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3656 = igen_1_io_fire ? _GEN_2632 : _GEN_1608; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3657 = igen_1_io_fire ? _GEN_2633 : _GEN_1609; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3658 = igen_1_io_fire ? _GEN_2634 : _GEN_1610; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3659 = igen_1_io_fire ? _GEN_2635 : _GEN_1611; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3660 = igen_1_io_fire ? _GEN_2636 : _GEN_1612; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3661 = igen_1_io_fire ? _GEN_2637 : _GEN_1613; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3662 = igen_1_io_fire ? _GEN_2638 : _GEN_1614; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3663 = igen_1_io_fire ? _GEN_2639 : _GEN_1615; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3664 = igen_1_io_fire ? _GEN_2640 : _GEN_1616; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3665 = igen_1_io_fire ? _GEN_2641 : _GEN_1617; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3666 = igen_1_io_fire ? _GEN_2642 : _GEN_1618; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3667 = igen_1_io_fire ? _GEN_2643 : _GEN_1619; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3668 = igen_1_io_fire ? _GEN_2644 : _GEN_1620; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3669 = igen_1_io_fire ? _GEN_2645 : _GEN_1621; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3670 = igen_1_io_fire ? _GEN_2646 : _GEN_1622; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3671 = igen_1_io_fire ? _GEN_2647 : _GEN_1623; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3672 = igen_1_io_fire ? _GEN_2648 : _GEN_1624; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3673 = igen_1_io_fire ? _GEN_2649 : _GEN_1625; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3674 = igen_1_io_fire ? _GEN_2650 : _GEN_1626; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3675 = igen_1_io_fire ? _GEN_2651 : _GEN_1627; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3676 = igen_1_io_fire ? _GEN_2652 : _GEN_1628; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3677 = igen_1_io_fire ? _GEN_2653 : _GEN_1629; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3678 = igen_1_io_fire ? _GEN_2654 : _GEN_1630; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3679 = igen_1_io_fire ? _GEN_2655 : _GEN_1631; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3680 = igen_1_io_fire ? _GEN_2656 : _GEN_1632; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3681 = igen_1_io_fire ? _GEN_2657 : _GEN_1633; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3682 = igen_1_io_fire ? _GEN_2658 : _GEN_1634; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3683 = igen_1_io_fire ? _GEN_2659 : _GEN_1635; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3684 = igen_1_io_fire ? _GEN_2660 : _GEN_1636; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3685 = igen_1_io_fire ? _GEN_2661 : _GEN_1637; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3686 = igen_1_io_fire ? _GEN_2662 : _GEN_1638; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3687 = igen_1_io_fire ? _GEN_2663 : _GEN_1639; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3688 = igen_1_io_fire ? _GEN_2664 : _GEN_1640; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3689 = igen_1_io_fire ? _GEN_2665 : _GEN_1641; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3690 = igen_1_io_fire ? _GEN_2666 : _GEN_1642; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3691 = igen_1_io_fire ? _GEN_2667 : _GEN_1643; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3692 = igen_1_io_fire ? _GEN_2668 : _GEN_1644; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3693 = igen_1_io_fire ? _GEN_2669 : _GEN_1645; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3694 = igen_1_io_fire ? _GEN_2670 : _GEN_1646; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3695 = igen_1_io_fire ? _GEN_2671 : _GEN_1647; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3696 = igen_1_io_fire ? _GEN_2672 : _GEN_1648; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3697 = igen_1_io_fire ? _GEN_2673 : _GEN_1649; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3698 = igen_1_io_fire ? _GEN_2674 : _GEN_1650; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3699 = igen_1_io_fire ? _GEN_2675 : _GEN_1651; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3700 = igen_1_io_fire ? _GEN_2676 : _GEN_1652; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3701 = igen_1_io_fire ? _GEN_2677 : _GEN_1653; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3702 = igen_1_io_fire ? _GEN_2678 : _GEN_1654; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3703 = igen_1_io_fire ? _GEN_2679 : _GEN_1655; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3704 = igen_1_io_fire ? _GEN_2680 : _GEN_1656; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3705 = igen_1_io_fire ? _GEN_2681 : _GEN_1657; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3706 = igen_1_io_fire ? _GEN_2682 : _GEN_1658; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3707 = igen_1_io_fire ? _GEN_2683 : _GEN_1659; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3708 = igen_1_io_fire ? _GEN_2684 : _GEN_1660; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3709 = igen_1_io_fire ? _GEN_2685 : _GEN_1661; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3710 = igen_1_io_fire ? _GEN_2686 : _GEN_1662; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3711 = igen_1_io_fire ? _GEN_2687 : _GEN_1663; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_3712 = igen_1_io_fire ? _GEN_2688 : _GEN_1664; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3713 = igen_1_io_fire ? _GEN_2689 : _GEN_1665; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3714 = igen_1_io_fire ? _GEN_2690 : _GEN_1666; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3715 = igen_1_io_fire ? _GEN_2691 : _GEN_1667; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3716 = igen_1_io_fire ? _GEN_2692 : _GEN_1668; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3717 = igen_1_io_fire ? _GEN_2693 : _GEN_1669; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3718 = igen_1_io_fire ? _GEN_2694 : _GEN_1670; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3719 = igen_1_io_fire ? _GEN_2695 : _GEN_1671; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3720 = igen_1_io_fire ? _GEN_2696 : _GEN_1672; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3721 = igen_1_io_fire ? _GEN_2697 : _GEN_1673; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3722 = igen_1_io_fire ? _GEN_2698 : _GEN_1674; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3723 = igen_1_io_fire ? _GEN_2699 : _GEN_1675; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3724 = igen_1_io_fire ? _GEN_2700 : _GEN_1676; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3725 = igen_1_io_fire ? _GEN_2701 : _GEN_1677; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3726 = igen_1_io_fire ? _GEN_2702 : _GEN_1678; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3727 = igen_1_io_fire ? _GEN_2703 : _GEN_1679; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3728 = igen_1_io_fire ? _GEN_2704 : _GEN_1680; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3729 = igen_1_io_fire ? _GEN_2705 : _GEN_1681; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3730 = igen_1_io_fire ? _GEN_2706 : _GEN_1682; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3731 = igen_1_io_fire ? _GEN_2707 : _GEN_1683; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3732 = igen_1_io_fire ? _GEN_2708 : _GEN_1684; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3733 = igen_1_io_fire ? _GEN_2709 : _GEN_1685; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3734 = igen_1_io_fire ? _GEN_2710 : _GEN_1686; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3735 = igen_1_io_fire ? _GEN_2711 : _GEN_1687; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3736 = igen_1_io_fire ? _GEN_2712 : _GEN_1688; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3737 = igen_1_io_fire ? _GEN_2713 : _GEN_1689; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3738 = igen_1_io_fire ? _GEN_2714 : _GEN_1690; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3739 = igen_1_io_fire ? _GEN_2715 : _GEN_1691; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3740 = igen_1_io_fire ? _GEN_2716 : _GEN_1692; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3741 = igen_1_io_fire ? _GEN_2717 : _GEN_1693; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3742 = igen_1_io_fire ? _GEN_2718 : _GEN_1694; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3743 = igen_1_io_fire ? _GEN_2719 : _GEN_1695; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3744 = igen_1_io_fire ? _GEN_2720 : _GEN_1696; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3745 = igen_1_io_fire ? _GEN_2721 : _GEN_1697; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3746 = igen_1_io_fire ? _GEN_2722 : _GEN_1698; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3747 = igen_1_io_fire ? _GEN_2723 : _GEN_1699; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3748 = igen_1_io_fire ? _GEN_2724 : _GEN_1700; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3749 = igen_1_io_fire ? _GEN_2725 : _GEN_1701; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3750 = igen_1_io_fire ? _GEN_2726 : _GEN_1702; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3751 = igen_1_io_fire ? _GEN_2727 : _GEN_1703; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3752 = igen_1_io_fire ? _GEN_2728 : _GEN_1704; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3753 = igen_1_io_fire ? _GEN_2729 : _GEN_1705; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3754 = igen_1_io_fire ? _GEN_2730 : _GEN_1706; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3755 = igen_1_io_fire ? _GEN_2731 : _GEN_1707; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3756 = igen_1_io_fire ? _GEN_2732 : _GEN_1708; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3757 = igen_1_io_fire ? _GEN_2733 : _GEN_1709; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3758 = igen_1_io_fire ? _GEN_2734 : _GEN_1710; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3759 = igen_1_io_fire ? _GEN_2735 : _GEN_1711; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3760 = igen_1_io_fire ? _GEN_2736 : _GEN_1712; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3761 = igen_1_io_fire ? _GEN_2737 : _GEN_1713; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3762 = igen_1_io_fire ? _GEN_2738 : _GEN_1714; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3763 = igen_1_io_fire ? _GEN_2739 : _GEN_1715; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3764 = igen_1_io_fire ? _GEN_2740 : _GEN_1716; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3765 = igen_1_io_fire ? _GEN_2741 : _GEN_1717; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3766 = igen_1_io_fire ? _GEN_2742 : _GEN_1718; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3767 = igen_1_io_fire ? _GEN_2743 : _GEN_1719; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3768 = igen_1_io_fire ? _GEN_2744 : _GEN_1720; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3769 = igen_1_io_fire ? _GEN_2745 : _GEN_1721; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3770 = igen_1_io_fire ? _GEN_2746 : _GEN_1722; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3771 = igen_1_io_fire ? _GEN_2747 : _GEN_1723; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3772 = igen_1_io_fire ? _GEN_2748 : _GEN_1724; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3773 = igen_1_io_fire ? _GEN_2749 : _GEN_1725; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3774 = igen_1_io_fire ? _GEN_2750 : _GEN_1726; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3775 = igen_1_io_fire ? _GEN_2751 : _GEN_1727; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3776 = igen_1_io_fire ? _GEN_2752 : _GEN_1728; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3777 = igen_1_io_fire ? _GEN_2753 : _GEN_1729; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3778 = igen_1_io_fire ? _GEN_2754 : _GEN_1730; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3779 = igen_1_io_fire ? _GEN_2755 : _GEN_1731; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3780 = igen_1_io_fire ? _GEN_2756 : _GEN_1732; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3781 = igen_1_io_fire ? _GEN_2757 : _GEN_1733; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3782 = igen_1_io_fire ? _GEN_2758 : _GEN_1734; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3783 = igen_1_io_fire ? _GEN_2759 : _GEN_1735; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3784 = igen_1_io_fire ? _GEN_2760 : _GEN_1736; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3785 = igen_1_io_fire ? _GEN_2761 : _GEN_1737; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3786 = igen_1_io_fire ? _GEN_2762 : _GEN_1738; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3787 = igen_1_io_fire ? _GEN_2763 : _GEN_1739; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3788 = igen_1_io_fire ? _GEN_2764 : _GEN_1740; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3789 = igen_1_io_fire ? _GEN_2765 : _GEN_1741; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3790 = igen_1_io_fire ? _GEN_2766 : _GEN_1742; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3791 = igen_1_io_fire ? _GEN_2767 : _GEN_1743; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3792 = igen_1_io_fire ? _GEN_2768 : _GEN_1744; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3793 = igen_1_io_fire ? _GEN_2769 : _GEN_1745; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3794 = igen_1_io_fire ? _GEN_2770 : _GEN_1746; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3795 = igen_1_io_fire ? _GEN_2771 : _GEN_1747; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3796 = igen_1_io_fire ? _GEN_2772 : _GEN_1748; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3797 = igen_1_io_fire ? _GEN_2773 : _GEN_1749; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3798 = igen_1_io_fire ? _GEN_2774 : _GEN_1750; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3799 = igen_1_io_fire ? _GEN_2775 : _GEN_1751; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3800 = igen_1_io_fire ? _GEN_2776 : _GEN_1752; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3801 = igen_1_io_fire ? _GEN_2777 : _GEN_1753; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3802 = igen_1_io_fire ? _GEN_2778 : _GEN_1754; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3803 = igen_1_io_fire ? _GEN_2779 : _GEN_1755; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3804 = igen_1_io_fire ? _GEN_2780 : _GEN_1756; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3805 = igen_1_io_fire ? _GEN_2781 : _GEN_1757; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3806 = igen_1_io_fire ? _GEN_2782 : _GEN_1758; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3807 = igen_1_io_fire ? _GEN_2783 : _GEN_1759; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3808 = igen_1_io_fire ? _GEN_2784 : _GEN_1760; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3809 = igen_1_io_fire ? _GEN_2785 : _GEN_1761; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3810 = igen_1_io_fire ? _GEN_2786 : _GEN_1762; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3811 = igen_1_io_fire ? _GEN_2787 : _GEN_1763; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3812 = igen_1_io_fire ? _GEN_2788 : _GEN_1764; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3813 = igen_1_io_fire ? _GEN_2789 : _GEN_1765; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3814 = igen_1_io_fire ? _GEN_2790 : _GEN_1766; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3815 = igen_1_io_fire ? _GEN_2791 : _GEN_1767; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3816 = igen_1_io_fire ? _GEN_2792 : _GEN_1768; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3817 = igen_1_io_fire ? _GEN_2793 : _GEN_1769; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3818 = igen_1_io_fire ? _GEN_2794 : _GEN_1770; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3819 = igen_1_io_fire ? _GEN_2795 : _GEN_1771; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3820 = igen_1_io_fire ? _GEN_2796 : _GEN_1772; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3821 = igen_1_io_fire ? _GEN_2797 : _GEN_1773; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3822 = igen_1_io_fire ? _GEN_2798 : _GEN_1774; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3823 = igen_1_io_fire ? _GEN_2799 : _GEN_1775; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3824 = igen_1_io_fire ? _GEN_2800 : _GEN_1776; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3825 = igen_1_io_fire ? _GEN_2801 : _GEN_1777; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3826 = igen_1_io_fire ? _GEN_2802 : _GEN_1778; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3827 = igen_1_io_fire ? _GEN_2803 : _GEN_1779; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3828 = igen_1_io_fire ? _GEN_2804 : _GEN_1780; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3829 = igen_1_io_fire ? _GEN_2805 : _GEN_1781; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3830 = igen_1_io_fire ? _GEN_2806 : _GEN_1782; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3831 = igen_1_io_fire ? _GEN_2807 : _GEN_1783; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3832 = igen_1_io_fire ? _GEN_2808 : _GEN_1784; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3833 = igen_1_io_fire ? _GEN_2809 : _GEN_1785; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3834 = igen_1_io_fire ? _GEN_2810 : _GEN_1786; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3835 = igen_1_io_fire ? _GEN_2811 : _GEN_1787; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3836 = igen_1_io_fire ? _GEN_2812 : _GEN_1788; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3837 = igen_1_io_fire ? _GEN_2813 : _GEN_1789; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3838 = igen_1_io_fire ? _GEN_2814 : _GEN_1790; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3839 = igen_1_io_fire ? _GEN_2815 : _GEN_1791; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3840 = igen_1_io_fire ? _GEN_2816 : _GEN_1792; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3841 = igen_1_io_fire ? _GEN_2817 : _GEN_1793; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3842 = igen_1_io_fire ? _GEN_2818 : _GEN_1794; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3843 = igen_1_io_fire ? _GEN_2819 : _GEN_1795; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3844 = igen_1_io_fire ? _GEN_2820 : _GEN_1796; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3845 = igen_1_io_fire ? _GEN_2821 : _GEN_1797; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3846 = igen_1_io_fire ? _GEN_2822 : _GEN_1798; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3847 = igen_1_io_fire ? _GEN_2823 : _GEN_1799; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3848 = igen_1_io_fire ? _GEN_2824 : _GEN_1800; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3849 = igen_1_io_fire ? _GEN_2825 : _GEN_1801; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3850 = igen_1_io_fire ? _GEN_2826 : _GEN_1802; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3851 = igen_1_io_fire ? _GEN_2827 : _GEN_1803; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3852 = igen_1_io_fire ? _GEN_2828 : _GEN_1804; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3853 = igen_1_io_fire ? _GEN_2829 : _GEN_1805; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3854 = igen_1_io_fire ? _GEN_2830 : _GEN_1806; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3855 = igen_1_io_fire ? _GEN_2831 : _GEN_1807; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3856 = igen_1_io_fire ? _GEN_2832 : _GEN_1808; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3857 = igen_1_io_fire ? _GEN_2833 : _GEN_1809; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3858 = igen_1_io_fire ? _GEN_2834 : _GEN_1810; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3859 = igen_1_io_fire ? _GEN_2835 : _GEN_1811; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3860 = igen_1_io_fire ? _GEN_2836 : _GEN_1812; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3861 = igen_1_io_fire ? _GEN_2837 : _GEN_1813; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3862 = igen_1_io_fire ? _GEN_2838 : _GEN_1814; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3863 = igen_1_io_fire ? _GEN_2839 : _GEN_1815; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3864 = igen_1_io_fire ? _GEN_2840 : _GEN_1816; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3865 = igen_1_io_fire ? _GEN_2841 : _GEN_1817; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3866 = igen_1_io_fire ? _GEN_2842 : _GEN_1818; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3867 = igen_1_io_fire ? _GEN_2843 : _GEN_1819; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3868 = igen_1_io_fire ? _GEN_2844 : _GEN_1820; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3869 = igen_1_io_fire ? _GEN_2845 : _GEN_1821; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3870 = igen_1_io_fire ? _GEN_2846 : _GEN_1822; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3871 = igen_1_io_fire ? _GEN_2847 : _GEN_1823; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3872 = igen_1_io_fire ? _GEN_2848 : _GEN_1824; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3873 = igen_1_io_fire ? _GEN_2849 : _GEN_1825; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3874 = igen_1_io_fire ? _GEN_2850 : _GEN_1826; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3875 = igen_1_io_fire ? _GEN_2851 : _GEN_1827; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3876 = igen_1_io_fire ? _GEN_2852 : _GEN_1828; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3877 = igen_1_io_fire ? _GEN_2853 : _GEN_1829; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3878 = igen_1_io_fire ? _GEN_2854 : _GEN_1830; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3879 = igen_1_io_fire ? _GEN_2855 : _GEN_1831; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3880 = igen_1_io_fire ? _GEN_2856 : _GEN_1832; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3881 = igen_1_io_fire ? _GEN_2857 : _GEN_1833; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3882 = igen_1_io_fire ? _GEN_2858 : _GEN_1834; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3883 = igen_1_io_fire ? _GEN_2859 : _GEN_1835; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3884 = igen_1_io_fire ? _GEN_2860 : _GEN_1836; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3885 = igen_1_io_fire ? _GEN_2861 : _GEN_1837; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3886 = igen_1_io_fire ? _GEN_2862 : _GEN_1838; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3887 = igen_1_io_fire ? _GEN_2863 : _GEN_1839; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3888 = igen_1_io_fire ? _GEN_2864 : _GEN_1840; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3889 = igen_1_io_fire ? _GEN_2865 : _GEN_1841; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3890 = igen_1_io_fire ? _GEN_2866 : _GEN_1842; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3891 = igen_1_io_fire ? _GEN_2867 : _GEN_1843; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3892 = igen_1_io_fire ? _GEN_2868 : _GEN_1844; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3893 = igen_1_io_fire ? _GEN_2869 : _GEN_1845; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3894 = igen_1_io_fire ? _GEN_2870 : _GEN_1846; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3895 = igen_1_io_fire ? _GEN_2871 : _GEN_1847; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3896 = igen_1_io_fire ? _GEN_2872 : _GEN_1848; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3897 = igen_1_io_fire ? _GEN_2873 : _GEN_1849; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3898 = igen_1_io_fire ? _GEN_2874 : _GEN_1850; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3899 = igen_1_io_fire ? _GEN_2875 : _GEN_1851; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3900 = igen_1_io_fire ? _GEN_2876 : _GEN_1852; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3901 = igen_1_io_fire ? _GEN_2877 : _GEN_1853; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3902 = igen_1_io_fire ? _GEN_2878 : _GEN_1854; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3903 = igen_1_io_fire ? _GEN_2879 : _GEN_1855; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3904 = igen_1_io_fire ? _GEN_2880 : _GEN_1856; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3905 = igen_1_io_fire ? _GEN_2881 : _GEN_1857; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3906 = igen_1_io_fire ? _GEN_2882 : _GEN_1858; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3907 = igen_1_io_fire ? _GEN_2883 : _GEN_1859; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3908 = igen_1_io_fire ? _GEN_2884 : _GEN_1860; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3909 = igen_1_io_fire ? _GEN_2885 : _GEN_1861; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3910 = igen_1_io_fire ? _GEN_2886 : _GEN_1862; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3911 = igen_1_io_fire ? _GEN_2887 : _GEN_1863; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3912 = igen_1_io_fire ? _GEN_2888 : _GEN_1864; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3913 = igen_1_io_fire ? _GEN_2889 : _GEN_1865; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3914 = igen_1_io_fire ? _GEN_2890 : _GEN_1866; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3915 = igen_1_io_fire ? _GEN_2891 : _GEN_1867; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3916 = igen_1_io_fire ? _GEN_2892 : _GEN_1868; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3917 = igen_1_io_fire ? _GEN_2893 : _GEN_1869; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3918 = igen_1_io_fire ? _GEN_2894 : _GEN_1870; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3919 = igen_1_io_fire ? _GEN_2895 : _GEN_1871; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3920 = igen_1_io_fire ? _GEN_2896 : _GEN_1872; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3921 = igen_1_io_fire ? _GEN_2897 : _GEN_1873; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3922 = igen_1_io_fire ? _GEN_2898 : _GEN_1874; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3923 = igen_1_io_fire ? _GEN_2899 : _GEN_1875; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3924 = igen_1_io_fire ? _GEN_2900 : _GEN_1876; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3925 = igen_1_io_fire ? _GEN_2901 : _GEN_1877; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3926 = igen_1_io_fire ? _GEN_2902 : _GEN_1878; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3927 = igen_1_io_fire ? _GEN_2903 : _GEN_1879; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3928 = igen_1_io_fire ? _GEN_2904 : _GEN_1880; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3929 = igen_1_io_fire ? _GEN_2905 : _GEN_1881; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3930 = igen_1_io_fire ? _GEN_2906 : _GEN_1882; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3931 = igen_1_io_fire ? _GEN_2907 : _GEN_1883; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3932 = igen_1_io_fire ? _GEN_2908 : _GEN_1884; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3933 = igen_1_io_fire ? _GEN_2909 : _GEN_1885; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3934 = igen_1_io_fire ? _GEN_2910 : _GEN_1886; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3935 = igen_1_io_fire ? _GEN_2911 : _GEN_1887; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3936 = igen_1_io_fire ? _GEN_2912 : _GEN_1888; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3937 = igen_1_io_fire ? _GEN_2913 : _GEN_1889; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3938 = igen_1_io_fire ? _GEN_2914 : _GEN_1890; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3939 = igen_1_io_fire ? _GEN_2915 : _GEN_1891; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3940 = igen_1_io_fire ? _GEN_2916 : _GEN_1892; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3941 = igen_1_io_fire ? _GEN_2917 : _GEN_1893; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3942 = igen_1_io_fire ? _GEN_2918 : _GEN_1894; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3943 = igen_1_io_fire ? _GEN_2919 : _GEN_1895; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3944 = igen_1_io_fire ? _GEN_2920 : _GEN_1896; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3945 = igen_1_io_fire ? _GEN_2921 : _GEN_1897; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3946 = igen_1_io_fire ? _GEN_2922 : _GEN_1898; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3947 = igen_1_io_fire ? _GEN_2923 : _GEN_1899; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3948 = igen_1_io_fire ? _GEN_2924 : _GEN_1900; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3949 = igen_1_io_fire ? _GEN_2925 : _GEN_1901; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3950 = igen_1_io_fire ? _GEN_2926 : _GEN_1902; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3951 = igen_1_io_fire ? _GEN_2927 : _GEN_1903; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3952 = igen_1_io_fire ? _GEN_2928 : _GEN_1904; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3953 = igen_1_io_fire ? _GEN_2929 : _GEN_1905; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3954 = igen_1_io_fire ? _GEN_2930 : _GEN_1906; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3955 = igen_1_io_fire ? _GEN_2931 : _GEN_1907; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3956 = igen_1_io_fire ? _GEN_2932 : _GEN_1908; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3957 = igen_1_io_fire ? _GEN_2933 : _GEN_1909; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3958 = igen_1_io_fire ? _GEN_2934 : _GEN_1910; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3959 = igen_1_io_fire ? _GEN_2935 : _GEN_1911; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3960 = igen_1_io_fire ? _GEN_2936 : _GEN_1912; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3961 = igen_1_io_fire ? _GEN_2937 : _GEN_1913; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3962 = igen_1_io_fire ? _GEN_2938 : _GEN_1914; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3963 = igen_1_io_fire ? _GEN_2939 : _GEN_1915; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3964 = igen_1_io_fire ? _GEN_2940 : _GEN_1916; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3965 = igen_1_io_fire ? _GEN_2941 : _GEN_1917; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3966 = igen_1_io_fire ? _GEN_2942 : _GEN_1918; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3967 = igen_1_io_fire ? _GEN_2943 : _GEN_1919; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3968 = igen_1_io_fire ? _GEN_2944 : _GEN_1920; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_3969 = igen_1_io_fire ? _GEN_2945 : _GEN_1921; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_3970 = igen_1_io_fire ? _GEN_2946 : _GEN_1922; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_3971 = igen_1_io_fire ? _GEN_2947 : _GEN_1923; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_3972 = igen_1_io_fire ? _GEN_2948 : _GEN_1924; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_3973 = igen_1_io_fire ? _GEN_2949 : _GEN_1925; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_3974 = igen_1_io_fire ? _GEN_2950 : _GEN_1926; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_3975 = igen_1_io_fire ? _GEN_2951 : _GEN_1927; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_3976 = igen_1_io_fire ? _GEN_2952 : _GEN_1928; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_3977 = igen_1_io_fire ? _GEN_2953 : _GEN_1929; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_3978 = igen_1_io_fire ? _GEN_2954 : _GEN_1930; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_3979 = igen_1_io_fire ? _GEN_2955 : _GEN_1931; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_3980 = igen_1_io_fire ? _GEN_2956 : _GEN_1932; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_3981 = igen_1_io_fire ? _GEN_2957 : _GEN_1933; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_3982 = igen_1_io_fire ? _GEN_2958 : _GEN_1934; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_3983 = igen_1_io_fire ? _GEN_2959 : _GEN_1935; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_3984 = igen_1_io_fire ? _GEN_2960 : _GEN_1936; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_3985 = igen_1_io_fire ? _GEN_2961 : _GEN_1937; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_3986 = igen_1_io_fire ? _GEN_2962 : _GEN_1938; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_3987 = igen_1_io_fire ? _GEN_2963 : _GEN_1939; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_3988 = igen_1_io_fire ? _GEN_2964 : _GEN_1940; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_3989 = igen_1_io_fire ? _GEN_2965 : _GEN_1941; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_3990 = igen_1_io_fire ? _GEN_2966 : _GEN_1942; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_3991 = igen_1_io_fire ? _GEN_2967 : _GEN_1943; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_3992 = igen_1_io_fire ? _GEN_2968 : _GEN_1944; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_3993 = igen_1_io_fire ? _GEN_2969 : _GEN_1945; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_3994 = igen_1_io_fire ? _GEN_2970 : _GEN_1946; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_3995 = igen_1_io_fire ? _GEN_2971 : _GEN_1947; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_3996 = igen_1_io_fire ? _GEN_2972 : _GEN_1948; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_3997 = igen_1_io_fire ? _GEN_2973 : _GEN_1949; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_3998 = igen_1_io_fire ? _GEN_2974 : _GEN_1950; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_3999 = igen_1_io_fire ? _GEN_2975 : _GEN_1951; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4000 = igen_1_io_fire ? _GEN_2976 : _GEN_1952; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4001 = igen_1_io_fire ? _GEN_2977 : _GEN_1953; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4002 = igen_1_io_fire ? _GEN_2978 : _GEN_1954; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4003 = igen_1_io_fire ? _GEN_2979 : _GEN_1955; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4004 = igen_1_io_fire ? _GEN_2980 : _GEN_1956; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4005 = igen_1_io_fire ? _GEN_2981 : _GEN_1957; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4006 = igen_1_io_fire ? _GEN_2982 : _GEN_1958; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4007 = igen_1_io_fire ? _GEN_2983 : _GEN_1959; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4008 = igen_1_io_fire ? _GEN_2984 : _GEN_1960; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4009 = igen_1_io_fire ? _GEN_2985 : _GEN_1961; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4010 = igen_1_io_fire ? _GEN_2986 : _GEN_1962; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4011 = igen_1_io_fire ? _GEN_2987 : _GEN_1963; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4012 = igen_1_io_fire ? _GEN_2988 : _GEN_1964; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4013 = igen_1_io_fire ? _GEN_2989 : _GEN_1965; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4014 = igen_1_io_fire ? _GEN_2990 : _GEN_1966; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4015 = igen_1_io_fire ? _GEN_2991 : _GEN_1967; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4016 = igen_1_io_fire ? _GEN_2992 : _GEN_1968; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4017 = igen_1_io_fire ? _GEN_2993 : _GEN_1969; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4018 = igen_1_io_fire ? _GEN_2994 : _GEN_1970; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4019 = igen_1_io_fire ? _GEN_2995 : _GEN_1971; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4020 = igen_1_io_fire ? _GEN_2996 : _GEN_1972; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4021 = igen_1_io_fire ? _GEN_2997 : _GEN_1973; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4022 = igen_1_io_fire ? _GEN_2998 : _GEN_1974; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4023 = igen_1_io_fire ? _GEN_2999 : _GEN_1975; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4024 = igen_1_io_fire ? _GEN_3000 : _GEN_1976; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4025 = igen_1_io_fire ? _GEN_3001 : _GEN_1977; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4026 = igen_1_io_fire ? _GEN_3002 : _GEN_1978; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4027 = igen_1_io_fire ? _GEN_3003 : _GEN_1979; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4028 = igen_1_io_fire ? _GEN_3004 : _GEN_1980; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4029 = igen_1_io_fire ? _GEN_3005 : _GEN_1981; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4030 = igen_1_io_fire ? _GEN_3006 : _GEN_1982; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4031 = igen_1_io_fire ? _GEN_3007 : _GEN_1983; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4032 = igen_1_io_fire ? _GEN_3008 : _GEN_1984; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4033 = igen_1_io_fire ? _GEN_3009 : _GEN_1985; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4034 = igen_1_io_fire ? _GEN_3010 : _GEN_1986; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4035 = igen_1_io_fire ? _GEN_3011 : _GEN_1987; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4036 = igen_1_io_fire ? _GEN_3012 : _GEN_1988; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4037 = igen_1_io_fire ? _GEN_3013 : _GEN_1989; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4038 = igen_1_io_fire ? _GEN_3014 : _GEN_1990; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4039 = igen_1_io_fire ? _GEN_3015 : _GEN_1991; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4040 = igen_1_io_fire ? _GEN_3016 : _GEN_1992; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4041 = igen_1_io_fire ? _GEN_3017 : _GEN_1993; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4042 = igen_1_io_fire ? _GEN_3018 : _GEN_1994; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4043 = igen_1_io_fire ? _GEN_3019 : _GEN_1995; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4044 = igen_1_io_fire ? _GEN_3020 : _GEN_1996; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4045 = igen_1_io_fire ? _GEN_3021 : _GEN_1997; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4046 = igen_1_io_fire ? _GEN_3022 : _GEN_1998; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4047 = igen_1_io_fire ? _GEN_3023 : _GEN_1999; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4048 = igen_1_io_fire ? _GEN_3024 : _GEN_2000; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4049 = igen_1_io_fire ? _GEN_3025 : _GEN_2001; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4050 = igen_1_io_fire ? _GEN_3026 : _GEN_2002; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4051 = igen_1_io_fire ? _GEN_3027 : _GEN_2003; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4052 = igen_1_io_fire ? _GEN_3028 : _GEN_2004; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4053 = igen_1_io_fire ? _GEN_3029 : _GEN_2005; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4054 = igen_1_io_fire ? _GEN_3030 : _GEN_2006; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4055 = igen_1_io_fire ? _GEN_3031 : _GEN_2007; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4056 = igen_1_io_fire ? _GEN_3032 : _GEN_2008; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4057 = igen_1_io_fire ? _GEN_3033 : _GEN_2009; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4058 = igen_1_io_fire ? _GEN_3034 : _GEN_2010; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4059 = igen_1_io_fire ? _GEN_3035 : _GEN_2011; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4060 = igen_1_io_fire ? _GEN_3036 : _GEN_2012; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4061 = igen_1_io_fire ? _GEN_3037 : _GEN_2013; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4062 = igen_1_io_fire ? _GEN_3038 : _GEN_2014; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4063 = igen_1_io_fire ? _GEN_3039 : _GEN_2015; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4064 = igen_1_io_fire ? _GEN_3040 : _GEN_2016; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4065 = igen_1_io_fire ? _GEN_3041 : _GEN_2017; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4066 = igen_1_io_fire ? _GEN_3042 : _GEN_2018; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4067 = igen_1_io_fire ? _GEN_3043 : _GEN_2019; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4068 = igen_1_io_fire ? _GEN_3044 : _GEN_2020; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4069 = igen_1_io_fire ? _GEN_3045 : _GEN_2021; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4070 = igen_1_io_fire ? _GEN_3046 : _GEN_2022; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4071 = igen_1_io_fire ? _GEN_3047 : _GEN_2023; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4072 = igen_1_io_fire ? _GEN_3048 : _GEN_2024; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4073 = igen_1_io_fire ? _GEN_3049 : _GEN_2025; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4074 = igen_1_io_fire ? _GEN_3050 : _GEN_2026; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4075 = igen_1_io_fire ? _GEN_3051 : _GEN_2027; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4076 = igen_1_io_fire ? _GEN_3052 : _GEN_2028; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4077 = igen_1_io_fire ? _GEN_3053 : _GEN_2029; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4078 = igen_1_io_fire ? _GEN_3054 : _GEN_2030; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4079 = igen_1_io_fire ? _GEN_3055 : _GEN_2031; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4080 = igen_1_io_fire ? _GEN_3056 : _GEN_2032; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4081 = igen_1_io_fire ? _GEN_3057 : _GEN_2033; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4082 = igen_1_io_fire ? _GEN_3058 : _GEN_2034; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4083 = igen_1_io_fire ? _GEN_3059 : _GEN_2035; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4084 = igen_1_io_fire ? _GEN_3060 : _GEN_2036; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4085 = igen_1_io_fire ? _GEN_3061 : _GEN_2037; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4086 = igen_1_io_fire ? _GEN_3062 : _GEN_2038; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4087 = igen_1_io_fire ? _GEN_3063 : _GEN_2039; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4088 = igen_1_io_fire ? _GEN_3064 : _GEN_2040; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4089 = igen_1_io_fire ? _GEN_3065 : _GEN_2041; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4090 = igen_1_io_fire ? _GEN_3066 : _GEN_2042; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4091 = igen_1_io_fire ? _GEN_3067 : _GEN_2043; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4092 = igen_1_io_fire ? _GEN_3068 : _GEN_2044; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4093 = igen_1_io_fire ? _GEN_3069 : _GEN_2045; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4094 = igen_1_io_fire ? _GEN_3070 : _GEN_2046; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4095 = igen_1_io_fire ? _GEN_3071 : _GEN_2047; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_4096 = igen_1_io_fire ? _GEN_3072 : _GEN_2048; // @[TestHarness.scala 178:25]
  wire  _igen_io_rob_ready_T_12 = rob_alloc_avail_2 & rob_alloc_fires_2 & _igen_io_rob_ready_T_1; // @[TestHarness.scala 174:72]
  wire [63:0] _rob_payload_WIRE_5 = igen_2_io_out_bits_payload; // @[TestHarness.scala 179:{72,72}]
  wire [31:0] _GEN_4097 = 7'h0 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3073; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4098 = 7'h1 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3074; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4099 = 7'h2 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3075; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4100 = 7'h3 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3076; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4101 = 7'h4 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3077; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4102 = 7'h5 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3078; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4103 = 7'h6 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3079; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4104 = 7'h7 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3080; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4105 = 7'h8 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3081; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4106 = 7'h9 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3082; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4107 = 7'ha == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3083; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4108 = 7'hb == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3084; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4109 = 7'hc == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3085; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4110 = 7'hd == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3086; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4111 = 7'he == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3087; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4112 = 7'hf == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3088; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4113 = 7'h10 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3089; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4114 = 7'h11 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3090; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4115 = 7'h12 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3091; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4116 = 7'h13 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3092; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4117 = 7'h14 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3093; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4118 = 7'h15 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3094; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4119 = 7'h16 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3095; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4120 = 7'h17 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3096; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4121 = 7'h18 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3097; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4122 = 7'h19 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3098; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4123 = 7'h1a == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3099; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4124 = 7'h1b == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3100; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4125 = 7'h1c == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3101; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4126 = 7'h1d == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3102; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4127 = 7'h1e == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3103; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4128 = 7'h1f == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3104; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4129 = 7'h20 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3105; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4130 = 7'h21 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3106; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4131 = 7'h22 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3107; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4132 = 7'h23 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3108; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4133 = 7'h24 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3109; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4134 = 7'h25 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3110; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4135 = 7'h26 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3111; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4136 = 7'h27 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3112; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4137 = 7'h28 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3113; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4138 = 7'h29 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3114; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4139 = 7'h2a == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3115; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4140 = 7'h2b == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3116; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4141 = 7'h2c == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3117; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4142 = 7'h2d == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3118; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4143 = 7'h2e == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3119; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4144 = 7'h2f == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3120; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4145 = 7'h30 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3121; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4146 = 7'h31 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3122; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4147 = 7'h32 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3123; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4148 = 7'h33 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3124; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4149 = 7'h34 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3125; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4150 = 7'h35 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3126; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4151 = 7'h36 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3127; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4152 = 7'h37 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3128; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4153 = 7'h38 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3129; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4154 = 7'h39 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3130; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4155 = 7'h3a == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3131; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4156 = 7'h3b == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3132; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4157 = 7'h3c == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3133; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4158 = 7'h3d == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3134; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4159 = 7'h3e == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3135; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4160 = 7'h3f == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3136; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4161 = 7'h40 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3137; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4162 = 7'h41 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3138; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4163 = 7'h42 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3139; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4164 = 7'h43 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3140; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4165 = 7'h44 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3141; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4166 = 7'h45 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3142; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4167 = 7'h46 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3143; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4168 = 7'h47 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3144; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4169 = 7'h48 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3145; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4170 = 7'h49 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3146; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4171 = 7'h4a == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3147; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4172 = 7'h4b == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3148; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4173 = 7'h4c == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3149; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4174 = 7'h4d == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3150; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4175 = 7'h4e == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3151; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4176 = 7'h4f == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3152; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4177 = 7'h50 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3153; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4178 = 7'h51 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3154; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4179 = 7'h52 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3155; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4180 = 7'h53 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3156; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4181 = 7'h54 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3157; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4182 = 7'h55 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3158; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4183 = 7'h56 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3159; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4184 = 7'h57 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3160; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4185 = 7'h58 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3161; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4186 = 7'h59 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3162; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4187 = 7'h5a == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3163; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4188 = 7'h5b == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3164; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4189 = 7'h5c == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3165; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4190 = 7'h5d == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3166; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4191 = 7'h5e == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3167; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4192 = 7'h5f == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3168; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4193 = 7'h60 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3169; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4194 = 7'h61 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3170; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4195 = 7'h62 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3171; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4196 = 7'h63 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3172; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4197 = 7'h64 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3173; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4198 = 7'h65 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3174; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4199 = 7'h66 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3175; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4200 = 7'h67 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3176; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4201 = 7'h68 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3177; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4202 = 7'h69 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3178; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4203 = 7'h6a == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3179; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4204 = 7'h6b == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3180; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4205 = 7'h6c == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3181; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4206 = 7'h6d == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3182; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4207 = 7'h6e == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3183; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4208 = 7'h6f == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3184; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4209 = 7'h70 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3185; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4210 = 7'h71 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3186; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4211 = 7'h72 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3187; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4212 = 7'h73 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3188; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4213 = 7'h74 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3189; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4214 = 7'h75 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3190; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4215 = 7'h76 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3191; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4216 = 7'h77 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3192; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4217 = 7'h78 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3193; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4218 = 7'h79 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3194; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4219 = 7'h7a == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3195; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4220 = 7'h7b == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3196; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4221 = 7'h7c == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3197; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4222 = 7'h7d == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3198; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4223 = 7'h7e == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3199; // @[TestHarness.scala 179:{36,36}]
  wire [31:0] _GEN_4224 = 7'h7f == rob_alloc_ids_2 ? _rob_payload_WIRE_5[63:32] : _GEN_3200; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4225 = 7'h0 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3201; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4226 = 7'h1 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3202; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4227 = 7'h2 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3203; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4228 = 7'h3 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3204; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4229 = 7'h4 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3205; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4230 = 7'h5 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3206; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4231 = 7'h6 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3207; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4232 = 7'h7 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3208; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4233 = 7'h8 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3209; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4234 = 7'h9 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3210; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4235 = 7'ha == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3211; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4236 = 7'hb == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3212; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4237 = 7'hc == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3213; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4238 = 7'hd == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3214; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4239 = 7'he == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3215; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4240 = 7'hf == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3216; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4241 = 7'h10 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3217; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4242 = 7'h11 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3218; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4243 = 7'h12 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3219; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4244 = 7'h13 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3220; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4245 = 7'h14 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3221; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4246 = 7'h15 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3222; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4247 = 7'h16 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3223; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4248 = 7'h17 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3224; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4249 = 7'h18 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3225; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4250 = 7'h19 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3226; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4251 = 7'h1a == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3227; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4252 = 7'h1b == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3228; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4253 = 7'h1c == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3229; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4254 = 7'h1d == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3230; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4255 = 7'h1e == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3231; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4256 = 7'h1f == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3232; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4257 = 7'h20 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3233; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4258 = 7'h21 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3234; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4259 = 7'h22 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3235; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4260 = 7'h23 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3236; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4261 = 7'h24 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3237; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4262 = 7'h25 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3238; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4263 = 7'h26 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3239; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4264 = 7'h27 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3240; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4265 = 7'h28 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3241; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4266 = 7'h29 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3242; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4267 = 7'h2a == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3243; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4268 = 7'h2b == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3244; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4269 = 7'h2c == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3245; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4270 = 7'h2d == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3246; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4271 = 7'h2e == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3247; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4272 = 7'h2f == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3248; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4273 = 7'h30 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3249; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4274 = 7'h31 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3250; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4275 = 7'h32 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3251; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4276 = 7'h33 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3252; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4277 = 7'h34 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3253; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4278 = 7'h35 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3254; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4279 = 7'h36 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3255; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4280 = 7'h37 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3256; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4281 = 7'h38 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3257; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4282 = 7'h39 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3258; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4283 = 7'h3a == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3259; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4284 = 7'h3b == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3260; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4285 = 7'h3c == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3261; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4286 = 7'h3d == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3262; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4287 = 7'h3e == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3263; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4288 = 7'h3f == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3264; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4289 = 7'h40 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3265; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4290 = 7'h41 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3266; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4291 = 7'h42 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3267; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4292 = 7'h43 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3268; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4293 = 7'h44 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3269; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4294 = 7'h45 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3270; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4295 = 7'h46 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3271; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4296 = 7'h47 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3272; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4297 = 7'h48 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3273; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4298 = 7'h49 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3274; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4299 = 7'h4a == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3275; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4300 = 7'h4b == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3276; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4301 = 7'h4c == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3277; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4302 = 7'h4d == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3278; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4303 = 7'h4e == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3279; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4304 = 7'h4f == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3280; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4305 = 7'h50 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3281; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4306 = 7'h51 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3282; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4307 = 7'h52 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3283; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4308 = 7'h53 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3284; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4309 = 7'h54 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3285; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4310 = 7'h55 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3286; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4311 = 7'h56 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3287; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4312 = 7'h57 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3288; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4313 = 7'h58 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3289; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4314 = 7'h59 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3290; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4315 = 7'h5a == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3291; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4316 = 7'h5b == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3292; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4317 = 7'h5c == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3293; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4318 = 7'h5d == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3294; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4319 = 7'h5e == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3295; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4320 = 7'h5f == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3296; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4321 = 7'h60 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3297; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4322 = 7'h61 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3298; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4323 = 7'h62 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3299; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4324 = 7'h63 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3300; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4325 = 7'h64 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3301; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4326 = 7'h65 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3302; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4327 = 7'h66 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3303; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4328 = 7'h67 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3304; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4329 = 7'h68 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3305; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4330 = 7'h69 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3306; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4331 = 7'h6a == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3307; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4332 = 7'h6b == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3308; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4333 = 7'h6c == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3309; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4334 = 7'h6d == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3310; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4335 = 7'h6e == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3311; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4336 = 7'h6f == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3312; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4337 = 7'h70 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3313; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4338 = 7'h71 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3314; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4339 = 7'h72 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3315; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4340 = 7'h73 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3316; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4341 = 7'h74 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3317; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4342 = 7'h75 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3318; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4343 = 7'h76 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3319; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4344 = 7'h77 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3320; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4345 = 7'h78 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3321; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4346 = 7'h79 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3322; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4347 = 7'h7a == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3323; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4348 = 7'h7b == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3324; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4349 = 7'h7c == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3325; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4350 = 7'h7d == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3326; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4351 = 7'h7e == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3327; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4352 = 7'h7f == rob_alloc_ids_2 ? _rob_payload_WIRE_5[31:16] : _GEN_3328; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4353 = 7'h0 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3329; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4354 = 7'h1 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3330; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4355 = 7'h2 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3331; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4356 = 7'h3 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3332; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4357 = 7'h4 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3333; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4358 = 7'h5 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3334; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4359 = 7'h6 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3335; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4360 = 7'h7 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3336; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4361 = 7'h8 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3337; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4362 = 7'h9 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3338; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4363 = 7'ha == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3339; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4364 = 7'hb == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3340; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4365 = 7'hc == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3341; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4366 = 7'hd == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3342; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4367 = 7'he == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3343; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4368 = 7'hf == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3344; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4369 = 7'h10 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3345; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4370 = 7'h11 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3346; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4371 = 7'h12 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3347; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4372 = 7'h13 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3348; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4373 = 7'h14 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3349; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4374 = 7'h15 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3350; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4375 = 7'h16 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3351; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4376 = 7'h17 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3352; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4377 = 7'h18 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3353; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4378 = 7'h19 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3354; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4379 = 7'h1a == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3355; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4380 = 7'h1b == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3356; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4381 = 7'h1c == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3357; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4382 = 7'h1d == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3358; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4383 = 7'h1e == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3359; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4384 = 7'h1f == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3360; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4385 = 7'h20 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3361; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4386 = 7'h21 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3362; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4387 = 7'h22 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3363; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4388 = 7'h23 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3364; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4389 = 7'h24 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3365; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4390 = 7'h25 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3366; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4391 = 7'h26 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3367; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4392 = 7'h27 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3368; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4393 = 7'h28 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3369; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4394 = 7'h29 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3370; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4395 = 7'h2a == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3371; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4396 = 7'h2b == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3372; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4397 = 7'h2c == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3373; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4398 = 7'h2d == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3374; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4399 = 7'h2e == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3375; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4400 = 7'h2f == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3376; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4401 = 7'h30 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3377; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4402 = 7'h31 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3378; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4403 = 7'h32 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3379; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4404 = 7'h33 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3380; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4405 = 7'h34 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3381; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4406 = 7'h35 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3382; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4407 = 7'h36 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3383; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4408 = 7'h37 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3384; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4409 = 7'h38 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3385; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4410 = 7'h39 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3386; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4411 = 7'h3a == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3387; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4412 = 7'h3b == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3388; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4413 = 7'h3c == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3389; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4414 = 7'h3d == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3390; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4415 = 7'h3e == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3391; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4416 = 7'h3f == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3392; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4417 = 7'h40 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3393; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4418 = 7'h41 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3394; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4419 = 7'h42 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3395; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4420 = 7'h43 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3396; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4421 = 7'h44 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3397; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4422 = 7'h45 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3398; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4423 = 7'h46 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3399; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4424 = 7'h47 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3400; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4425 = 7'h48 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3401; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4426 = 7'h49 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3402; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4427 = 7'h4a == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3403; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4428 = 7'h4b == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3404; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4429 = 7'h4c == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3405; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4430 = 7'h4d == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3406; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4431 = 7'h4e == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3407; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4432 = 7'h4f == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3408; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4433 = 7'h50 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3409; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4434 = 7'h51 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3410; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4435 = 7'h52 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3411; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4436 = 7'h53 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3412; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4437 = 7'h54 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3413; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4438 = 7'h55 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3414; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4439 = 7'h56 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3415; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4440 = 7'h57 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3416; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4441 = 7'h58 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3417; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4442 = 7'h59 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3418; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4443 = 7'h5a == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3419; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4444 = 7'h5b == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3420; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4445 = 7'h5c == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3421; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4446 = 7'h5d == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3422; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4447 = 7'h5e == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3423; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4448 = 7'h5f == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3424; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4449 = 7'h60 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3425; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4450 = 7'h61 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3426; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4451 = 7'h62 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3427; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4452 = 7'h63 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3428; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4453 = 7'h64 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3429; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4454 = 7'h65 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3430; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4455 = 7'h66 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3431; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4456 = 7'h67 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3432; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4457 = 7'h68 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3433; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4458 = 7'h69 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3434; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4459 = 7'h6a == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3435; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4460 = 7'h6b == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3436; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4461 = 7'h6c == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3437; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4462 = 7'h6d == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3438; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4463 = 7'h6e == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3439; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4464 = 7'h6f == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3440; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4465 = 7'h70 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3441; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4466 = 7'h71 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3442; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4467 = 7'h72 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3443; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4468 = 7'h73 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3444; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4469 = 7'h74 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3445; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4470 = 7'h75 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3446; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4471 = 7'h76 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3447; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4472 = 7'h77 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3448; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4473 = 7'h78 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3449; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4474 = 7'h79 == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3450; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4475 = 7'h7a == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3451; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4476 = 7'h7b == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3452; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4477 = 7'h7c == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3453; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4478 = 7'h7d == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3454; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4479 = 7'h7e == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3455; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_4480 = 7'h7f == rob_alloc_ids_2 ? _rob_payload_WIRE_5[15:0] : _GEN_3456; // @[TestHarness.scala 179:{36,36}]
  wire [1:0] _rob_egress_id_T_51 = igen_2_io_out_bits_egress_id; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4481 = 7'h0 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3457; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4482 = 7'h1 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3458; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4483 = 7'h2 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3459; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4484 = 7'h3 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3460; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4485 = 7'h4 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3461; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4486 = 7'h5 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3462; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4487 = 7'h6 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3463; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4488 = 7'h7 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3464; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4489 = 7'h8 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3465; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4490 = 7'h9 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3466; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4491 = 7'ha == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3467; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4492 = 7'hb == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3468; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4493 = 7'hc == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3469; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4494 = 7'hd == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3470; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4495 = 7'he == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3471; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4496 = 7'hf == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3472; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4497 = 7'h10 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3473; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4498 = 7'h11 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3474; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4499 = 7'h12 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3475; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4500 = 7'h13 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3476; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4501 = 7'h14 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3477; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4502 = 7'h15 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3478; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4503 = 7'h16 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3479; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4504 = 7'h17 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3480; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4505 = 7'h18 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3481; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4506 = 7'h19 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3482; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4507 = 7'h1a == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3483; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4508 = 7'h1b == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3484; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4509 = 7'h1c == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3485; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4510 = 7'h1d == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3486; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4511 = 7'h1e == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3487; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4512 = 7'h1f == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3488; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4513 = 7'h20 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3489; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4514 = 7'h21 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3490; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4515 = 7'h22 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3491; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4516 = 7'h23 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3492; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4517 = 7'h24 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3493; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4518 = 7'h25 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3494; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4519 = 7'h26 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3495; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4520 = 7'h27 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3496; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4521 = 7'h28 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3497; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4522 = 7'h29 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3498; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4523 = 7'h2a == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3499; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4524 = 7'h2b == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3500; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4525 = 7'h2c == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3501; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4526 = 7'h2d == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3502; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4527 = 7'h2e == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3503; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4528 = 7'h2f == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3504; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4529 = 7'h30 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3505; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4530 = 7'h31 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3506; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4531 = 7'h32 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3507; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4532 = 7'h33 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3508; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4533 = 7'h34 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3509; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4534 = 7'h35 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3510; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4535 = 7'h36 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3511; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4536 = 7'h37 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3512; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4537 = 7'h38 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3513; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4538 = 7'h39 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3514; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4539 = 7'h3a == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3515; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4540 = 7'h3b == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3516; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4541 = 7'h3c == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3517; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4542 = 7'h3d == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3518; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4543 = 7'h3e == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3519; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4544 = 7'h3f == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3520; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4545 = 7'h40 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3521; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4546 = 7'h41 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3522; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4547 = 7'h42 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3523; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4548 = 7'h43 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3524; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4549 = 7'h44 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3525; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4550 = 7'h45 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3526; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4551 = 7'h46 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3527; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4552 = 7'h47 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3528; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4553 = 7'h48 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3529; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4554 = 7'h49 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3530; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4555 = 7'h4a == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3531; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4556 = 7'h4b == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3532; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4557 = 7'h4c == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3533; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4558 = 7'h4d == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3534; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4559 = 7'h4e == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3535; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4560 = 7'h4f == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3536; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4561 = 7'h50 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3537; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4562 = 7'h51 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3538; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4563 = 7'h52 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3539; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4564 = 7'h53 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3540; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4565 = 7'h54 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3541; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4566 = 7'h55 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3542; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4567 = 7'h56 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3543; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4568 = 7'h57 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3544; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4569 = 7'h58 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3545; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4570 = 7'h59 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3546; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4571 = 7'h5a == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3547; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4572 = 7'h5b == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3548; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4573 = 7'h5c == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3549; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4574 = 7'h5d == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3550; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4575 = 7'h5e == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3551; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4576 = 7'h5f == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3552; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4577 = 7'h60 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3553; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4578 = 7'h61 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3554; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4579 = 7'h62 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3555; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4580 = 7'h63 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3556; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4581 = 7'h64 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3557; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4582 = 7'h65 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3558; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4583 = 7'h66 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3559; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4584 = 7'h67 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3560; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4585 = 7'h68 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3561; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4586 = 7'h69 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3562; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4587 = 7'h6a == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3563; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4588 = 7'h6b == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3564; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4589 = 7'h6c == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3565; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4590 = 7'h6d == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3566; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4591 = 7'h6e == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3567; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4592 = 7'h6f == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3568; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4593 = 7'h70 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3569; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4594 = 7'h71 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3570; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4595 = 7'h72 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3571; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4596 = 7'h73 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3572; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4597 = 7'h74 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3573; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4598 = 7'h75 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3574; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4599 = 7'h76 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3575; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4600 = 7'h77 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3576; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4601 = 7'h78 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3577; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4602 = 7'h79 == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3578; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4603 = 7'h7a == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3579; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4604 = 7'h7b == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3580; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4605 = 7'h7c == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3581; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4606 = 7'h7d == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3582; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4607 = 7'h7e == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3583; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4608 = 7'h7f == rob_alloc_ids_2 ? _rob_egress_id_T_51 : _GEN_3584; // @[TestHarness.scala 180:{36,36}]
  wire [1:0] _GEN_4609 = 7'h0 == rob_alloc_ids_2 ? 2'h2 : _GEN_3585; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4610 = 7'h1 == rob_alloc_ids_2 ? 2'h2 : _GEN_3586; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4611 = 7'h2 == rob_alloc_ids_2 ? 2'h2 : _GEN_3587; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4612 = 7'h3 == rob_alloc_ids_2 ? 2'h2 : _GEN_3588; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4613 = 7'h4 == rob_alloc_ids_2 ? 2'h2 : _GEN_3589; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4614 = 7'h5 == rob_alloc_ids_2 ? 2'h2 : _GEN_3590; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4615 = 7'h6 == rob_alloc_ids_2 ? 2'h2 : _GEN_3591; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4616 = 7'h7 == rob_alloc_ids_2 ? 2'h2 : _GEN_3592; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4617 = 7'h8 == rob_alloc_ids_2 ? 2'h2 : _GEN_3593; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4618 = 7'h9 == rob_alloc_ids_2 ? 2'h2 : _GEN_3594; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4619 = 7'ha == rob_alloc_ids_2 ? 2'h2 : _GEN_3595; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4620 = 7'hb == rob_alloc_ids_2 ? 2'h2 : _GEN_3596; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4621 = 7'hc == rob_alloc_ids_2 ? 2'h2 : _GEN_3597; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4622 = 7'hd == rob_alloc_ids_2 ? 2'h2 : _GEN_3598; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4623 = 7'he == rob_alloc_ids_2 ? 2'h2 : _GEN_3599; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4624 = 7'hf == rob_alloc_ids_2 ? 2'h2 : _GEN_3600; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4625 = 7'h10 == rob_alloc_ids_2 ? 2'h2 : _GEN_3601; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4626 = 7'h11 == rob_alloc_ids_2 ? 2'h2 : _GEN_3602; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4627 = 7'h12 == rob_alloc_ids_2 ? 2'h2 : _GEN_3603; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4628 = 7'h13 == rob_alloc_ids_2 ? 2'h2 : _GEN_3604; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4629 = 7'h14 == rob_alloc_ids_2 ? 2'h2 : _GEN_3605; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4630 = 7'h15 == rob_alloc_ids_2 ? 2'h2 : _GEN_3606; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4631 = 7'h16 == rob_alloc_ids_2 ? 2'h2 : _GEN_3607; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4632 = 7'h17 == rob_alloc_ids_2 ? 2'h2 : _GEN_3608; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4633 = 7'h18 == rob_alloc_ids_2 ? 2'h2 : _GEN_3609; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4634 = 7'h19 == rob_alloc_ids_2 ? 2'h2 : _GEN_3610; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4635 = 7'h1a == rob_alloc_ids_2 ? 2'h2 : _GEN_3611; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4636 = 7'h1b == rob_alloc_ids_2 ? 2'h2 : _GEN_3612; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4637 = 7'h1c == rob_alloc_ids_2 ? 2'h2 : _GEN_3613; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4638 = 7'h1d == rob_alloc_ids_2 ? 2'h2 : _GEN_3614; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4639 = 7'h1e == rob_alloc_ids_2 ? 2'h2 : _GEN_3615; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4640 = 7'h1f == rob_alloc_ids_2 ? 2'h2 : _GEN_3616; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4641 = 7'h20 == rob_alloc_ids_2 ? 2'h2 : _GEN_3617; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4642 = 7'h21 == rob_alloc_ids_2 ? 2'h2 : _GEN_3618; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4643 = 7'h22 == rob_alloc_ids_2 ? 2'h2 : _GEN_3619; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4644 = 7'h23 == rob_alloc_ids_2 ? 2'h2 : _GEN_3620; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4645 = 7'h24 == rob_alloc_ids_2 ? 2'h2 : _GEN_3621; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4646 = 7'h25 == rob_alloc_ids_2 ? 2'h2 : _GEN_3622; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4647 = 7'h26 == rob_alloc_ids_2 ? 2'h2 : _GEN_3623; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4648 = 7'h27 == rob_alloc_ids_2 ? 2'h2 : _GEN_3624; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4649 = 7'h28 == rob_alloc_ids_2 ? 2'h2 : _GEN_3625; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4650 = 7'h29 == rob_alloc_ids_2 ? 2'h2 : _GEN_3626; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4651 = 7'h2a == rob_alloc_ids_2 ? 2'h2 : _GEN_3627; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4652 = 7'h2b == rob_alloc_ids_2 ? 2'h2 : _GEN_3628; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4653 = 7'h2c == rob_alloc_ids_2 ? 2'h2 : _GEN_3629; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4654 = 7'h2d == rob_alloc_ids_2 ? 2'h2 : _GEN_3630; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4655 = 7'h2e == rob_alloc_ids_2 ? 2'h2 : _GEN_3631; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4656 = 7'h2f == rob_alloc_ids_2 ? 2'h2 : _GEN_3632; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4657 = 7'h30 == rob_alloc_ids_2 ? 2'h2 : _GEN_3633; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4658 = 7'h31 == rob_alloc_ids_2 ? 2'h2 : _GEN_3634; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4659 = 7'h32 == rob_alloc_ids_2 ? 2'h2 : _GEN_3635; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4660 = 7'h33 == rob_alloc_ids_2 ? 2'h2 : _GEN_3636; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4661 = 7'h34 == rob_alloc_ids_2 ? 2'h2 : _GEN_3637; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4662 = 7'h35 == rob_alloc_ids_2 ? 2'h2 : _GEN_3638; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4663 = 7'h36 == rob_alloc_ids_2 ? 2'h2 : _GEN_3639; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4664 = 7'h37 == rob_alloc_ids_2 ? 2'h2 : _GEN_3640; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4665 = 7'h38 == rob_alloc_ids_2 ? 2'h2 : _GEN_3641; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4666 = 7'h39 == rob_alloc_ids_2 ? 2'h2 : _GEN_3642; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4667 = 7'h3a == rob_alloc_ids_2 ? 2'h2 : _GEN_3643; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4668 = 7'h3b == rob_alloc_ids_2 ? 2'h2 : _GEN_3644; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4669 = 7'h3c == rob_alloc_ids_2 ? 2'h2 : _GEN_3645; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4670 = 7'h3d == rob_alloc_ids_2 ? 2'h2 : _GEN_3646; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4671 = 7'h3e == rob_alloc_ids_2 ? 2'h2 : _GEN_3647; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4672 = 7'h3f == rob_alloc_ids_2 ? 2'h2 : _GEN_3648; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4673 = 7'h40 == rob_alloc_ids_2 ? 2'h2 : _GEN_3649; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4674 = 7'h41 == rob_alloc_ids_2 ? 2'h2 : _GEN_3650; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4675 = 7'h42 == rob_alloc_ids_2 ? 2'h2 : _GEN_3651; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4676 = 7'h43 == rob_alloc_ids_2 ? 2'h2 : _GEN_3652; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4677 = 7'h44 == rob_alloc_ids_2 ? 2'h2 : _GEN_3653; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4678 = 7'h45 == rob_alloc_ids_2 ? 2'h2 : _GEN_3654; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4679 = 7'h46 == rob_alloc_ids_2 ? 2'h2 : _GEN_3655; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4680 = 7'h47 == rob_alloc_ids_2 ? 2'h2 : _GEN_3656; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4681 = 7'h48 == rob_alloc_ids_2 ? 2'h2 : _GEN_3657; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4682 = 7'h49 == rob_alloc_ids_2 ? 2'h2 : _GEN_3658; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4683 = 7'h4a == rob_alloc_ids_2 ? 2'h2 : _GEN_3659; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4684 = 7'h4b == rob_alloc_ids_2 ? 2'h2 : _GEN_3660; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4685 = 7'h4c == rob_alloc_ids_2 ? 2'h2 : _GEN_3661; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4686 = 7'h4d == rob_alloc_ids_2 ? 2'h2 : _GEN_3662; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4687 = 7'h4e == rob_alloc_ids_2 ? 2'h2 : _GEN_3663; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4688 = 7'h4f == rob_alloc_ids_2 ? 2'h2 : _GEN_3664; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4689 = 7'h50 == rob_alloc_ids_2 ? 2'h2 : _GEN_3665; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4690 = 7'h51 == rob_alloc_ids_2 ? 2'h2 : _GEN_3666; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4691 = 7'h52 == rob_alloc_ids_2 ? 2'h2 : _GEN_3667; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4692 = 7'h53 == rob_alloc_ids_2 ? 2'h2 : _GEN_3668; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4693 = 7'h54 == rob_alloc_ids_2 ? 2'h2 : _GEN_3669; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4694 = 7'h55 == rob_alloc_ids_2 ? 2'h2 : _GEN_3670; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4695 = 7'h56 == rob_alloc_ids_2 ? 2'h2 : _GEN_3671; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4696 = 7'h57 == rob_alloc_ids_2 ? 2'h2 : _GEN_3672; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4697 = 7'h58 == rob_alloc_ids_2 ? 2'h2 : _GEN_3673; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4698 = 7'h59 == rob_alloc_ids_2 ? 2'h2 : _GEN_3674; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4699 = 7'h5a == rob_alloc_ids_2 ? 2'h2 : _GEN_3675; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4700 = 7'h5b == rob_alloc_ids_2 ? 2'h2 : _GEN_3676; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4701 = 7'h5c == rob_alloc_ids_2 ? 2'h2 : _GEN_3677; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4702 = 7'h5d == rob_alloc_ids_2 ? 2'h2 : _GEN_3678; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4703 = 7'h5e == rob_alloc_ids_2 ? 2'h2 : _GEN_3679; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4704 = 7'h5f == rob_alloc_ids_2 ? 2'h2 : _GEN_3680; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4705 = 7'h60 == rob_alloc_ids_2 ? 2'h2 : _GEN_3681; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4706 = 7'h61 == rob_alloc_ids_2 ? 2'h2 : _GEN_3682; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4707 = 7'h62 == rob_alloc_ids_2 ? 2'h2 : _GEN_3683; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4708 = 7'h63 == rob_alloc_ids_2 ? 2'h2 : _GEN_3684; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4709 = 7'h64 == rob_alloc_ids_2 ? 2'h2 : _GEN_3685; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4710 = 7'h65 == rob_alloc_ids_2 ? 2'h2 : _GEN_3686; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4711 = 7'h66 == rob_alloc_ids_2 ? 2'h2 : _GEN_3687; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4712 = 7'h67 == rob_alloc_ids_2 ? 2'h2 : _GEN_3688; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4713 = 7'h68 == rob_alloc_ids_2 ? 2'h2 : _GEN_3689; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4714 = 7'h69 == rob_alloc_ids_2 ? 2'h2 : _GEN_3690; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4715 = 7'h6a == rob_alloc_ids_2 ? 2'h2 : _GEN_3691; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4716 = 7'h6b == rob_alloc_ids_2 ? 2'h2 : _GEN_3692; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4717 = 7'h6c == rob_alloc_ids_2 ? 2'h2 : _GEN_3693; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4718 = 7'h6d == rob_alloc_ids_2 ? 2'h2 : _GEN_3694; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4719 = 7'h6e == rob_alloc_ids_2 ? 2'h2 : _GEN_3695; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4720 = 7'h6f == rob_alloc_ids_2 ? 2'h2 : _GEN_3696; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4721 = 7'h70 == rob_alloc_ids_2 ? 2'h2 : _GEN_3697; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4722 = 7'h71 == rob_alloc_ids_2 ? 2'h2 : _GEN_3698; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4723 = 7'h72 == rob_alloc_ids_2 ? 2'h2 : _GEN_3699; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4724 = 7'h73 == rob_alloc_ids_2 ? 2'h2 : _GEN_3700; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4725 = 7'h74 == rob_alloc_ids_2 ? 2'h2 : _GEN_3701; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4726 = 7'h75 == rob_alloc_ids_2 ? 2'h2 : _GEN_3702; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4727 = 7'h76 == rob_alloc_ids_2 ? 2'h2 : _GEN_3703; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4728 = 7'h77 == rob_alloc_ids_2 ? 2'h2 : _GEN_3704; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4729 = 7'h78 == rob_alloc_ids_2 ? 2'h2 : _GEN_3705; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4730 = 7'h79 == rob_alloc_ids_2 ? 2'h2 : _GEN_3706; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4731 = 7'h7a == rob_alloc_ids_2 ? 2'h2 : _GEN_3707; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4732 = 7'h7b == rob_alloc_ids_2 ? 2'h2 : _GEN_3708; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4733 = 7'h7c == rob_alloc_ids_2 ? 2'h2 : _GEN_3709; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4734 = 7'h7d == rob_alloc_ids_2 ? 2'h2 : _GEN_3710; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4735 = 7'h7e == rob_alloc_ids_2 ? 2'h2 : _GEN_3711; // @[TestHarness.scala 181:{36,36}]
  wire [1:0] _GEN_4736 = 7'h7f == rob_alloc_ids_2 ? 2'h2 : _GEN_3712; // @[TestHarness.scala 181:{36,36}]
  wire [3:0] _rob_n_flits_T_55 = igen_2_io_n_flits; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4737 = 7'h0 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3713; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4738 = 7'h1 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3714; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4739 = 7'h2 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3715; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4740 = 7'h3 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3716; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4741 = 7'h4 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3717; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4742 = 7'h5 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3718; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4743 = 7'h6 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3719; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4744 = 7'h7 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3720; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4745 = 7'h8 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3721; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4746 = 7'h9 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3722; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4747 = 7'ha == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3723; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4748 = 7'hb == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3724; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4749 = 7'hc == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3725; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4750 = 7'hd == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3726; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4751 = 7'he == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3727; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4752 = 7'hf == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3728; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4753 = 7'h10 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3729; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4754 = 7'h11 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3730; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4755 = 7'h12 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3731; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4756 = 7'h13 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3732; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4757 = 7'h14 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3733; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4758 = 7'h15 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3734; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4759 = 7'h16 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3735; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4760 = 7'h17 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3736; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4761 = 7'h18 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3737; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4762 = 7'h19 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3738; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4763 = 7'h1a == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3739; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4764 = 7'h1b == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3740; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4765 = 7'h1c == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3741; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4766 = 7'h1d == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3742; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4767 = 7'h1e == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3743; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4768 = 7'h1f == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3744; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4769 = 7'h20 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3745; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4770 = 7'h21 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3746; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4771 = 7'h22 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3747; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4772 = 7'h23 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3748; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4773 = 7'h24 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3749; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4774 = 7'h25 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3750; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4775 = 7'h26 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3751; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4776 = 7'h27 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3752; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4777 = 7'h28 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3753; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4778 = 7'h29 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3754; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4779 = 7'h2a == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3755; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4780 = 7'h2b == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3756; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4781 = 7'h2c == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3757; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4782 = 7'h2d == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3758; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4783 = 7'h2e == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3759; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4784 = 7'h2f == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3760; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4785 = 7'h30 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3761; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4786 = 7'h31 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3762; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4787 = 7'h32 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3763; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4788 = 7'h33 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3764; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4789 = 7'h34 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3765; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4790 = 7'h35 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3766; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4791 = 7'h36 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3767; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4792 = 7'h37 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3768; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4793 = 7'h38 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3769; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4794 = 7'h39 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3770; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4795 = 7'h3a == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3771; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4796 = 7'h3b == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3772; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4797 = 7'h3c == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3773; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4798 = 7'h3d == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3774; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4799 = 7'h3e == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3775; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4800 = 7'h3f == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3776; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4801 = 7'h40 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3777; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4802 = 7'h41 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3778; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4803 = 7'h42 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3779; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4804 = 7'h43 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3780; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4805 = 7'h44 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3781; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4806 = 7'h45 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3782; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4807 = 7'h46 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3783; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4808 = 7'h47 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3784; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4809 = 7'h48 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3785; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4810 = 7'h49 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3786; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4811 = 7'h4a == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3787; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4812 = 7'h4b == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3788; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4813 = 7'h4c == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3789; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4814 = 7'h4d == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3790; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4815 = 7'h4e == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3791; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4816 = 7'h4f == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3792; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4817 = 7'h50 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3793; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4818 = 7'h51 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3794; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4819 = 7'h52 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3795; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4820 = 7'h53 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3796; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4821 = 7'h54 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3797; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4822 = 7'h55 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3798; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4823 = 7'h56 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3799; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4824 = 7'h57 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3800; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4825 = 7'h58 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3801; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4826 = 7'h59 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3802; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4827 = 7'h5a == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3803; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4828 = 7'h5b == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3804; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4829 = 7'h5c == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3805; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4830 = 7'h5d == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3806; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4831 = 7'h5e == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3807; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4832 = 7'h5f == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3808; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4833 = 7'h60 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3809; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4834 = 7'h61 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3810; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4835 = 7'h62 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3811; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4836 = 7'h63 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3812; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4837 = 7'h64 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3813; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4838 = 7'h65 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3814; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4839 = 7'h66 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3815; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4840 = 7'h67 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3816; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4841 = 7'h68 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3817; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4842 = 7'h69 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3818; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4843 = 7'h6a == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3819; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4844 = 7'h6b == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3820; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4845 = 7'h6c == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3821; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4846 = 7'h6d == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3822; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4847 = 7'h6e == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3823; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4848 = 7'h6f == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3824; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4849 = 7'h70 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3825; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4850 = 7'h71 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3826; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4851 = 7'h72 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3827; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4852 = 7'h73 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3828; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4853 = 7'h74 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3829; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4854 = 7'h75 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3830; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4855 = 7'h76 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3831; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4856 = 7'h77 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3832; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4857 = 7'h78 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3833; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4858 = 7'h79 == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3834; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4859 = 7'h7a == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3835; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4860 = 7'h7b == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3836; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4861 = 7'h7c == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3837; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4862 = 7'h7d == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3838; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4863 = 7'h7e == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3839; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4864 = 7'h7f == rob_alloc_ids_2 ? _rob_n_flits_T_55 : _GEN_3840; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_4865 = 7'h0 == rob_alloc_ids_2 ? 4'h0 : _GEN_3841; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4866 = 7'h1 == rob_alloc_ids_2 ? 4'h0 : _GEN_3842; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4867 = 7'h2 == rob_alloc_ids_2 ? 4'h0 : _GEN_3843; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4868 = 7'h3 == rob_alloc_ids_2 ? 4'h0 : _GEN_3844; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4869 = 7'h4 == rob_alloc_ids_2 ? 4'h0 : _GEN_3845; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4870 = 7'h5 == rob_alloc_ids_2 ? 4'h0 : _GEN_3846; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4871 = 7'h6 == rob_alloc_ids_2 ? 4'h0 : _GEN_3847; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4872 = 7'h7 == rob_alloc_ids_2 ? 4'h0 : _GEN_3848; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4873 = 7'h8 == rob_alloc_ids_2 ? 4'h0 : _GEN_3849; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4874 = 7'h9 == rob_alloc_ids_2 ? 4'h0 : _GEN_3850; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4875 = 7'ha == rob_alloc_ids_2 ? 4'h0 : _GEN_3851; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4876 = 7'hb == rob_alloc_ids_2 ? 4'h0 : _GEN_3852; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4877 = 7'hc == rob_alloc_ids_2 ? 4'h0 : _GEN_3853; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4878 = 7'hd == rob_alloc_ids_2 ? 4'h0 : _GEN_3854; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4879 = 7'he == rob_alloc_ids_2 ? 4'h0 : _GEN_3855; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4880 = 7'hf == rob_alloc_ids_2 ? 4'h0 : _GEN_3856; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4881 = 7'h10 == rob_alloc_ids_2 ? 4'h0 : _GEN_3857; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4882 = 7'h11 == rob_alloc_ids_2 ? 4'h0 : _GEN_3858; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4883 = 7'h12 == rob_alloc_ids_2 ? 4'h0 : _GEN_3859; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4884 = 7'h13 == rob_alloc_ids_2 ? 4'h0 : _GEN_3860; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4885 = 7'h14 == rob_alloc_ids_2 ? 4'h0 : _GEN_3861; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4886 = 7'h15 == rob_alloc_ids_2 ? 4'h0 : _GEN_3862; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4887 = 7'h16 == rob_alloc_ids_2 ? 4'h0 : _GEN_3863; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4888 = 7'h17 == rob_alloc_ids_2 ? 4'h0 : _GEN_3864; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4889 = 7'h18 == rob_alloc_ids_2 ? 4'h0 : _GEN_3865; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4890 = 7'h19 == rob_alloc_ids_2 ? 4'h0 : _GEN_3866; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4891 = 7'h1a == rob_alloc_ids_2 ? 4'h0 : _GEN_3867; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4892 = 7'h1b == rob_alloc_ids_2 ? 4'h0 : _GEN_3868; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4893 = 7'h1c == rob_alloc_ids_2 ? 4'h0 : _GEN_3869; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4894 = 7'h1d == rob_alloc_ids_2 ? 4'h0 : _GEN_3870; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4895 = 7'h1e == rob_alloc_ids_2 ? 4'h0 : _GEN_3871; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4896 = 7'h1f == rob_alloc_ids_2 ? 4'h0 : _GEN_3872; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4897 = 7'h20 == rob_alloc_ids_2 ? 4'h0 : _GEN_3873; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4898 = 7'h21 == rob_alloc_ids_2 ? 4'h0 : _GEN_3874; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4899 = 7'h22 == rob_alloc_ids_2 ? 4'h0 : _GEN_3875; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4900 = 7'h23 == rob_alloc_ids_2 ? 4'h0 : _GEN_3876; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4901 = 7'h24 == rob_alloc_ids_2 ? 4'h0 : _GEN_3877; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4902 = 7'h25 == rob_alloc_ids_2 ? 4'h0 : _GEN_3878; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4903 = 7'h26 == rob_alloc_ids_2 ? 4'h0 : _GEN_3879; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4904 = 7'h27 == rob_alloc_ids_2 ? 4'h0 : _GEN_3880; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4905 = 7'h28 == rob_alloc_ids_2 ? 4'h0 : _GEN_3881; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4906 = 7'h29 == rob_alloc_ids_2 ? 4'h0 : _GEN_3882; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4907 = 7'h2a == rob_alloc_ids_2 ? 4'h0 : _GEN_3883; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4908 = 7'h2b == rob_alloc_ids_2 ? 4'h0 : _GEN_3884; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4909 = 7'h2c == rob_alloc_ids_2 ? 4'h0 : _GEN_3885; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4910 = 7'h2d == rob_alloc_ids_2 ? 4'h0 : _GEN_3886; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4911 = 7'h2e == rob_alloc_ids_2 ? 4'h0 : _GEN_3887; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4912 = 7'h2f == rob_alloc_ids_2 ? 4'h0 : _GEN_3888; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4913 = 7'h30 == rob_alloc_ids_2 ? 4'h0 : _GEN_3889; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4914 = 7'h31 == rob_alloc_ids_2 ? 4'h0 : _GEN_3890; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4915 = 7'h32 == rob_alloc_ids_2 ? 4'h0 : _GEN_3891; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4916 = 7'h33 == rob_alloc_ids_2 ? 4'h0 : _GEN_3892; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4917 = 7'h34 == rob_alloc_ids_2 ? 4'h0 : _GEN_3893; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4918 = 7'h35 == rob_alloc_ids_2 ? 4'h0 : _GEN_3894; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4919 = 7'h36 == rob_alloc_ids_2 ? 4'h0 : _GEN_3895; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4920 = 7'h37 == rob_alloc_ids_2 ? 4'h0 : _GEN_3896; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4921 = 7'h38 == rob_alloc_ids_2 ? 4'h0 : _GEN_3897; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4922 = 7'h39 == rob_alloc_ids_2 ? 4'h0 : _GEN_3898; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4923 = 7'h3a == rob_alloc_ids_2 ? 4'h0 : _GEN_3899; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4924 = 7'h3b == rob_alloc_ids_2 ? 4'h0 : _GEN_3900; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4925 = 7'h3c == rob_alloc_ids_2 ? 4'h0 : _GEN_3901; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4926 = 7'h3d == rob_alloc_ids_2 ? 4'h0 : _GEN_3902; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4927 = 7'h3e == rob_alloc_ids_2 ? 4'h0 : _GEN_3903; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4928 = 7'h3f == rob_alloc_ids_2 ? 4'h0 : _GEN_3904; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4929 = 7'h40 == rob_alloc_ids_2 ? 4'h0 : _GEN_3905; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4930 = 7'h41 == rob_alloc_ids_2 ? 4'h0 : _GEN_3906; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4931 = 7'h42 == rob_alloc_ids_2 ? 4'h0 : _GEN_3907; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4932 = 7'h43 == rob_alloc_ids_2 ? 4'h0 : _GEN_3908; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4933 = 7'h44 == rob_alloc_ids_2 ? 4'h0 : _GEN_3909; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4934 = 7'h45 == rob_alloc_ids_2 ? 4'h0 : _GEN_3910; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4935 = 7'h46 == rob_alloc_ids_2 ? 4'h0 : _GEN_3911; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4936 = 7'h47 == rob_alloc_ids_2 ? 4'h0 : _GEN_3912; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4937 = 7'h48 == rob_alloc_ids_2 ? 4'h0 : _GEN_3913; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4938 = 7'h49 == rob_alloc_ids_2 ? 4'h0 : _GEN_3914; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4939 = 7'h4a == rob_alloc_ids_2 ? 4'h0 : _GEN_3915; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4940 = 7'h4b == rob_alloc_ids_2 ? 4'h0 : _GEN_3916; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4941 = 7'h4c == rob_alloc_ids_2 ? 4'h0 : _GEN_3917; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4942 = 7'h4d == rob_alloc_ids_2 ? 4'h0 : _GEN_3918; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4943 = 7'h4e == rob_alloc_ids_2 ? 4'h0 : _GEN_3919; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4944 = 7'h4f == rob_alloc_ids_2 ? 4'h0 : _GEN_3920; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4945 = 7'h50 == rob_alloc_ids_2 ? 4'h0 : _GEN_3921; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4946 = 7'h51 == rob_alloc_ids_2 ? 4'h0 : _GEN_3922; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4947 = 7'h52 == rob_alloc_ids_2 ? 4'h0 : _GEN_3923; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4948 = 7'h53 == rob_alloc_ids_2 ? 4'h0 : _GEN_3924; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4949 = 7'h54 == rob_alloc_ids_2 ? 4'h0 : _GEN_3925; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4950 = 7'h55 == rob_alloc_ids_2 ? 4'h0 : _GEN_3926; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4951 = 7'h56 == rob_alloc_ids_2 ? 4'h0 : _GEN_3927; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4952 = 7'h57 == rob_alloc_ids_2 ? 4'h0 : _GEN_3928; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4953 = 7'h58 == rob_alloc_ids_2 ? 4'h0 : _GEN_3929; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4954 = 7'h59 == rob_alloc_ids_2 ? 4'h0 : _GEN_3930; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4955 = 7'h5a == rob_alloc_ids_2 ? 4'h0 : _GEN_3931; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4956 = 7'h5b == rob_alloc_ids_2 ? 4'h0 : _GEN_3932; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4957 = 7'h5c == rob_alloc_ids_2 ? 4'h0 : _GEN_3933; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4958 = 7'h5d == rob_alloc_ids_2 ? 4'h0 : _GEN_3934; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4959 = 7'h5e == rob_alloc_ids_2 ? 4'h0 : _GEN_3935; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4960 = 7'h5f == rob_alloc_ids_2 ? 4'h0 : _GEN_3936; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4961 = 7'h60 == rob_alloc_ids_2 ? 4'h0 : _GEN_3937; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4962 = 7'h61 == rob_alloc_ids_2 ? 4'h0 : _GEN_3938; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4963 = 7'h62 == rob_alloc_ids_2 ? 4'h0 : _GEN_3939; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4964 = 7'h63 == rob_alloc_ids_2 ? 4'h0 : _GEN_3940; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4965 = 7'h64 == rob_alloc_ids_2 ? 4'h0 : _GEN_3941; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4966 = 7'h65 == rob_alloc_ids_2 ? 4'h0 : _GEN_3942; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4967 = 7'h66 == rob_alloc_ids_2 ? 4'h0 : _GEN_3943; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4968 = 7'h67 == rob_alloc_ids_2 ? 4'h0 : _GEN_3944; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4969 = 7'h68 == rob_alloc_ids_2 ? 4'h0 : _GEN_3945; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4970 = 7'h69 == rob_alloc_ids_2 ? 4'h0 : _GEN_3946; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4971 = 7'h6a == rob_alloc_ids_2 ? 4'h0 : _GEN_3947; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4972 = 7'h6b == rob_alloc_ids_2 ? 4'h0 : _GEN_3948; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4973 = 7'h6c == rob_alloc_ids_2 ? 4'h0 : _GEN_3949; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4974 = 7'h6d == rob_alloc_ids_2 ? 4'h0 : _GEN_3950; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4975 = 7'h6e == rob_alloc_ids_2 ? 4'h0 : _GEN_3951; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4976 = 7'h6f == rob_alloc_ids_2 ? 4'h0 : _GEN_3952; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4977 = 7'h70 == rob_alloc_ids_2 ? 4'h0 : _GEN_3953; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4978 = 7'h71 == rob_alloc_ids_2 ? 4'h0 : _GEN_3954; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4979 = 7'h72 == rob_alloc_ids_2 ? 4'h0 : _GEN_3955; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4980 = 7'h73 == rob_alloc_ids_2 ? 4'h0 : _GEN_3956; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4981 = 7'h74 == rob_alloc_ids_2 ? 4'h0 : _GEN_3957; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4982 = 7'h75 == rob_alloc_ids_2 ? 4'h0 : _GEN_3958; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4983 = 7'h76 == rob_alloc_ids_2 ? 4'h0 : _GEN_3959; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4984 = 7'h77 == rob_alloc_ids_2 ? 4'h0 : _GEN_3960; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4985 = 7'h78 == rob_alloc_ids_2 ? 4'h0 : _GEN_3961; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4986 = 7'h79 == rob_alloc_ids_2 ? 4'h0 : _GEN_3962; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4987 = 7'h7a == rob_alloc_ids_2 ? 4'h0 : _GEN_3963; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4988 = 7'h7b == rob_alloc_ids_2 ? 4'h0 : _GEN_3964; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4989 = 7'h7c == rob_alloc_ids_2 ? 4'h0 : _GEN_3965; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4990 = 7'h7d == rob_alloc_ids_2 ? 4'h0 : _GEN_3966; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4991 = 7'h7e == rob_alloc_ids_2 ? 4'h0 : _GEN_3967; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_4992 = 7'h7f == rob_alloc_ids_2 ? 4'h0 : _GEN_3968; // @[TestHarness.scala 183:{36,36}]
  wire [63:0] _GEN_4993 = 7'h0 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_3969; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_4994 = 7'h1 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_3970; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_4995 = 7'h2 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_3971; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_4996 = 7'h3 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_3972; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_4997 = 7'h4 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_3973; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_4998 = 7'h5 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_3974; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_4999 = 7'h6 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_3975; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5000 = 7'h7 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_3976; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5001 = 7'h8 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_3977; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5002 = 7'h9 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_3978; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5003 = 7'ha == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_3979; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5004 = 7'hb == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_3980; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5005 = 7'hc == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_3981; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5006 = 7'hd == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_3982; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5007 = 7'he == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_3983; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5008 = 7'hf == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_3984; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5009 = 7'h10 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_3985; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5010 = 7'h11 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_3986; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5011 = 7'h12 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_3987; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5012 = 7'h13 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_3988; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5013 = 7'h14 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_3989; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5014 = 7'h15 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_3990; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5015 = 7'h16 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_3991; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5016 = 7'h17 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_3992; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5017 = 7'h18 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_3993; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5018 = 7'h19 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_3994; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5019 = 7'h1a == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_3995; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5020 = 7'h1b == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_3996; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5021 = 7'h1c == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_3997; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5022 = 7'h1d == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_3998; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5023 = 7'h1e == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_3999; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5024 = 7'h1f == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4000; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5025 = 7'h20 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4001; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5026 = 7'h21 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4002; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5027 = 7'h22 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4003; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5028 = 7'h23 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4004; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5029 = 7'h24 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4005; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5030 = 7'h25 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4006; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5031 = 7'h26 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4007; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5032 = 7'h27 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4008; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5033 = 7'h28 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4009; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5034 = 7'h29 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4010; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5035 = 7'h2a == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4011; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5036 = 7'h2b == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4012; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5037 = 7'h2c == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4013; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5038 = 7'h2d == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4014; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5039 = 7'h2e == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4015; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5040 = 7'h2f == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4016; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5041 = 7'h30 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4017; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5042 = 7'h31 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4018; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5043 = 7'h32 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4019; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5044 = 7'h33 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4020; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5045 = 7'h34 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4021; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5046 = 7'h35 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4022; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5047 = 7'h36 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4023; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5048 = 7'h37 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4024; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5049 = 7'h38 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4025; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5050 = 7'h39 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4026; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5051 = 7'h3a == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4027; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5052 = 7'h3b == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4028; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5053 = 7'h3c == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4029; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5054 = 7'h3d == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4030; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5055 = 7'h3e == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4031; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5056 = 7'h3f == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4032; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5057 = 7'h40 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4033; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5058 = 7'h41 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4034; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5059 = 7'h42 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4035; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5060 = 7'h43 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4036; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5061 = 7'h44 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4037; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5062 = 7'h45 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4038; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5063 = 7'h46 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4039; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5064 = 7'h47 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4040; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5065 = 7'h48 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4041; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5066 = 7'h49 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4042; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5067 = 7'h4a == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4043; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5068 = 7'h4b == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4044; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5069 = 7'h4c == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4045; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5070 = 7'h4d == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4046; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5071 = 7'h4e == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4047; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5072 = 7'h4f == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4048; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5073 = 7'h50 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4049; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5074 = 7'h51 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4050; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5075 = 7'h52 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4051; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5076 = 7'h53 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4052; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5077 = 7'h54 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4053; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5078 = 7'h55 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4054; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5079 = 7'h56 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4055; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5080 = 7'h57 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4056; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5081 = 7'h58 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4057; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5082 = 7'h59 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4058; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5083 = 7'h5a == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4059; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5084 = 7'h5b == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4060; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5085 = 7'h5c == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4061; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5086 = 7'h5d == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4062; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5087 = 7'h5e == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4063; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5088 = 7'h5f == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4064; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5089 = 7'h60 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4065; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5090 = 7'h61 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4066; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5091 = 7'h62 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4067; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5092 = 7'h63 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4068; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5093 = 7'h64 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4069; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5094 = 7'h65 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4070; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5095 = 7'h66 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4071; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5096 = 7'h67 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4072; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5097 = 7'h68 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4073; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5098 = 7'h69 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4074; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5099 = 7'h6a == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4075; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5100 = 7'h6b == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4076; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5101 = 7'h6c == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4077; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5102 = 7'h6d == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4078; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5103 = 7'h6e == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4079; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5104 = 7'h6f == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4080; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5105 = 7'h70 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4081; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5106 = 7'h71 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4082; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5107 = 7'h72 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4083; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5108 = 7'h73 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4084; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5109 = 7'h74 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4085; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5110 = 7'h75 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4086; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5111 = 7'h76 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4087; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5112 = 7'h77 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4088; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5113 = 7'h78 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4089; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5114 = 7'h79 == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4090; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5115 = 7'h7a == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4091; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5116 = 7'h7b == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4092; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5117 = 7'h7c == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4093; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5118 = 7'h7d == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4094; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5119 = 7'h7e == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4095; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_5120 = 7'h7f == rob_alloc_ids_2 ? _rob_tscs_T_31 : _GEN_4096; // @[TestHarness.scala 184:{36,36}]
  wire [31:0] _GEN_5121 = igen_2_io_fire ? _GEN_4097 : _GEN_3073; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5122 = igen_2_io_fire ? _GEN_4098 : _GEN_3074; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5123 = igen_2_io_fire ? _GEN_4099 : _GEN_3075; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5124 = igen_2_io_fire ? _GEN_4100 : _GEN_3076; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5125 = igen_2_io_fire ? _GEN_4101 : _GEN_3077; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5126 = igen_2_io_fire ? _GEN_4102 : _GEN_3078; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5127 = igen_2_io_fire ? _GEN_4103 : _GEN_3079; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5128 = igen_2_io_fire ? _GEN_4104 : _GEN_3080; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5129 = igen_2_io_fire ? _GEN_4105 : _GEN_3081; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5130 = igen_2_io_fire ? _GEN_4106 : _GEN_3082; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5131 = igen_2_io_fire ? _GEN_4107 : _GEN_3083; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5132 = igen_2_io_fire ? _GEN_4108 : _GEN_3084; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5133 = igen_2_io_fire ? _GEN_4109 : _GEN_3085; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5134 = igen_2_io_fire ? _GEN_4110 : _GEN_3086; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5135 = igen_2_io_fire ? _GEN_4111 : _GEN_3087; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5136 = igen_2_io_fire ? _GEN_4112 : _GEN_3088; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5137 = igen_2_io_fire ? _GEN_4113 : _GEN_3089; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5138 = igen_2_io_fire ? _GEN_4114 : _GEN_3090; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5139 = igen_2_io_fire ? _GEN_4115 : _GEN_3091; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5140 = igen_2_io_fire ? _GEN_4116 : _GEN_3092; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5141 = igen_2_io_fire ? _GEN_4117 : _GEN_3093; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5142 = igen_2_io_fire ? _GEN_4118 : _GEN_3094; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5143 = igen_2_io_fire ? _GEN_4119 : _GEN_3095; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5144 = igen_2_io_fire ? _GEN_4120 : _GEN_3096; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5145 = igen_2_io_fire ? _GEN_4121 : _GEN_3097; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5146 = igen_2_io_fire ? _GEN_4122 : _GEN_3098; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5147 = igen_2_io_fire ? _GEN_4123 : _GEN_3099; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5148 = igen_2_io_fire ? _GEN_4124 : _GEN_3100; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5149 = igen_2_io_fire ? _GEN_4125 : _GEN_3101; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5150 = igen_2_io_fire ? _GEN_4126 : _GEN_3102; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5151 = igen_2_io_fire ? _GEN_4127 : _GEN_3103; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5152 = igen_2_io_fire ? _GEN_4128 : _GEN_3104; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5153 = igen_2_io_fire ? _GEN_4129 : _GEN_3105; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5154 = igen_2_io_fire ? _GEN_4130 : _GEN_3106; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5155 = igen_2_io_fire ? _GEN_4131 : _GEN_3107; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5156 = igen_2_io_fire ? _GEN_4132 : _GEN_3108; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5157 = igen_2_io_fire ? _GEN_4133 : _GEN_3109; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5158 = igen_2_io_fire ? _GEN_4134 : _GEN_3110; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5159 = igen_2_io_fire ? _GEN_4135 : _GEN_3111; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5160 = igen_2_io_fire ? _GEN_4136 : _GEN_3112; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5161 = igen_2_io_fire ? _GEN_4137 : _GEN_3113; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5162 = igen_2_io_fire ? _GEN_4138 : _GEN_3114; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5163 = igen_2_io_fire ? _GEN_4139 : _GEN_3115; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5164 = igen_2_io_fire ? _GEN_4140 : _GEN_3116; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5165 = igen_2_io_fire ? _GEN_4141 : _GEN_3117; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5166 = igen_2_io_fire ? _GEN_4142 : _GEN_3118; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5167 = igen_2_io_fire ? _GEN_4143 : _GEN_3119; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5168 = igen_2_io_fire ? _GEN_4144 : _GEN_3120; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5169 = igen_2_io_fire ? _GEN_4145 : _GEN_3121; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5170 = igen_2_io_fire ? _GEN_4146 : _GEN_3122; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5171 = igen_2_io_fire ? _GEN_4147 : _GEN_3123; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5172 = igen_2_io_fire ? _GEN_4148 : _GEN_3124; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5173 = igen_2_io_fire ? _GEN_4149 : _GEN_3125; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5174 = igen_2_io_fire ? _GEN_4150 : _GEN_3126; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5175 = igen_2_io_fire ? _GEN_4151 : _GEN_3127; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5176 = igen_2_io_fire ? _GEN_4152 : _GEN_3128; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5177 = igen_2_io_fire ? _GEN_4153 : _GEN_3129; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5178 = igen_2_io_fire ? _GEN_4154 : _GEN_3130; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5179 = igen_2_io_fire ? _GEN_4155 : _GEN_3131; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5180 = igen_2_io_fire ? _GEN_4156 : _GEN_3132; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5181 = igen_2_io_fire ? _GEN_4157 : _GEN_3133; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5182 = igen_2_io_fire ? _GEN_4158 : _GEN_3134; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5183 = igen_2_io_fire ? _GEN_4159 : _GEN_3135; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5184 = igen_2_io_fire ? _GEN_4160 : _GEN_3136; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5185 = igen_2_io_fire ? _GEN_4161 : _GEN_3137; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5186 = igen_2_io_fire ? _GEN_4162 : _GEN_3138; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5187 = igen_2_io_fire ? _GEN_4163 : _GEN_3139; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5188 = igen_2_io_fire ? _GEN_4164 : _GEN_3140; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5189 = igen_2_io_fire ? _GEN_4165 : _GEN_3141; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5190 = igen_2_io_fire ? _GEN_4166 : _GEN_3142; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5191 = igen_2_io_fire ? _GEN_4167 : _GEN_3143; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5192 = igen_2_io_fire ? _GEN_4168 : _GEN_3144; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5193 = igen_2_io_fire ? _GEN_4169 : _GEN_3145; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5194 = igen_2_io_fire ? _GEN_4170 : _GEN_3146; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5195 = igen_2_io_fire ? _GEN_4171 : _GEN_3147; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5196 = igen_2_io_fire ? _GEN_4172 : _GEN_3148; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5197 = igen_2_io_fire ? _GEN_4173 : _GEN_3149; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5198 = igen_2_io_fire ? _GEN_4174 : _GEN_3150; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5199 = igen_2_io_fire ? _GEN_4175 : _GEN_3151; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5200 = igen_2_io_fire ? _GEN_4176 : _GEN_3152; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5201 = igen_2_io_fire ? _GEN_4177 : _GEN_3153; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5202 = igen_2_io_fire ? _GEN_4178 : _GEN_3154; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5203 = igen_2_io_fire ? _GEN_4179 : _GEN_3155; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5204 = igen_2_io_fire ? _GEN_4180 : _GEN_3156; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5205 = igen_2_io_fire ? _GEN_4181 : _GEN_3157; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5206 = igen_2_io_fire ? _GEN_4182 : _GEN_3158; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5207 = igen_2_io_fire ? _GEN_4183 : _GEN_3159; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5208 = igen_2_io_fire ? _GEN_4184 : _GEN_3160; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5209 = igen_2_io_fire ? _GEN_4185 : _GEN_3161; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5210 = igen_2_io_fire ? _GEN_4186 : _GEN_3162; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5211 = igen_2_io_fire ? _GEN_4187 : _GEN_3163; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5212 = igen_2_io_fire ? _GEN_4188 : _GEN_3164; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5213 = igen_2_io_fire ? _GEN_4189 : _GEN_3165; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5214 = igen_2_io_fire ? _GEN_4190 : _GEN_3166; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5215 = igen_2_io_fire ? _GEN_4191 : _GEN_3167; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5216 = igen_2_io_fire ? _GEN_4192 : _GEN_3168; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5217 = igen_2_io_fire ? _GEN_4193 : _GEN_3169; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5218 = igen_2_io_fire ? _GEN_4194 : _GEN_3170; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5219 = igen_2_io_fire ? _GEN_4195 : _GEN_3171; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5220 = igen_2_io_fire ? _GEN_4196 : _GEN_3172; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5221 = igen_2_io_fire ? _GEN_4197 : _GEN_3173; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5222 = igen_2_io_fire ? _GEN_4198 : _GEN_3174; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5223 = igen_2_io_fire ? _GEN_4199 : _GEN_3175; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5224 = igen_2_io_fire ? _GEN_4200 : _GEN_3176; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5225 = igen_2_io_fire ? _GEN_4201 : _GEN_3177; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5226 = igen_2_io_fire ? _GEN_4202 : _GEN_3178; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5227 = igen_2_io_fire ? _GEN_4203 : _GEN_3179; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5228 = igen_2_io_fire ? _GEN_4204 : _GEN_3180; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5229 = igen_2_io_fire ? _GEN_4205 : _GEN_3181; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5230 = igen_2_io_fire ? _GEN_4206 : _GEN_3182; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5231 = igen_2_io_fire ? _GEN_4207 : _GEN_3183; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5232 = igen_2_io_fire ? _GEN_4208 : _GEN_3184; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5233 = igen_2_io_fire ? _GEN_4209 : _GEN_3185; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5234 = igen_2_io_fire ? _GEN_4210 : _GEN_3186; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5235 = igen_2_io_fire ? _GEN_4211 : _GEN_3187; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5236 = igen_2_io_fire ? _GEN_4212 : _GEN_3188; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5237 = igen_2_io_fire ? _GEN_4213 : _GEN_3189; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5238 = igen_2_io_fire ? _GEN_4214 : _GEN_3190; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5239 = igen_2_io_fire ? _GEN_4215 : _GEN_3191; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5240 = igen_2_io_fire ? _GEN_4216 : _GEN_3192; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5241 = igen_2_io_fire ? _GEN_4217 : _GEN_3193; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5242 = igen_2_io_fire ? _GEN_4218 : _GEN_3194; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5243 = igen_2_io_fire ? _GEN_4219 : _GEN_3195; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5244 = igen_2_io_fire ? _GEN_4220 : _GEN_3196; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5245 = igen_2_io_fire ? _GEN_4221 : _GEN_3197; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5246 = igen_2_io_fire ? _GEN_4222 : _GEN_3198; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5247 = igen_2_io_fire ? _GEN_4223 : _GEN_3199; // @[TestHarness.scala 178:25]
  wire [31:0] _GEN_5248 = igen_2_io_fire ? _GEN_4224 : _GEN_3200; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5249 = igen_2_io_fire ? _GEN_4225 : _GEN_3201; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5250 = igen_2_io_fire ? _GEN_4226 : _GEN_3202; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5251 = igen_2_io_fire ? _GEN_4227 : _GEN_3203; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5252 = igen_2_io_fire ? _GEN_4228 : _GEN_3204; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5253 = igen_2_io_fire ? _GEN_4229 : _GEN_3205; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5254 = igen_2_io_fire ? _GEN_4230 : _GEN_3206; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5255 = igen_2_io_fire ? _GEN_4231 : _GEN_3207; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5256 = igen_2_io_fire ? _GEN_4232 : _GEN_3208; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5257 = igen_2_io_fire ? _GEN_4233 : _GEN_3209; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5258 = igen_2_io_fire ? _GEN_4234 : _GEN_3210; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5259 = igen_2_io_fire ? _GEN_4235 : _GEN_3211; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5260 = igen_2_io_fire ? _GEN_4236 : _GEN_3212; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5261 = igen_2_io_fire ? _GEN_4237 : _GEN_3213; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5262 = igen_2_io_fire ? _GEN_4238 : _GEN_3214; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5263 = igen_2_io_fire ? _GEN_4239 : _GEN_3215; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5264 = igen_2_io_fire ? _GEN_4240 : _GEN_3216; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5265 = igen_2_io_fire ? _GEN_4241 : _GEN_3217; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5266 = igen_2_io_fire ? _GEN_4242 : _GEN_3218; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5267 = igen_2_io_fire ? _GEN_4243 : _GEN_3219; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5268 = igen_2_io_fire ? _GEN_4244 : _GEN_3220; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5269 = igen_2_io_fire ? _GEN_4245 : _GEN_3221; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5270 = igen_2_io_fire ? _GEN_4246 : _GEN_3222; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5271 = igen_2_io_fire ? _GEN_4247 : _GEN_3223; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5272 = igen_2_io_fire ? _GEN_4248 : _GEN_3224; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5273 = igen_2_io_fire ? _GEN_4249 : _GEN_3225; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5274 = igen_2_io_fire ? _GEN_4250 : _GEN_3226; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5275 = igen_2_io_fire ? _GEN_4251 : _GEN_3227; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5276 = igen_2_io_fire ? _GEN_4252 : _GEN_3228; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5277 = igen_2_io_fire ? _GEN_4253 : _GEN_3229; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5278 = igen_2_io_fire ? _GEN_4254 : _GEN_3230; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5279 = igen_2_io_fire ? _GEN_4255 : _GEN_3231; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5280 = igen_2_io_fire ? _GEN_4256 : _GEN_3232; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5281 = igen_2_io_fire ? _GEN_4257 : _GEN_3233; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5282 = igen_2_io_fire ? _GEN_4258 : _GEN_3234; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5283 = igen_2_io_fire ? _GEN_4259 : _GEN_3235; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5284 = igen_2_io_fire ? _GEN_4260 : _GEN_3236; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5285 = igen_2_io_fire ? _GEN_4261 : _GEN_3237; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5286 = igen_2_io_fire ? _GEN_4262 : _GEN_3238; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5287 = igen_2_io_fire ? _GEN_4263 : _GEN_3239; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5288 = igen_2_io_fire ? _GEN_4264 : _GEN_3240; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5289 = igen_2_io_fire ? _GEN_4265 : _GEN_3241; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5290 = igen_2_io_fire ? _GEN_4266 : _GEN_3242; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5291 = igen_2_io_fire ? _GEN_4267 : _GEN_3243; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5292 = igen_2_io_fire ? _GEN_4268 : _GEN_3244; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5293 = igen_2_io_fire ? _GEN_4269 : _GEN_3245; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5294 = igen_2_io_fire ? _GEN_4270 : _GEN_3246; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5295 = igen_2_io_fire ? _GEN_4271 : _GEN_3247; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5296 = igen_2_io_fire ? _GEN_4272 : _GEN_3248; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5297 = igen_2_io_fire ? _GEN_4273 : _GEN_3249; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5298 = igen_2_io_fire ? _GEN_4274 : _GEN_3250; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5299 = igen_2_io_fire ? _GEN_4275 : _GEN_3251; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5300 = igen_2_io_fire ? _GEN_4276 : _GEN_3252; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5301 = igen_2_io_fire ? _GEN_4277 : _GEN_3253; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5302 = igen_2_io_fire ? _GEN_4278 : _GEN_3254; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5303 = igen_2_io_fire ? _GEN_4279 : _GEN_3255; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5304 = igen_2_io_fire ? _GEN_4280 : _GEN_3256; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5305 = igen_2_io_fire ? _GEN_4281 : _GEN_3257; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5306 = igen_2_io_fire ? _GEN_4282 : _GEN_3258; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5307 = igen_2_io_fire ? _GEN_4283 : _GEN_3259; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5308 = igen_2_io_fire ? _GEN_4284 : _GEN_3260; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5309 = igen_2_io_fire ? _GEN_4285 : _GEN_3261; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5310 = igen_2_io_fire ? _GEN_4286 : _GEN_3262; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5311 = igen_2_io_fire ? _GEN_4287 : _GEN_3263; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5312 = igen_2_io_fire ? _GEN_4288 : _GEN_3264; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5313 = igen_2_io_fire ? _GEN_4289 : _GEN_3265; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5314 = igen_2_io_fire ? _GEN_4290 : _GEN_3266; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5315 = igen_2_io_fire ? _GEN_4291 : _GEN_3267; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5316 = igen_2_io_fire ? _GEN_4292 : _GEN_3268; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5317 = igen_2_io_fire ? _GEN_4293 : _GEN_3269; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5318 = igen_2_io_fire ? _GEN_4294 : _GEN_3270; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5319 = igen_2_io_fire ? _GEN_4295 : _GEN_3271; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5320 = igen_2_io_fire ? _GEN_4296 : _GEN_3272; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5321 = igen_2_io_fire ? _GEN_4297 : _GEN_3273; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5322 = igen_2_io_fire ? _GEN_4298 : _GEN_3274; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5323 = igen_2_io_fire ? _GEN_4299 : _GEN_3275; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5324 = igen_2_io_fire ? _GEN_4300 : _GEN_3276; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5325 = igen_2_io_fire ? _GEN_4301 : _GEN_3277; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5326 = igen_2_io_fire ? _GEN_4302 : _GEN_3278; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5327 = igen_2_io_fire ? _GEN_4303 : _GEN_3279; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5328 = igen_2_io_fire ? _GEN_4304 : _GEN_3280; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5329 = igen_2_io_fire ? _GEN_4305 : _GEN_3281; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5330 = igen_2_io_fire ? _GEN_4306 : _GEN_3282; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5331 = igen_2_io_fire ? _GEN_4307 : _GEN_3283; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5332 = igen_2_io_fire ? _GEN_4308 : _GEN_3284; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5333 = igen_2_io_fire ? _GEN_4309 : _GEN_3285; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5334 = igen_2_io_fire ? _GEN_4310 : _GEN_3286; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5335 = igen_2_io_fire ? _GEN_4311 : _GEN_3287; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5336 = igen_2_io_fire ? _GEN_4312 : _GEN_3288; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5337 = igen_2_io_fire ? _GEN_4313 : _GEN_3289; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5338 = igen_2_io_fire ? _GEN_4314 : _GEN_3290; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5339 = igen_2_io_fire ? _GEN_4315 : _GEN_3291; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5340 = igen_2_io_fire ? _GEN_4316 : _GEN_3292; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5341 = igen_2_io_fire ? _GEN_4317 : _GEN_3293; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5342 = igen_2_io_fire ? _GEN_4318 : _GEN_3294; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5343 = igen_2_io_fire ? _GEN_4319 : _GEN_3295; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5344 = igen_2_io_fire ? _GEN_4320 : _GEN_3296; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5345 = igen_2_io_fire ? _GEN_4321 : _GEN_3297; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5346 = igen_2_io_fire ? _GEN_4322 : _GEN_3298; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5347 = igen_2_io_fire ? _GEN_4323 : _GEN_3299; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5348 = igen_2_io_fire ? _GEN_4324 : _GEN_3300; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5349 = igen_2_io_fire ? _GEN_4325 : _GEN_3301; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5350 = igen_2_io_fire ? _GEN_4326 : _GEN_3302; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5351 = igen_2_io_fire ? _GEN_4327 : _GEN_3303; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5352 = igen_2_io_fire ? _GEN_4328 : _GEN_3304; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5353 = igen_2_io_fire ? _GEN_4329 : _GEN_3305; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5354 = igen_2_io_fire ? _GEN_4330 : _GEN_3306; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5355 = igen_2_io_fire ? _GEN_4331 : _GEN_3307; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5356 = igen_2_io_fire ? _GEN_4332 : _GEN_3308; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5357 = igen_2_io_fire ? _GEN_4333 : _GEN_3309; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5358 = igen_2_io_fire ? _GEN_4334 : _GEN_3310; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5359 = igen_2_io_fire ? _GEN_4335 : _GEN_3311; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5360 = igen_2_io_fire ? _GEN_4336 : _GEN_3312; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5361 = igen_2_io_fire ? _GEN_4337 : _GEN_3313; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5362 = igen_2_io_fire ? _GEN_4338 : _GEN_3314; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5363 = igen_2_io_fire ? _GEN_4339 : _GEN_3315; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5364 = igen_2_io_fire ? _GEN_4340 : _GEN_3316; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5365 = igen_2_io_fire ? _GEN_4341 : _GEN_3317; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5366 = igen_2_io_fire ? _GEN_4342 : _GEN_3318; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5367 = igen_2_io_fire ? _GEN_4343 : _GEN_3319; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5368 = igen_2_io_fire ? _GEN_4344 : _GEN_3320; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5369 = igen_2_io_fire ? _GEN_4345 : _GEN_3321; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5370 = igen_2_io_fire ? _GEN_4346 : _GEN_3322; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5371 = igen_2_io_fire ? _GEN_4347 : _GEN_3323; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5372 = igen_2_io_fire ? _GEN_4348 : _GEN_3324; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5373 = igen_2_io_fire ? _GEN_4349 : _GEN_3325; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5374 = igen_2_io_fire ? _GEN_4350 : _GEN_3326; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5375 = igen_2_io_fire ? _GEN_4351 : _GEN_3327; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5376 = igen_2_io_fire ? _GEN_4352 : _GEN_3328; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5377 = igen_2_io_fire ? _GEN_4353 : _GEN_3329; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5378 = igen_2_io_fire ? _GEN_4354 : _GEN_3330; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5379 = igen_2_io_fire ? _GEN_4355 : _GEN_3331; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5380 = igen_2_io_fire ? _GEN_4356 : _GEN_3332; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5381 = igen_2_io_fire ? _GEN_4357 : _GEN_3333; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5382 = igen_2_io_fire ? _GEN_4358 : _GEN_3334; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5383 = igen_2_io_fire ? _GEN_4359 : _GEN_3335; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5384 = igen_2_io_fire ? _GEN_4360 : _GEN_3336; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5385 = igen_2_io_fire ? _GEN_4361 : _GEN_3337; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5386 = igen_2_io_fire ? _GEN_4362 : _GEN_3338; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5387 = igen_2_io_fire ? _GEN_4363 : _GEN_3339; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5388 = igen_2_io_fire ? _GEN_4364 : _GEN_3340; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5389 = igen_2_io_fire ? _GEN_4365 : _GEN_3341; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5390 = igen_2_io_fire ? _GEN_4366 : _GEN_3342; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5391 = igen_2_io_fire ? _GEN_4367 : _GEN_3343; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5392 = igen_2_io_fire ? _GEN_4368 : _GEN_3344; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5393 = igen_2_io_fire ? _GEN_4369 : _GEN_3345; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5394 = igen_2_io_fire ? _GEN_4370 : _GEN_3346; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5395 = igen_2_io_fire ? _GEN_4371 : _GEN_3347; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5396 = igen_2_io_fire ? _GEN_4372 : _GEN_3348; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5397 = igen_2_io_fire ? _GEN_4373 : _GEN_3349; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5398 = igen_2_io_fire ? _GEN_4374 : _GEN_3350; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5399 = igen_2_io_fire ? _GEN_4375 : _GEN_3351; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5400 = igen_2_io_fire ? _GEN_4376 : _GEN_3352; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5401 = igen_2_io_fire ? _GEN_4377 : _GEN_3353; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5402 = igen_2_io_fire ? _GEN_4378 : _GEN_3354; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5403 = igen_2_io_fire ? _GEN_4379 : _GEN_3355; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5404 = igen_2_io_fire ? _GEN_4380 : _GEN_3356; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5405 = igen_2_io_fire ? _GEN_4381 : _GEN_3357; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5406 = igen_2_io_fire ? _GEN_4382 : _GEN_3358; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5407 = igen_2_io_fire ? _GEN_4383 : _GEN_3359; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5408 = igen_2_io_fire ? _GEN_4384 : _GEN_3360; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5409 = igen_2_io_fire ? _GEN_4385 : _GEN_3361; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5410 = igen_2_io_fire ? _GEN_4386 : _GEN_3362; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5411 = igen_2_io_fire ? _GEN_4387 : _GEN_3363; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5412 = igen_2_io_fire ? _GEN_4388 : _GEN_3364; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5413 = igen_2_io_fire ? _GEN_4389 : _GEN_3365; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5414 = igen_2_io_fire ? _GEN_4390 : _GEN_3366; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5415 = igen_2_io_fire ? _GEN_4391 : _GEN_3367; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5416 = igen_2_io_fire ? _GEN_4392 : _GEN_3368; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5417 = igen_2_io_fire ? _GEN_4393 : _GEN_3369; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5418 = igen_2_io_fire ? _GEN_4394 : _GEN_3370; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5419 = igen_2_io_fire ? _GEN_4395 : _GEN_3371; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5420 = igen_2_io_fire ? _GEN_4396 : _GEN_3372; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5421 = igen_2_io_fire ? _GEN_4397 : _GEN_3373; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5422 = igen_2_io_fire ? _GEN_4398 : _GEN_3374; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5423 = igen_2_io_fire ? _GEN_4399 : _GEN_3375; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5424 = igen_2_io_fire ? _GEN_4400 : _GEN_3376; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5425 = igen_2_io_fire ? _GEN_4401 : _GEN_3377; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5426 = igen_2_io_fire ? _GEN_4402 : _GEN_3378; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5427 = igen_2_io_fire ? _GEN_4403 : _GEN_3379; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5428 = igen_2_io_fire ? _GEN_4404 : _GEN_3380; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5429 = igen_2_io_fire ? _GEN_4405 : _GEN_3381; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5430 = igen_2_io_fire ? _GEN_4406 : _GEN_3382; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5431 = igen_2_io_fire ? _GEN_4407 : _GEN_3383; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5432 = igen_2_io_fire ? _GEN_4408 : _GEN_3384; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5433 = igen_2_io_fire ? _GEN_4409 : _GEN_3385; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5434 = igen_2_io_fire ? _GEN_4410 : _GEN_3386; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5435 = igen_2_io_fire ? _GEN_4411 : _GEN_3387; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5436 = igen_2_io_fire ? _GEN_4412 : _GEN_3388; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5437 = igen_2_io_fire ? _GEN_4413 : _GEN_3389; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5438 = igen_2_io_fire ? _GEN_4414 : _GEN_3390; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5439 = igen_2_io_fire ? _GEN_4415 : _GEN_3391; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5440 = igen_2_io_fire ? _GEN_4416 : _GEN_3392; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5441 = igen_2_io_fire ? _GEN_4417 : _GEN_3393; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5442 = igen_2_io_fire ? _GEN_4418 : _GEN_3394; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5443 = igen_2_io_fire ? _GEN_4419 : _GEN_3395; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5444 = igen_2_io_fire ? _GEN_4420 : _GEN_3396; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5445 = igen_2_io_fire ? _GEN_4421 : _GEN_3397; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5446 = igen_2_io_fire ? _GEN_4422 : _GEN_3398; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5447 = igen_2_io_fire ? _GEN_4423 : _GEN_3399; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5448 = igen_2_io_fire ? _GEN_4424 : _GEN_3400; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5449 = igen_2_io_fire ? _GEN_4425 : _GEN_3401; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5450 = igen_2_io_fire ? _GEN_4426 : _GEN_3402; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5451 = igen_2_io_fire ? _GEN_4427 : _GEN_3403; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5452 = igen_2_io_fire ? _GEN_4428 : _GEN_3404; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5453 = igen_2_io_fire ? _GEN_4429 : _GEN_3405; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5454 = igen_2_io_fire ? _GEN_4430 : _GEN_3406; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5455 = igen_2_io_fire ? _GEN_4431 : _GEN_3407; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5456 = igen_2_io_fire ? _GEN_4432 : _GEN_3408; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5457 = igen_2_io_fire ? _GEN_4433 : _GEN_3409; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5458 = igen_2_io_fire ? _GEN_4434 : _GEN_3410; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5459 = igen_2_io_fire ? _GEN_4435 : _GEN_3411; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5460 = igen_2_io_fire ? _GEN_4436 : _GEN_3412; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5461 = igen_2_io_fire ? _GEN_4437 : _GEN_3413; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5462 = igen_2_io_fire ? _GEN_4438 : _GEN_3414; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5463 = igen_2_io_fire ? _GEN_4439 : _GEN_3415; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5464 = igen_2_io_fire ? _GEN_4440 : _GEN_3416; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5465 = igen_2_io_fire ? _GEN_4441 : _GEN_3417; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5466 = igen_2_io_fire ? _GEN_4442 : _GEN_3418; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5467 = igen_2_io_fire ? _GEN_4443 : _GEN_3419; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5468 = igen_2_io_fire ? _GEN_4444 : _GEN_3420; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5469 = igen_2_io_fire ? _GEN_4445 : _GEN_3421; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5470 = igen_2_io_fire ? _GEN_4446 : _GEN_3422; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5471 = igen_2_io_fire ? _GEN_4447 : _GEN_3423; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5472 = igen_2_io_fire ? _GEN_4448 : _GEN_3424; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5473 = igen_2_io_fire ? _GEN_4449 : _GEN_3425; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5474 = igen_2_io_fire ? _GEN_4450 : _GEN_3426; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5475 = igen_2_io_fire ? _GEN_4451 : _GEN_3427; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5476 = igen_2_io_fire ? _GEN_4452 : _GEN_3428; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5477 = igen_2_io_fire ? _GEN_4453 : _GEN_3429; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5478 = igen_2_io_fire ? _GEN_4454 : _GEN_3430; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5479 = igen_2_io_fire ? _GEN_4455 : _GEN_3431; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5480 = igen_2_io_fire ? _GEN_4456 : _GEN_3432; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5481 = igen_2_io_fire ? _GEN_4457 : _GEN_3433; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5482 = igen_2_io_fire ? _GEN_4458 : _GEN_3434; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5483 = igen_2_io_fire ? _GEN_4459 : _GEN_3435; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5484 = igen_2_io_fire ? _GEN_4460 : _GEN_3436; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5485 = igen_2_io_fire ? _GEN_4461 : _GEN_3437; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5486 = igen_2_io_fire ? _GEN_4462 : _GEN_3438; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5487 = igen_2_io_fire ? _GEN_4463 : _GEN_3439; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5488 = igen_2_io_fire ? _GEN_4464 : _GEN_3440; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5489 = igen_2_io_fire ? _GEN_4465 : _GEN_3441; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5490 = igen_2_io_fire ? _GEN_4466 : _GEN_3442; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5491 = igen_2_io_fire ? _GEN_4467 : _GEN_3443; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5492 = igen_2_io_fire ? _GEN_4468 : _GEN_3444; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5493 = igen_2_io_fire ? _GEN_4469 : _GEN_3445; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5494 = igen_2_io_fire ? _GEN_4470 : _GEN_3446; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5495 = igen_2_io_fire ? _GEN_4471 : _GEN_3447; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5496 = igen_2_io_fire ? _GEN_4472 : _GEN_3448; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5497 = igen_2_io_fire ? _GEN_4473 : _GEN_3449; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5498 = igen_2_io_fire ? _GEN_4474 : _GEN_3450; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5499 = igen_2_io_fire ? _GEN_4475 : _GEN_3451; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5500 = igen_2_io_fire ? _GEN_4476 : _GEN_3452; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5501 = igen_2_io_fire ? _GEN_4477 : _GEN_3453; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5502 = igen_2_io_fire ? _GEN_4478 : _GEN_3454; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5503 = igen_2_io_fire ? _GEN_4479 : _GEN_3455; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_5504 = igen_2_io_fire ? _GEN_4480 : _GEN_3456; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5505 = igen_2_io_fire ? _GEN_4481 : _GEN_3457; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5506 = igen_2_io_fire ? _GEN_4482 : _GEN_3458; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5507 = igen_2_io_fire ? _GEN_4483 : _GEN_3459; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5508 = igen_2_io_fire ? _GEN_4484 : _GEN_3460; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5509 = igen_2_io_fire ? _GEN_4485 : _GEN_3461; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5510 = igen_2_io_fire ? _GEN_4486 : _GEN_3462; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5511 = igen_2_io_fire ? _GEN_4487 : _GEN_3463; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5512 = igen_2_io_fire ? _GEN_4488 : _GEN_3464; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5513 = igen_2_io_fire ? _GEN_4489 : _GEN_3465; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5514 = igen_2_io_fire ? _GEN_4490 : _GEN_3466; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5515 = igen_2_io_fire ? _GEN_4491 : _GEN_3467; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5516 = igen_2_io_fire ? _GEN_4492 : _GEN_3468; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5517 = igen_2_io_fire ? _GEN_4493 : _GEN_3469; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5518 = igen_2_io_fire ? _GEN_4494 : _GEN_3470; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5519 = igen_2_io_fire ? _GEN_4495 : _GEN_3471; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5520 = igen_2_io_fire ? _GEN_4496 : _GEN_3472; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5521 = igen_2_io_fire ? _GEN_4497 : _GEN_3473; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5522 = igen_2_io_fire ? _GEN_4498 : _GEN_3474; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5523 = igen_2_io_fire ? _GEN_4499 : _GEN_3475; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5524 = igen_2_io_fire ? _GEN_4500 : _GEN_3476; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5525 = igen_2_io_fire ? _GEN_4501 : _GEN_3477; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5526 = igen_2_io_fire ? _GEN_4502 : _GEN_3478; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5527 = igen_2_io_fire ? _GEN_4503 : _GEN_3479; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5528 = igen_2_io_fire ? _GEN_4504 : _GEN_3480; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5529 = igen_2_io_fire ? _GEN_4505 : _GEN_3481; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5530 = igen_2_io_fire ? _GEN_4506 : _GEN_3482; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5531 = igen_2_io_fire ? _GEN_4507 : _GEN_3483; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5532 = igen_2_io_fire ? _GEN_4508 : _GEN_3484; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5533 = igen_2_io_fire ? _GEN_4509 : _GEN_3485; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5534 = igen_2_io_fire ? _GEN_4510 : _GEN_3486; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5535 = igen_2_io_fire ? _GEN_4511 : _GEN_3487; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5536 = igen_2_io_fire ? _GEN_4512 : _GEN_3488; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5537 = igen_2_io_fire ? _GEN_4513 : _GEN_3489; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5538 = igen_2_io_fire ? _GEN_4514 : _GEN_3490; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5539 = igen_2_io_fire ? _GEN_4515 : _GEN_3491; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5540 = igen_2_io_fire ? _GEN_4516 : _GEN_3492; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5541 = igen_2_io_fire ? _GEN_4517 : _GEN_3493; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5542 = igen_2_io_fire ? _GEN_4518 : _GEN_3494; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5543 = igen_2_io_fire ? _GEN_4519 : _GEN_3495; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5544 = igen_2_io_fire ? _GEN_4520 : _GEN_3496; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5545 = igen_2_io_fire ? _GEN_4521 : _GEN_3497; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5546 = igen_2_io_fire ? _GEN_4522 : _GEN_3498; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5547 = igen_2_io_fire ? _GEN_4523 : _GEN_3499; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5548 = igen_2_io_fire ? _GEN_4524 : _GEN_3500; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5549 = igen_2_io_fire ? _GEN_4525 : _GEN_3501; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5550 = igen_2_io_fire ? _GEN_4526 : _GEN_3502; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5551 = igen_2_io_fire ? _GEN_4527 : _GEN_3503; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5552 = igen_2_io_fire ? _GEN_4528 : _GEN_3504; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5553 = igen_2_io_fire ? _GEN_4529 : _GEN_3505; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5554 = igen_2_io_fire ? _GEN_4530 : _GEN_3506; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5555 = igen_2_io_fire ? _GEN_4531 : _GEN_3507; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5556 = igen_2_io_fire ? _GEN_4532 : _GEN_3508; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5557 = igen_2_io_fire ? _GEN_4533 : _GEN_3509; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5558 = igen_2_io_fire ? _GEN_4534 : _GEN_3510; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5559 = igen_2_io_fire ? _GEN_4535 : _GEN_3511; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5560 = igen_2_io_fire ? _GEN_4536 : _GEN_3512; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5561 = igen_2_io_fire ? _GEN_4537 : _GEN_3513; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5562 = igen_2_io_fire ? _GEN_4538 : _GEN_3514; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5563 = igen_2_io_fire ? _GEN_4539 : _GEN_3515; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5564 = igen_2_io_fire ? _GEN_4540 : _GEN_3516; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5565 = igen_2_io_fire ? _GEN_4541 : _GEN_3517; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5566 = igen_2_io_fire ? _GEN_4542 : _GEN_3518; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5567 = igen_2_io_fire ? _GEN_4543 : _GEN_3519; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5568 = igen_2_io_fire ? _GEN_4544 : _GEN_3520; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5569 = igen_2_io_fire ? _GEN_4545 : _GEN_3521; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5570 = igen_2_io_fire ? _GEN_4546 : _GEN_3522; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5571 = igen_2_io_fire ? _GEN_4547 : _GEN_3523; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5572 = igen_2_io_fire ? _GEN_4548 : _GEN_3524; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5573 = igen_2_io_fire ? _GEN_4549 : _GEN_3525; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5574 = igen_2_io_fire ? _GEN_4550 : _GEN_3526; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5575 = igen_2_io_fire ? _GEN_4551 : _GEN_3527; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5576 = igen_2_io_fire ? _GEN_4552 : _GEN_3528; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5577 = igen_2_io_fire ? _GEN_4553 : _GEN_3529; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5578 = igen_2_io_fire ? _GEN_4554 : _GEN_3530; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5579 = igen_2_io_fire ? _GEN_4555 : _GEN_3531; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5580 = igen_2_io_fire ? _GEN_4556 : _GEN_3532; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5581 = igen_2_io_fire ? _GEN_4557 : _GEN_3533; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5582 = igen_2_io_fire ? _GEN_4558 : _GEN_3534; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5583 = igen_2_io_fire ? _GEN_4559 : _GEN_3535; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5584 = igen_2_io_fire ? _GEN_4560 : _GEN_3536; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5585 = igen_2_io_fire ? _GEN_4561 : _GEN_3537; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5586 = igen_2_io_fire ? _GEN_4562 : _GEN_3538; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5587 = igen_2_io_fire ? _GEN_4563 : _GEN_3539; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5588 = igen_2_io_fire ? _GEN_4564 : _GEN_3540; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5589 = igen_2_io_fire ? _GEN_4565 : _GEN_3541; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5590 = igen_2_io_fire ? _GEN_4566 : _GEN_3542; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5591 = igen_2_io_fire ? _GEN_4567 : _GEN_3543; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5592 = igen_2_io_fire ? _GEN_4568 : _GEN_3544; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5593 = igen_2_io_fire ? _GEN_4569 : _GEN_3545; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5594 = igen_2_io_fire ? _GEN_4570 : _GEN_3546; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5595 = igen_2_io_fire ? _GEN_4571 : _GEN_3547; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5596 = igen_2_io_fire ? _GEN_4572 : _GEN_3548; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5597 = igen_2_io_fire ? _GEN_4573 : _GEN_3549; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5598 = igen_2_io_fire ? _GEN_4574 : _GEN_3550; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5599 = igen_2_io_fire ? _GEN_4575 : _GEN_3551; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5600 = igen_2_io_fire ? _GEN_4576 : _GEN_3552; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5601 = igen_2_io_fire ? _GEN_4577 : _GEN_3553; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5602 = igen_2_io_fire ? _GEN_4578 : _GEN_3554; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5603 = igen_2_io_fire ? _GEN_4579 : _GEN_3555; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5604 = igen_2_io_fire ? _GEN_4580 : _GEN_3556; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5605 = igen_2_io_fire ? _GEN_4581 : _GEN_3557; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5606 = igen_2_io_fire ? _GEN_4582 : _GEN_3558; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5607 = igen_2_io_fire ? _GEN_4583 : _GEN_3559; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5608 = igen_2_io_fire ? _GEN_4584 : _GEN_3560; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5609 = igen_2_io_fire ? _GEN_4585 : _GEN_3561; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5610 = igen_2_io_fire ? _GEN_4586 : _GEN_3562; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5611 = igen_2_io_fire ? _GEN_4587 : _GEN_3563; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5612 = igen_2_io_fire ? _GEN_4588 : _GEN_3564; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5613 = igen_2_io_fire ? _GEN_4589 : _GEN_3565; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5614 = igen_2_io_fire ? _GEN_4590 : _GEN_3566; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5615 = igen_2_io_fire ? _GEN_4591 : _GEN_3567; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5616 = igen_2_io_fire ? _GEN_4592 : _GEN_3568; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5617 = igen_2_io_fire ? _GEN_4593 : _GEN_3569; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5618 = igen_2_io_fire ? _GEN_4594 : _GEN_3570; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5619 = igen_2_io_fire ? _GEN_4595 : _GEN_3571; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5620 = igen_2_io_fire ? _GEN_4596 : _GEN_3572; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5621 = igen_2_io_fire ? _GEN_4597 : _GEN_3573; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5622 = igen_2_io_fire ? _GEN_4598 : _GEN_3574; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5623 = igen_2_io_fire ? _GEN_4599 : _GEN_3575; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5624 = igen_2_io_fire ? _GEN_4600 : _GEN_3576; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5625 = igen_2_io_fire ? _GEN_4601 : _GEN_3577; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5626 = igen_2_io_fire ? _GEN_4602 : _GEN_3578; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5627 = igen_2_io_fire ? _GEN_4603 : _GEN_3579; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5628 = igen_2_io_fire ? _GEN_4604 : _GEN_3580; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5629 = igen_2_io_fire ? _GEN_4605 : _GEN_3581; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5630 = igen_2_io_fire ? _GEN_4606 : _GEN_3582; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5631 = igen_2_io_fire ? _GEN_4607 : _GEN_3583; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5632 = igen_2_io_fire ? _GEN_4608 : _GEN_3584; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5633 = igen_2_io_fire ? _GEN_4609 : _GEN_3585; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5634 = igen_2_io_fire ? _GEN_4610 : _GEN_3586; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5635 = igen_2_io_fire ? _GEN_4611 : _GEN_3587; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5636 = igen_2_io_fire ? _GEN_4612 : _GEN_3588; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5637 = igen_2_io_fire ? _GEN_4613 : _GEN_3589; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5638 = igen_2_io_fire ? _GEN_4614 : _GEN_3590; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5639 = igen_2_io_fire ? _GEN_4615 : _GEN_3591; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5640 = igen_2_io_fire ? _GEN_4616 : _GEN_3592; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5641 = igen_2_io_fire ? _GEN_4617 : _GEN_3593; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5642 = igen_2_io_fire ? _GEN_4618 : _GEN_3594; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5643 = igen_2_io_fire ? _GEN_4619 : _GEN_3595; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5644 = igen_2_io_fire ? _GEN_4620 : _GEN_3596; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5645 = igen_2_io_fire ? _GEN_4621 : _GEN_3597; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5646 = igen_2_io_fire ? _GEN_4622 : _GEN_3598; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5647 = igen_2_io_fire ? _GEN_4623 : _GEN_3599; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5648 = igen_2_io_fire ? _GEN_4624 : _GEN_3600; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5649 = igen_2_io_fire ? _GEN_4625 : _GEN_3601; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5650 = igen_2_io_fire ? _GEN_4626 : _GEN_3602; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5651 = igen_2_io_fire ? _GEN_4627 : _GEN_3603; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5652 = igen_2_io_fire ? _GEN_4628 : _GEN_3604; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5653 = igen_2_io_fire ? _GEN_4629 : _GEN_3605; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5654 = igen_2_io_fire ? _GEN_4630 : _GEN_3606; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5655 = igen_2_io_fire ? _GEN_4631 : _GEN_3607; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5656 = igen_2_io_fire ? _GEN_4632 : _GEN_3608; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5657 = igen_2_io_fire ? _GEN_4633 : _GEN_3609; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5658 = igen_2_io_fire ? _GEN_4634 : _GEN_3610; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5659 = igen_2_io_fire ? _GEN_4635 : _GEN_3611; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5660 = igen_2_io_fire ? _GEN_4636 : _GEN_3612; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5661 = igen_2_io_fire ? _GEN_4637 : _GEN_3613; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5662 = igen_2_io_fire ? _GEN_4638 : _GEN_3614; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5663 = igen_2_io_fire ? _GEN_4639 : _GEN_3615; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5664 = igen_2_io_fire ? _GEN_4640 : _GEN_3616; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5665 = igen_2_io_fire ? _GEN_4641 : _GEN_3617; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5666 = igen_2_io_fire ? _GEN_4642 : _GEN_3618; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5667 = igen_2_io_fire ? _GEN_4643 : _GEN_3619; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5668 = igen_2_io_fire ? _GEN_4644 : _GEN_3620; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5669 = igen_2_io_fire ? _GEN_4645 : _GEN_3621; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5670 = igen_2_io_fire ? _GEN_4646 : _GEN_3622; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5671 = igen_2_io_fire ? _GEN_4647 : _GEN_3623; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5672 = igen_2_io_fire ? _GEN_4648 : _GEN_3624; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5673 = igen_2_io_fire ? _GEN_4649 : _GEN_3625; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5674 = igen_2_io_fire ? _GEN_4650 : _GEN_3626; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5675 = igen_2_io_fire ? _GEN_4651 : _GEN_3627; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5676 = igen_2_io_fire ? _GEN_4652 : _GEN_3628; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5677 = igen_2_io_fire ? _GEN_4653 : _GEN_3629; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5678 = igen_2_io_fire ? _GEN_4654 : _GEN_3630; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5679 = igen_2_io_fire ? _GEN_4655 : _GEN_3631; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5680 = igen_2_io_fire ? _GEN_4656 : _GEN_3632; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5681 = igen_2_io_fire ? _GEN_4657 : _GEN_3633; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5682 = igen_2_io_fire ? _GEN_4658 : _GEN_3634; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5683 = igen_2_io_fire ? _GEN_4659 : _GEN_3635; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5684 = igen_2_io_fire ? _GEN_4660 : _GEN_3636; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5685 = igen_2_io_fire ? _GEN_4661 : _GEN_3637; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5686 = igen_2_io_fire ? _GEN_4662 : _GEN_3638; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5687 = igen_2_io_fire ? _GEN_4663 : _GEN_3639; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5688 = igen_2_io_fire ? _GEN_4664 : _GEN_3640; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5689 = igen_2_io_fire ? _GEN_4665 : _GEN_3641; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5690 = igen_2_io_fire ? _GEN_4666 : _GEN_3642; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5691 = igen_2_io_fire ? _GEN_4667 : _GEN_3643; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5692 = igen_2_io_fire ? _GEN_4668 : _GEN_3644; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5693 = igen_2_io_fire ? _GEN_4669 : _GEN_3645; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5694 = igen_2_io_fire ? _GEN_4670 : _GEN_3646; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5695 = igen_2_io_fire ? _GEN_4671 : _GEN_3647; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5696 = igen_2_io_fire ? _GEN_4672 : _GEN_3648; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5697 = igen_2_io_fire ? _GEN_4673 : _GEN_3649; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5698 = igen_2_io_fire ? _GEN_4674 : _GEN_3650; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5699 = igen_2_io_fire ? _GEN_4675 : _GEN_3651; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5700 = igen_2_io_fire ? _GEN_4676 : _GEN_3652; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5701 = igen_2_io_fire ? _GEN_4677 : _GEN_3653; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5702 = igen_2_io_fire ? _GEN_4678 : _GEN_3654; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5703 = igen_2_io_fire ? _GEN_4679 : _GEN_3655; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5704 = igen_2_io_fire ? _GEN_4680 : _GEN_3656; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5705 = igen_2_io_fire ? _GEN_4681 : _GEN_3657; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5706 = igen_2_io_fire ? _GEN_4682 : _GEN_3658; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5707 = igen_2_io_fire ? _GEN_4683 : _GEN_3659; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5708 = igen_2_io_fire ? _GEN_4684 : _GEN_3660; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5709 = igen_2_io_fire ? _GEN_4685 : _GEN_3661; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5710 = igen_2_io_fire ? _GEN_4686 : _GEN_3662; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5711 = igen_2_io_fire ? _GEN_4687 : _GEN_3663; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5712 = igen_2_io_fire ? _GEN_4688 : _GEN_3664; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5713 = igen_2_io_fire ? _GEN_4689 : _GEN_3665; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5714 = igen_2_io_fire ? _GEN_4690 : _GEN_3666; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5715 = igen_2_io_fire ? _GEN_4691 : _GEN_3667; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5716 = igen_2_io_fire ? _GEN_4692 : _GEN_3668; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5717 = igen_2_io_fire ? _GEN_4693 : _GEN_3669; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5718 = igen_2_io_fire ? _GEN_4694 : _GEN_3670; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5719 = igen_2_io_fire ? _GEN_4695 : _GEN_3671; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5720 = igen_2_io_fire ? _GEN_4696 : _GEN_3672; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5721 = igen_2_io_fire ? _GEN_4697 : _GEN_3673; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5722 = igen_2_io_fire ? _GEN_4698 : _GEN_3674; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5723 = igen_2_io_fire ? _GEN_4699 : _GEN_3675; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5724 = igen_2_io_fire ? _GEN_4700 : _GEN_3676; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5725 = igen_2_io_fire ? _GEN_4701 : _GEN_3677; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5726 = igen_2_io_fire ? _GEN_4702 : _GEN_3678; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5727 = igen_2_io_fire ? _GEN_4703 : _GEN_3679; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5728 = igen_2_io_fire ? _GEN_4704 : _GEN_3680; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5729 = igen_2_io_fire ? _GEN_4705 : _GEN_3681; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5730 = igen_2_io_fire ? _GEN_4706 : _GEN_3682; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5731 = igen_2_io_fire ? _GEN_4707 : _GEN_3683; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5732 = igen_2_io_fire ? _GEN_4708 : _GEN_3684; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5733 = igen_2_io_fire ? _GEN_4709 : _GEN_3685; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5734 = igen_2_io_fire ? _GEN_4710 : _GEN_3686; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5735 = igen_2_io_fire ? _GEN_4711 : _GEN_3687; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5736 = igen_2_io_fire ? _GEN_4712 : _GEN_3688; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5737 = igen_2_io_fire ? _GEN_4713 : _GEN_3689; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5738 = igen_2_io_fire ? _GEN_4714 : _GEN_3690; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5739 = igen_2_io_fire ? _GEN_4715 : _GEN_3691; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5740 = igen_2_io_fire ? _GEN_4716 : _GEN_3692; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5741 = igen_2_io_fire ? _GEN_4717 : _GEN_3693; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5742 = igen_2_io_fire ? _GEN_4718 : _GEN_3694; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5743 = igen_2_io_fire ? _GEN_4719 : _GEN_3695; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5744 = igen_2_io_fire ? _GEN_4720 : _GEN_3696; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5745 = igen_2_io_fire ? _GEN_4721 : _GEN_3697; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5746 = igen_2_io_fire ? _GEN_4722 : _GEN_3698; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5747 = igen_2_io_fire ? _GEN_4723 : _GEN_3699; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5748 = igen_2_io_fire ? _GEN_4724 : _GEN_3700; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5749 = igen_2_io_fire ? _GEN_4725 : _GEN_3701; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5750 = igen_2_io_fire ? _GEN_4726 : _GEN_3702; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5751 = igen_2_io_fire ? _GEN_4727 : _GEN_3703; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5752 = igen_2_io_fire ? _GEN_4728 : _GEN_3704; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5753 = igen_2_io_fire ? _GEN_4729 : _GEN_3705; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5754 = igen_2_io_fire ? _GEN_4730 : _GEN_3706; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5755 = igen_2_io_fire ? _GEN_4731 : _GEN_3707; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5756 = igen_2_io_fire ? _GEN_4732 : _GEN_3708; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5757 = igen_2_io_fire ? _GEN_4733 : _GEN_3709; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5758 = igen_2_io_fire ? _GEN_4734 : _GEN_3710; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5759 = igen_2_io_fire ? _GEN_4735 : _GEN_3711; // @[TestHarness.scala 178:25]
  wire [1:0] _GEN_5760 = igen_2_io_fire ? _GEN_4736 : _GEN_3712; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5761 = igen_2_io_fire ? _GEN_4737 : _GEN_3713; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5762 = igen_2_io_fire ? _GEN_4738 : _GEN_3714; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5763 = igen_2_io_fire ? _GEN_4739 : _GEN_3715; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5764 = igen_2_io_fire ? _GEN_4740 : _GEN_3716; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5765 = igen_2_io_fire ? _GEN_4741 : _GEN_3717; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5766 = igen_2_io_fire ? _GEN_4742 : _GEN_3718; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5767 = igen_2_io_fire ? _GEN_4743 : _GEN_3719; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5768 = igen_2_io_fire ? _GEN_4744 : _GEN_3720; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5769 = igen_2_io_fire ? _GEN_4745 : _GEN_3721; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5770 = igen_2_io_fire ? _GEN_4746 : _GEN_3722; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5771 = igen_2_io_fire ? _GEN_4747 : _GEN_3723; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5772 = igen_2_io_fire ? _GEN_4748 : _GEN_3724; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5773 = igen_2_io_fire ? _GEN_4749 : _GEN_3725; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5774 = igen_2_io_fire ? _GEN_4750 : _GEN_3726; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5775 = igen_2_io_fire ? _GEN_4751 : _GEN_3727; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5776 = igen_2_io_fire ? _GEN_4752 : _GEN_3728; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5777 = igen_2_io_fire ? _GEN_4753 : _GEN_3729; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5778 = igen_2_io_fire ? _GEN_4754 : _GEN_3730; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5779 = igen_2_io_fire ? _GEN_4755 : _GEN_3731; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5780 = igen_2_io_fire ? _GEN_4756 : _GEN_3732; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5781 = igen_2_io_fire ? _GEN_4757 : _GEN_3733; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5782 = igen_2_io_fire ? _GEN_4758 : _GEN_3734; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5783 = igen_2_io_fire ? _GEN_4759 : _GEN_3735; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5784 = igen_2_io_fire ? _GEN_4760 : _GEN_3736; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5785 = igen_2_io_fire ? _GEN_4761 : _GEN_3737; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5786 = igen_2_io_fire ? _GEN_4762 : _GEN_3738; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5787 = igen_2_io_fire ? _GEN_4763 : _GEN_3739; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5788 = igen_2_io_fire ? _GEN_4764 : _GEN_3740; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5789 = igen_2_io_fire ? _GEN_4765 : _GEN_3741; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5790 = igen_2_io_fire ? _GEN_4766 : _GEN_3742; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5791 = igen_2_io_fire ? _GEN_4767 : _GEN_3743; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5792 = igen_2_io_fire ? _GEN_4768 : _GEN_3744; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5793 = igen_2_io_fire ? _GEN_4769 : _GEN_3745; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5794 = igen_2_io_fire ? _GEN_4770 : _GEN_3746; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5795 = igen_2_io_fire ? _GEN_4771 : _GEN_3747; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5796 = igen_2_io_fire ? _GEN_4772 : _GEN_3748; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5797 = igen_2_io_fire ? _GEN_4773 : _GEN_3749; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5798 = igen_2_io_fire ? _GEN_4774 : _GEN_3750; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5799 = igen_2_io_fire ? _GEN_4775 : _GEN_3751; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5800 = igen_2_io_fire ? _GEN_4776 : _GEN_3752; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5801 = igen_2_io_fire ? _GEN_4777 : _GEN_3753; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5802 = igen_2_io_fire ? _GEN_4778 : _GEN_3754; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5803 = igen_2_io_fire ? _GEN_4779 : _GEN_3755; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5804 = igen_2_io_fire ? _GEN_4780 : _GEN_3756; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5805 = igen_2_io_fire ? _GEN_4781 : _GEN_3757; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5806 = igen_2_io_fire ? _GEN_4782 : _GEN_3758; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5807 = igen_2_io_fire ? _GEN_4783 : _GEN_3759; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5808 = igen_2_io_fire ? _GEN_4784 : _GEN_3760; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5809 = igen_2_io_fire ? _GEN_4785 : _GEN_3761; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5810 = igen_2_io_fire ? _GEN_4786 : _GEN_3762; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5811 = igen_2_io_fire ? _GEN_4787 : _GEN_3763; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5812 = igen_2_io_fire ? _GEN_4788 : _GEN_3764; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5813 = igen_2_io_fire ? _GEN_4789 : _GEN_3765; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5814 = igen_2_io_fire ? _GEN_4790 : _GEN_3766; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5815 = igen_2_io_fire ? _GEN_4791 : _GEN_3767; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5816 = igen_2_io_fire ? _GEN_4792 : _GEN_3768; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5817 = igen_2_io_fire ? _GEN_4793 : _GEN_3769; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5818 = igen_2_io_fire ? _GEN_4794 : _GEN_3770; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5819 = igen_2_io_fire ? _GEN_4795 : _GEN_3771; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5820 = igen_2_io_fire ? _GEN_4796 : _GEN_3772; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5821 = igen_2_io_fire ? _GEN_4797 : _GEN_3773; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5822 = igen_2_io_fire ? _GEN_4798 : _GEN_3774; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5823 = igen_2_io_fire ? _GEN_4799 : _GEN_3775; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5824 = igen_2_io_fire ? _GEN_4800 : _GEN_3776; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5825 = igen_2_io_fire ? _GEN_4801 : _GEN_3777; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5826 = igen_2_io_fire ? _GEN_4802 : _GEN_3778; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5827 = igen_2_io_fire ? _GEN_4803 : _GEN_3779; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5828 = igen_2_io_fire ? _GEN_4804 : _GEN_3780; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5829 = igen_2_io_fire ? _GEN_4805 : _GEN_3781; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5830 = igen_2_io_fire ? _GEN_4806 : _GEN_3782; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5831 = igen_2_io_fire ? _GEN_4807 : _GEN_3783; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5832 = igen_2_io_fire ? _GEN_4808 : _GEN_3784; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5833 = igen_2_io_fire ? _GEN_4809 : _GEN_3785; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5834 = igen_2_io_fire ? _GEN_4810 : _GEN_3786; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5835 = igen_2_io_fire ? _GEN_4811 : _GEN_3787; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5836 = igen_2_io_fire ? _GEN_4812 : _GEN_3788; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5837 = igen_2_io_fire ? _GEN_4813 : _GEN_3789; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5838 = igen_2_io_fire ? _GEN_4814 : _GEN_3790; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5839 = igen_2_io_fire ? _GEN_4815 : _GEN_3791; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5840 = igen_2_io_fire ? _GEN_4816 : _GEN_3792; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5841 = igen_2_io_fire ? _GEN_4817 : _GEN_3793; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5842 = igen_2_io_fire ? _GEN_4818 : _GEN_3794; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5843 = igen_2_io_fire ? _GEN_4819 : _GEN_3795; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5844 = igen_2_io_fire ? _GEN_4820 : _GEN_3796; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5845 = igen_2_io_fire ? _GEN_4821 : _GEN_3797; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5846 = igen_2_io_fire ? _GEN_4822 : _GEN_3798; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5847 = igen_2_io_fire ? _GEN_4823 : _GEN_3799; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5848 = igen_2_io_fire ? _GEN_4824 : _GEN_3800; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5849 = igen_2_io_fire ? _GEN_4825 : _GEN_3801; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5850 = igen_2_io_fire ? _GEN_4826 : _GEN_3802; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5851 = igen_2_io_fire ? _GEN_4827 : _GEN_3803; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5852 = igen_2_io_fire ? _GEN_4828 : _GEN_3804; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5853 = igen_2_io_fire ? _GEN_4829 : _GEN_3805; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5854 = igen_2_io_fire ? _GEN_4830 : _GEN_3806; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5855 = igen_2_io_fire ? _GEN_4831 : _GEN_3807; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5856 = igen_2_io_fire ? _GEN_4832 : _GEN_3808; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5857 = igen_2_io_fire ? _GEN_4833 : _GEN_3809; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5858 = igen_2_io_fire ? _GEN_4834 : _GEN_3810; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5859 = igen_2_io_fire ? _GEN_4835 : _GEN_3811; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5860 = igen_2_io_fire ? _GEN_4836 : _GEN_3812; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5861 = igen_2_io_fire ? _GEN_4837 : _GEN_3813; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5862 = igen_2_io_fire ? _GEN_4838 : _GEN_3814; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5863 = igen_2_io_fire ? _GEN_4839 : _GEN_3815; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5864 = igen_2_io_fire ? _GEN_4840 : _GEN_3816; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5865 = igen_2_io_fire ? _GEN_4841 : _GEN_3817; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5866 = igen_2_io_fire ? _GEN_4842 : _GEN_3818; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5867 = igen_2_io_fire ? _GEN_4843 : _GEN_3819; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5868 = igen_2_io_fire ? _GEN_4844 : _GEN_3820; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5869 = igen_2_io_fire ? _GEN_4845 : _GEN_3821; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5870 = igen_2_io_fire ? _GEN_4846 : _GEN_3822; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5871 = igen_2_io_fire ? _GEN_4847 : _GEN_3823; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5872 = igen_2_io_fire ? _GEN_4848 : _GEN_3824; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5873 = igen_2_io_fire ? _GEN_4849 : _GEN_3825; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5874 = igen_2_io_fire ? _GEN_4850 : _GEN_3826; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5875 = igen_2_io_fire ? _GEN_4851 : _GEN_3827; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5876 = igen_2_io_fire ? _GEN_4852 : _GEN_3828; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5877 = igen_2_io_fire ? _GEN_4853 : _GEN_3829; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5878 = igen_2_io_fire ? _GEN_4854 : _GEN_3830; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5879 = igen_2_io_fire ? _GEN_4855 : _GEN_3831; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5880 = igen_2_io_fire ? _GEN_4856 : _GEN_3832; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5881 = igen_2_io_fire ? _GEN_4857 : _GEN_3833; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5882 = igen_2_io_fire ? _GEN_4858 : _GEN_3834; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5883 = igen_2_io_fire ? _GEN_4859 : _GEN_3835; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5884 = igen_2_io_fire ? _GEN_4860 : _GEN_3836; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5885 = igen_2_io_fire ? _GEN_4861 : _GEN_3837; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5886 = igen_2_io_fire ? _GEN_4862 : _GEN_3838; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5887 = igen_2_io_fire ? _GEN_4863 : _GEN_3839; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5888 = igen_2_io_fire ? _GEN_4864 : _GEN_3840; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5889 = igen_2_io_fire ? _GEN_4865 : _GEN_3841; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5890 = igen_2_io_fire ? _GEN_4866 : _GEN_3842; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5891 = igen_2_io_fire ? _GEN_4867 : _GEN_3843; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5892 = igen_2_io_fire ? _GEN_4868 : _GEN_3844; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5893 = igen_2_io_fire ? _GEN_4869 : _GEN_3845; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5894 = igen_2_io_fire ? _GEN_4870 : _GEN_3846; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5895 = igen_2_io_fire ? _GEN_4871 : _GEN_3847; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5896 = igen_2_io_fire ? _GEN_4872 : _GEN_3848; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5897 = igen_2_io_fire ? _GEN_4873 : _GEN_3849; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5898 = igen_2_io_fire ? _GEN_4874 : _GEN_3850; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5899 = igen_2_io_fire ? _GEN_4875 : _GEN_3851; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5900 = igen_2_io_fire ? _GEN_4876 : _GEN_3852; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5901 = igen_2_io_fire ? _GEN_4877 : _GEN_3853; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5902 = igen_2_io_fire ? _GEN_4878 : _GEN_3854; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5903 = igen_2_io_fire ? _GEN_4879 : _GEN_3855; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5904 = igen_2_io_fire ? _GEN_4880 : _GEN_3856; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5905 = igen_2_io_fire ? _GEN_4881 : _GEN_3857; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5906 = igen_2_io_fire ? _GEN_4882 : _GEN_3858; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5907 = igen_2_io_fire ? _GEN_4883 : _GEN_3859; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5908 = igen_2_io_fire ? _GEN_4884 : _GEN_3860; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5909 = igen_2_io_fire ? _GEN_4885 : _GEN_3861; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5910 = igen_2_io_fire ? _GEN_4886 : _GEN_3862; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5911 = igen_2_io_fire ? _GEN_4887 : _GEN_3863; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5912 = igen_2_io_fire ? _GEN_4888 : _GEN_3864; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5913 = igen_2_io_fire ? _GEN_4889 : _GEN_3865; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5914 = igen_2_io_fire ? _GEN_4890 : _GEN_3866; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5915 = igen_2_io_fire ? _GEN_4891 : _GEN_3867; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5916 = igen_2_io_fire ? _GEN_4892 : _GEN_3868; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5917 = igen_2_io_fire ? _GEN_4893 : _GEN_3869; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5918 = igen_2_io_fire ? _GEN_4894 : _GEN_3870; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5919 = igen_2_io_fire ? _GEN_4895 : _GEN_3871; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5920 = igen_2_io_fire ? _GEN_4896 : _GEN_3872; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5921 = igen_2_io_fire ? _GEN_4897 : _GEN_3873; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5922 = igen_2_io_fire ? _GEN_4898 : _GEN_3874; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5923 = igen_2_io_fire ? _GEN_4899 : _GEN_3875; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5924 = igen_2_io_fire ? _GEN_4900 : _GEN_3876; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5925 = igen_2_io_fire ? _GEN_4901 : _GEN_3877; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5926 = igen_2_io_fire ? _GEN_4902 : _GEN_3878; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5927 = igen_2_io_fire ? _GEN_4903 : _GEN_3879; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5928 = igen_2_io_fire ? _GEN_4904 : _GEN_3880; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5929 = igen_2_io_fire ? _GEN_4905 : _GEN_3881; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5930 = igen_2_io_fire ? _GEN_4906 : _GEN_3882; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5931 = igen_2_io_fire ? _GEN_4907 : _GEN_3883; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5932 = igen_2_io_fire ? _GEN_4908 : _GEN_3884; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5933 = igen_2_io_fire ? _GEN_4909 : _GEN_3885; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5934 = igen_2_io_fire ? _GEN_4910 : _GEN_3886; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5935 = igen_2_io_fire ? _GEN_4911 : _GEN_3887; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5936 = igen_2_io_fire ? _GEN_4912 : _GEN_3888; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5937 = igen_2_io_fire ? _GEN_4913 : _GEN_3889; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5938 = igen_2_io_fire ? _GEN_4914 : _GEN_3890; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5939 = igen_2_io_fire ? _GEN_4915 : _GEN_3891; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5940 = igen_2_io_fire ? _GEN_4916 : _GEN_3892; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5941 = igen_2_io_fire ? _GEN_4917 : _GEN_3893; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5942 = igen_2_io_fire ? _GEN_4918 : _GEN_3894; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5943 = igen_2_io_fire ? _GEN_4919 : _GEN_3895; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5944 = igen_2_io_fire ? _GEN_4920 : _GEN_3896; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5945 = igen_2_io_fire ? _GEN_4921 : _GEN_3897; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5946 = igen_2_io_fire ? _GEN_4922 : _GEN_3898; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5947 = igen_2_io_fire ? _GEN_4923 : _GEN_3899; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5948 = igen_2_io_fire ? _GEN_4924 : _GEN_3900; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5949 = igen_2_io_fire ? _GEN_4925 : _GEN_3901; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5950 = igen_2_io_fire ? _GEN_4926 : _GEN_3902; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5951 = igen_2_io_fire ? _GEN_4927 : _GEN_3903; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5952 = igen_2_io_fire ? _GEN_4928 : _GEN_3904; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5953 = igen_2_io_fire ? _GEN_4929 : _GEN_3905; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5954 = igen_2_io_fire ? _GEN_4930 : _GEN_3906; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5955 = igen_2_io_fire ? _GEN_4931 : _GEN_3907; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5956 = igen_2_io_fire ? _GEN_4932 : _GEN_3908; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5957 = igen_2_io_fire ? _GEN_4933 : _GEN_3909; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5958 = igen_2_io_fire ? _GEN_4934 : _GEN_3910; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5959 = igen_2_io_fire ? _GEN_4935 : _GEN_3911; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5960 = igen_2_io_fire ? _GEN_4936 : _GEN_3912; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5961 = igen_2_io_fire ? _GEN_4937 : _GEN_3913; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5962 = igen_2_io_fire ? _GEN_4938 : _GEN_3914; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5963 = igen_2_io_fire ? _GEN_4939 : _GEN_3915; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5964 = igen_2_io_fire ? _GEN_4940 : _GEN_3916; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5965 = igen_2_io_fire ? _GEN_4941 : _GEN_3917; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5966 = igen_2_io_fire ? _GEN_4942 : _GEN_3918; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5967 = igen_2_io_fire ? _GEN_4943 : _GEN_3919; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5968 = igen_2_io_fire ? _GEN_4944 : _GEN_3920; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5969 = igen_2_io_fire ? _GEN_4945 : _GEN_3921; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5970 = igen_2_io_fire ? _GEN_4946 : _GEN_3922; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5971 = igen_2_io_fire ? _GEN_4947 : _GEN_3923; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5972 = igen_2_io_fire ? _GEN_4948 : _GEN_3924; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5973 = igen_2_io_fire ? _GEN_4949 : _GEN_3925; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5974 = igen_2_io_fire ? _GEN_4950 : _GEN_3926; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5975 = igen_2_io_fire ? _GEN_4951 : _GEN_3927; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5976 = igen_2_io_fire ? _GEN_4952 : _GEN_3928; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5977 = igen_2_io_fire ? _GEN_4953 : _GEN_3929; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5978 = igen_2_io_fire ? _GEN_4954 : _GEN_3930; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5979 = igen_2_io_fire ? _GEN_4955 : _GEN_3931; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5980 = igen_2_io_fire ? _GEN_4956 : _GEN_3932; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5981 = igen_2_io_fire ? _GEN_4957 : _GEN_3933; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5982 = igen_2_io_fire ? _GEN_4958 : _GEN_3934; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5983 = igen_2_io_fire ? _GEN_4959 : _GEN_3935; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5984 = igen_2_io_fire ? _GEN_4960 : _GEN_3936; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5985 = igen_2_io_fire ? _GEN_4961 : _GEN_3937; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5986 = igen_2_io_fire ? _GEN_4962 : _GEN_3938; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5987 = igen_2_io_fire ? _GEN_4963 : _GEN_3939; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5988 = igen_2_io_fire ? _GEN_4964 : _GEN_3940; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5989 = igen_2_io_fire ? _GEN_4965 : _GEN_3941; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5990 = igen_2_io_fire ? _GEN_4966 : _GEN_3942; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5991 = igen_2_io_fire ? _GEN_4967 : _GEN_3943; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5992 = igen_2_io_fire ? _GEN_4968 : _GEN_3944; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5993 = igen_2_io_fire ? _GEN_4969 : _GEN_3945; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5994 = igen_2_io_fire ? _GEN_4970 : _GEN_3946; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5995 = igen_2_io_fire ? _GEN_4971 : _GEN_3947; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5996 = igen_2_io_fire ? _GEN_4972 : _GEN_3948; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5997 = igen_2_io_fire ? _GEN_4973 : _GEN_3949; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5998 = igen_2_io_fire ? _GEN_4974 : _GEN_3950; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_5999 = igen_2_io_fire ? _GEN_4975 : _GEN_3951; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_6000 = igen_2_io_fire ? _GEN_4976 : _GEN_3952; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_6001 = igen_2_io_fire ? _GEN_4977 : _GEN_3953; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_6002 = igen_2_io_fire ? _GEN_4978 : _GEN_3954; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_6003 = igen_2_io_fire ? _GEN_4979 : _GEN_3955; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_6004 = igen_2_io_fire ? _GEN_4980 : _GEN_3956; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_6005 = igen_2_io_fire ? _GEN_4981 : _GEN_3957; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_6006 = igen_2_io_fire ? _GEN_4982 : _GEN_3958; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_6007 = igen_2_io_fire ? _GEN_4983 : _GEN_3959; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_6008 = igen_2_io_fire ? _GEN_4984 : _GEN_3960; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_6009 = igen_2_io_fire ? _GEN_4985 : _GEN_3961; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_6010 = igen_2_io_fire ? _GEN_4986 : _GEN_3962; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_6011 = igen_2_io_fire ? _GEN_4987 : _GEN_3963; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_6012 = igen_2_io_fire ? _GEN_4988 : _GEN_3964; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_6013 = igen_2_io_fire ? _GEN_4989 : _GEN_3965; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_6014 = igen_2_io_fire ? _GEN_4990 : _GEN_3966; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_6015 = igen_2_io_fire ? _GEN_4991 : _GEN_3967; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_6016 = igen_2_io_fire ? _GEN_4992 : _GEN_3968; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6017 = igen_2_io_fire ? _GEN_4993 : _GEN_3969; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6018 = igen_2_io_fire ? _GEN_4994 : _GEN_3970; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6019 = igen_2_io_fire ? _GEN_4995 : _GEN_3971; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6020 = igen_2_io_fire ? _GEN_4996 : _GEN_3972; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6021 = igen_2_io_fire ? _GEN_4997 : _GEN_3973; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6022 = igen_2_io_fire ? _GEN_4998 : _GEN_3974; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6023 = igen_2_io_fire ? _GEN_4999 : _GEN_3975; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6024 = igen_2_io_fire ? _GEN_5000 : _GEN_3976; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6025 = igen_2_io_fire ? _GEN_5001 : _GEN_3977; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6026 = igen_2_io_fire ? _GEN_5002 : _GEN_3978; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6027 = igen_2_io_fire ? _GEN_5003 : _GEN_3979; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6028 = igen_2_io_fire ? _GEN_5004 : _GEN_3980; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6029 = igen_2_io_fire ? _GEN_5005 : _GEN_3981; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6030 = igen_2_io_fire ? _GEN_5006 : _GEN_3982; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6031 = igen_2_io_fire ? _GEN_5007 : _GEN_3983; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6032 = igen_2_io_fire ? _GEN_5008 : _GEN_3984; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6033 = igen_2_io_fire ? _GEN_5009 : _GEN_3985; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6034 = igen_2_io_fire ? _GEN_5010 : _GEN_3986; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6035 = igen_2_io_fire ? _GEN_5011 : _GEN_3987; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6036 = igen_2_io_fire ? _GEN_5012 : _GEN_3988; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6037 = igen_2_io_fire ? _GEN_5013 : _GEN_3989; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6038 = igen_2_io_fire ? _GEN_5014 : _GEN_3990; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6039 = igen_2_io_fire ? _GEN_5015 : _GEN_3991; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6040 = igen_2_io_fire ? _GEN_5016 : _GEN_3992; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6041 = igen_2_io_fire ? _GEN_5017 : _GEN_3993; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6042 = igen_2_io_fire ? _GEN_5018 : _GEN_3994; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6043 = igen_2_io_fire ? _GEN_5019 : _GEN_3995; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6044 = igen_2_io_fire ? _GEN_5020 : _GEN_3996; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6045 = igen_2_io_fire ? _GEN_5021 : _GEN_3997; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6046 = igen_2_io_fire ? _GEN_5022 : _GEN_3998; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6047 = igen_2_io_fire ? _GEN_5023 : _GEN_3999; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6048 = igen_2_io_fire ? _GEN_5024 : _GEN_4000; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6049 = igen_2_io_fire ? _GEN_5025 : _GEN_4001; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6050 = igen_2_io_fire ? _GEN_5026 : _GEN_4002; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6051 = igen_2_io_fire ? _GEN_5027 : _GEN_4003; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6052 = igen_2_io_fire ? _GEN_5028 : _GEN_4004; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6053 = igen_2_io_fire ? _GEN_5029 : _GEN_4005; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6054 = igen_2_io_fire ? _GEN_5030 : _GEN_4006; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6055 = igen_2_io_fire ? _GEN_5031 : _GEN_4007; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6056 = igen_2_io_fire ? _GEN_5032 : _GEN_4008; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6057 = igen_2_io_fire ? _GEN_5033 : _GEN_4009; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6058 = igen_2_io_fire ? _GEN_5034 : _GEN_4010; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6059 = igen_2_io_fire ? _GEN_5035 : _GEN_4011; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6060 = igen_2_io_fire ? _GEN_5036 : _GEN_4012; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6061 = igen_2_io_fire ? _GEN_5037 : _GEN_4013; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6062 = igen_2_io_fire ? _GEN_5038 : _GEN_4014; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6063 = igen_2_io_fire ? _GEN_5039 : _GEN_4015; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6064 = igen_2_io_fire ? _GEN_5040 : _GEN_4016; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6065 = igen_2_io_fire ? _GEN_5041 : _GEN_4017; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6066 = igen_2_io_fire ? _GEN_5042 : _GEN_4018; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6067 = igen_2_io_fire ? _GEN_5043 : _GEN_4019; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6068 = igen_2_io_fire ? _GEN_5044 : _GEN_4020; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6069 = igen_2_io_fire ? _GEN_5045 : _GEN_4021; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6070 = igen_2_io_fire ? _GEN_5046 : _GEN_4022; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6071 = igen_2_io_fire ? _GEN_5047 : _GEN_4023; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6072 = igen_2_io_fire ? _GEN_5048 : _GEN_4024; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6073 = igen_2_io_fire ? _GEN_5049 : _GEN_4025; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6074 = igen_2_io_fire ? _GEN_5050 : _GEN_4026; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6075 = igen_2_io_fire ? _GEN_5051 : _GEN_4027; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6076 = igen_2_io_fire ? _GEN_5052 : _GEN_4028; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6077 = igen_2_io_fire ? _GEN_5053 : _GEN_4029; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6078 = igen_2_io_fire ? _GEN_5054 : _GEN_4030; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6079 = igen_2_io_fire ? _GEN_5055 : _GEN_4031; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6080 = igen_2_io_fire ? _GEN_5056 : _GEN_4032; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6081 = igen_2_io_fire ? _GEN_5057 : _GEN_4033; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6082 = igen_2_io_fire ? _GEN_5058 : _GEN_4034; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6083 = igen_2_io_fire ? _GEN_5059 : _GEN_4035; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6084 = igen_2_io_fire ? _GEN_5060 : _GEN_4036; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6085 = igen_2_io_fire ? _GEN_5061 : _GEN_4037; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6086 = igen_2_io_fire ? _GEN_5062 : _GEN_4038; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6087 = igen_2_io_fire ? _GEN_5063 : _GEN_4039; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6088 = igen_2_io_fire ? _GEN_5064 : _GEN_4040; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6089 = igen_2_io_fire ? _GEN_5065 : _GEN_4041; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6090 = igen_2_io_fire ? _GEN_5066 : _GEN_4042; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6091 = igen_2_io_fire ? _GEN_5067 : _GEN_4043; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6092 = igen_2_io_fire ? _GEN_5068 : _GEN_4044; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6093 = igen_2_io_fire ? _GEN_5069 : _GEN_4045; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6094 = igen_2_io_fire ? _GEN_5070 : _GEN_4046; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6095 = igen_2_io_fire ? _GEN_5071 : _GEN_4047; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6096 = igen_2_io_fire ? _GEN_5072 : _GEN_4048; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6097 = igen_2_io_fire ? _GEN_5073 : _GEN_4049; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6098 = igen_2_io_fire ? _GEN_5074 : _GEN_4050; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6099 = igen_2_io_fire ? _GEN_5075 : _GEN_4051; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6100 = igen_2_io_fire ? _GEN_5076 : _GEN_4052; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6101 = igen_2_io_fire ? _GEN_5077 : _GEN_4053; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6102 = igen_2_io_fire ? _GEN_5078 : _GEN_4054; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6103 = igen_2_io_fire ? _GEN_5079 : _GEN_4055; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6104 = igen_2_io_fire ? _GEN_5080 : _GEN_4056; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6105 = igen_2_io_fire ? _GEN_5081 : _GEN_4057; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6106 = igen_2_io_fire ? _GEN_5082 : _GEN_4058; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6107 = igen_2_io_fire ? _GEN_5083 : _GEN_4059; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6108 = igen_2_io_fire ? _GEN_5084 : _GEN_4060; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6109 = igen_2_io_fire ? _GEN_5085 : _GEN_4061; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6110 = igen_2_io_fire ? _GEN_5086 : _GEN_4062; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6111 = igen_2_io_fire ? _GEN_5087 : _GEN_4063; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6112 = igen_2_io_fire ? _GEN_5088 : _GEN_4064; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6113 = igen_2_io_fire ? _GEN_5089 : _GEN_4065; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6114 = igen_2_io_fire ? _GEN_5090 : _GEN_4066; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6115 = igen_2_io_fire ? _GEN_5091 : _GEN_4067; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6116 = igen_2_io_fire ? _GEN_5092 : _GEN_4068; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6117 = igen_2_io_fire ? _GEN_5093 : _GEN_4069; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6118 = igen_2_io_fire ? _GEN_5094 : _GEN_4070; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6119 = igen_2_io_fire ? _GEN_5095 : _GEN_4071; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6120 = igen_2_io_fire ? _GEN_5096 : _GEN_4072; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6121 = igen_2_io_fire ? _GEN_5097 : _GEN_4073; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6122 = igen_2_io_fire ? _GEN_5098 : _GEN_4074; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6123 = igen_2_io_fire ? _GEN_5099 : _GEN_4075; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6124 = igen_2_io_fire ? _GEN_5100 : _GEN_4076; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6125 = igen_2_io_fire ? _GEN_5101 : _GEN_4077; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6126 = igen_2_io_fire ? _GEN_5102 : _GEN_4078; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6127 = igen_2_io_fire ? _GEN_5103 : _GEN_4079; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6128 = igen_2_io_fire ? _GEN_5104 : _GEN_4080; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6129 = igen_2_io_fire ? _GEN_5105 : _GEN_4081; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6130 = igen_2_io_fire ? _GEN_5106 : _GEN_4082; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6131 = igen_2_io_fire ? _GEN_5107 : _GEN_4083; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6132 = igen_2_io_fire ? _GEN_5108 : _GEN_4084; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6133 = igen_2_io_fire ? _GEN_5109 : _GEN_4085; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6134 = igen_2_io_fire ? _GEN_5110 : _GEN_4086; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6135 = igen_2_io_fire ? _GEN_5111 : _GEN_4087; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6136 = igen_2_io_fire ? _GEN_5112 : _GEN_4088; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6137 = igen_2_io_fire ? _GEN_5113 : _GEN_4089; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6138 = igen_2_io_fire ? _GEN_5114 : _GEN_4090; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6139 = igen_2_io_fire ? _GEN_5115 : _GEN_4091; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6140 = igen_2_io_fire ? _GEN_5116 : _GEN_4092; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6141 = igen_2_io_fire ? _GEN_5117 : _GEN_4093; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6142 = igen_2_io_fire ? _GEN_5118 : _GEN_4094; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6143 = igen_2_io_fire ? _GEN_5119 : _GEN_4095; // @[TestHarness.scala 178:25]
  wire [63:0] _GEN_6144 = igen_2_io_fire ? _GEN_5120 : _GEN_4096; // @[TestHarness.scala 178:25]
  wire  _igen_io_rob_ready_T_17 = rob_alloc_avail_3 & rob_alloc_fires_3 & _igen_io_rob_ready_T_1; // @[TestHarness.scala 174:72]
  wire [63:0] _rob_payload_WIRE_7 = igen_3_io_out_bits_payload; // @[TestHarness.scala 179:{72,72}]
  wire [15:0] _GEN_6401 = 7'h0 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5377; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6402 = 7'h1 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5378; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6403 = 7'h2 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5379; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6404 = 7'h3 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5380; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6405 = 7'h4 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5381; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6406 = 7'h5 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5382; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6407 = 7'h6 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5383; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6408 = 7'h7 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5384; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6409 = 7'h8 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5385; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6410 = 7'h9 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5386; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6411 = 7'ha == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5387; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6412 = 7'hb == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5388; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6413 = 7'hc == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5389; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6414 = 7'hd == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5390; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6415 = 7'he == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5391; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6416 = 7'hf == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5392; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6417 = 7'h10 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5393; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6418 = 7'h11 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5394; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6419 = 7'h12 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5395; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6420 = 7'h13 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5396; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6421 = 7'h14 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5397; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6422 = 7'h15 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5398; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6423 = 7'h16 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5399; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6424 = 7'h17 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5400; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6425 = 7'h18 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5401; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6426 = 7'h19 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5402; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6427 = 7'h1a == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5403; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6428 = 7'h1b == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5404; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6429 = 7'h1c == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5405; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6430 = 7'h1d == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5406; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6431 = 7'h1e == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5407; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6432 = 7'h1f == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5408; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6433 = 7'h20 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5409; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6434 = 7'h21 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5410; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6435 = 7'h22 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5411; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6436 = 7'h23 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5412; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6437 = 7'h24 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5413; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6438 = 7'h25 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5414; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6439 = 7'h26 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5415; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6440 = 7'h27 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5416; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6441 = 7'h28 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5417; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6442 = 7'h29 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5418; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6443 = 7'h2a == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5419; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6444 = 7'h2b == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5420; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6445 = 7'h2c == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5421; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6446 = 7'h2d == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5422; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6447 = 7'h2e == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5423; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6448 = 7'h2f == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5424; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6449 = 7'h30 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5425; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6450 = 7'h31 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5426; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6451 = 7'h32 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5427; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6452 = 7'h33 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5428; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6453 = 7'h34 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5429; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6454 = 7'h35 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5430; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6455 = 7'h36 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5431; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6456 = 7'h37 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5432; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6457 = 7'h38 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5433; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6458 = 7'h39 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5434; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6459 = 7'h3a == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5435; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6460 = 7'h3b == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5436; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6461 = 7'h3c == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5437; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6462 = 7'h3d == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5438; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6463 = 7'h3e == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5439; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6464 = 7'h3f == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5440; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6465 = 7'h40 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5441; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6466 = 7'h41 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5442; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6467 = 7'h42 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5443; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6468 = 7'h43 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5444; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6469 = 7'h44 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5445; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6470 = 7'h45 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5446; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6471 = 7'h46 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5447; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6472 = 7'h47 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5448; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6473 = 7'h48 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5449; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6474 = 7'h49 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5450; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6475 = 7'h4a == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5451; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6476 = 7'h4b == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5452; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6477 = 7'h4c == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5453; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6478 = 7'h4d == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5454; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6479 = 7'h4e == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5455; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6480 = 7'h4f == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5456; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6481 = 7'h50 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5457; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6482 = 7'h51 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5458; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6483 = 7'h52 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5459; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6484 = 7'h53 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5460; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6485 = 7'h54 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5461; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6486 = 7'h55 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5462; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6487 = 7'h56 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5463; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6488 = 7'h57 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5464; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6489 = 7'h58 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5465; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6490 = 7'h59 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5466; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6491 = 7'h5a == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5467; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6492 = 7'h5b == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5468; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6493 = 7'h5c == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5469; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6494 = 7'h5d == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5470; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6495 = 7'h5e == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5471; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6496 = 7'h5f == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5472; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6497 = 7'h60 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5473; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6498 = 7'h61 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5474; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6499 = 7'h62 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5475; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6500 = 7'h63 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5476; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6501 = 7'h64 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5477; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6502 = 7'h65 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5478; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6503 = 7'h66 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5479; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6504 = 7'h67 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5480; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6505 = 7'h68 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5481; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6506 = 7'h69 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5482; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6507 = 7'h6a == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5483; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6508 = 7'h6b == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5484; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6509 = 7'h6c == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5485; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6510 = 7'h6d == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5486; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6511 = 7'h6e == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5487; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6512 = 7'h6f == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5488; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6513 = 7'h70 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5489; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6514 = 7'h71 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5490; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6515 = 7'h72 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5491; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6516 = 7'h73 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5492; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6517 = 7'h74 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5493; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6518 = 7'h75 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5494; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6519 = 7'h76 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5495; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6520 = 7'h77 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5496; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6521 = 7'h78 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5497; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6522 = 7'h79 == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5498; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6523 = 7'h7a == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5499; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6524 = 7'h7b == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5500; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6525 = 7'h7c == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5501; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6526 = 7'h7d == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5502; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6527 = 7'h7e == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5503; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_6528 = 7'h7f == rob_alloc_ids_3 ? _rob_payload_WIRE_7[15:0] : _GEN_5504; // @[TestHarness.scala 179:{36,36}]
  wire [1:0] _rob_egress_id_T_65 = igen_3_io_out_bits_egress_id; // @[TestHarness.scala 180:{36,36}]
  wire [3:0] _rob_n_flits_T_69 = igen_3_io_n_flits; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_6913 = 7'h0 == rob_alloc_ids_3 ? 4'h0 : _GEN_5889; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6914 = 7'h1 == rob_alloc_ids_3 ? 4'h0 : _GEN_5890; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6915 = 7'h2 == rob_alloc_ids_3 ? 4'h0 : _GEN_5891; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6916 = 7'h3 == rob_alloc_ids_3 ? 4'h0 : _GEN_5892; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6917 = 7'h4 == rob_alloc_ids_3 ? 4'h0 : _GEN_5893; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6918 = 7'h5 == rob_alloc_ids_3 ? 4'h0 : _GEN_5894; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6919 = 7'h6 == rob_alloc_ids_3 ? 4'h0 : _GEN_5895; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6920 = 7'h7 == rob_alloc_ids_3 ? 4'h0 : _GEN_5896; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6921 = 7'h8 == rob_alloc_ids_3 ? 4'h0 : _GEN_5897; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6922 = 7'h9 == rob_alloc_ids_3 ? 4'h0 : _GEN_5898; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6923 = 7'ha == rob_alloc_ids_3 ? 4'h0 : _GEN_5899; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6924 = 7'hb == rob_alloc_ids_3 ? 4'h0 : _GEN_5900; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6925 = 7'hc == rob_alloc_ids_3 ? 4'h0 : _GEN_5901; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6926 = 7'hd == rob_alloc_ids_3 ? 4'h0 : _GEN_5902; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6927 = 7'he == rob_alloc_ids_3 ? 4'h0 : _GEN_5903; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6928 = 7'hf == rob_alloc_ids_3 ? 4'h0 : _GEN_5904; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6929 = 7'h10 == rob_alloc_ids_3 ? 4'h0 : _GEN_5905; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6930 = 7'h11 == rob_alloc_ids_3 ? 4'h0 : _GEN_5906; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6931 = 7'h12 == rob_alloc_ids_3 ? 4'h0 : _GEN_5907; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6932 = 7'h13 == rob_alloc_ids_3 ? 4'h0 : _GEN_5908; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6933 = 7'h14 == rob_alloc_ids_3 ? 4'h0 : _GEN_5909; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6934 = 7'h15 == rob_alloc_ids_3 ? 4'h0 : _GEN_5910; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6935 = 7'h16 == rob_alloc_ids_3 ? 4'h0 : _GEN_5911; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6936 = 7'h17 == rob_alloc_ids_3 ? 4'h0 : _GEN_5912; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6937 = 7'h18 == rob_alloc_ids_3 ? 4'h0 : _GEN_5913; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6938 = 7'h19 == rob_alloc_ids_3 ? 4'h0 : _GEN_5914; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6939 = 7'h1a == rob_alloc_ids_3 ? 4'h0 : _GEN_5915; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6940 = 7'h1b == rob_alloc_ids_3 ? 4'h0 : _GEN_5916; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6941 = 7'h1c == rob_alloc_ids_3 ? 4'h0 : _GEN_5917; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6942 = 7'h1d == rob_alloc_ids_3 ? 4'h0 : _GEN_5918; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6943 = 7'h1e == rob_alloc_ids_3 ? 4'h0 : _GEN_5919; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6944 = 7'h1f == rob_alloc_ids_3 ? 4'h0 : _GEN_5920; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6945 = 7'h20 == rob_alloc_ids_3 ? 4'h0 : _GEN_5921; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6946 = 7'h21 == rob_alloc_ids_3 ? 4'h0 : _GEN_5922; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6947 = 7'h22 == rob_alloc_ids_3 ? 4'h0 : _GEN_5923; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6948 = 7'h23 == rob_alloc_ids_3 ? 4'h0 : _GEN_5924; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6949 = 7'h24 == rob_alloc_ids_3 ? 4'h0 : _GEN_5925; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6950 = 7'h25 == rob_alloc_ids_3 ? 4'h0 : _GEN_5926; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6951 = 7'h26 == rob_alloc_ids_3 ? 4'h0 : _GEN_5927; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6952 = 7'h27 == rob_alloc_ids_3 ? 4'h0 : _GEN_5928; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6953 = 7'h28 == rob_alloc_ids_3 ? 4'h0 : _GEN_5929; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6954 = 7'h29 == rob_alloc_ids_3 ? 4'h0 : _GEN_5930; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6955 = 7'h2a == rob_alloc_ids_3 ? 4'h0 : _GEN_5931; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6956 = 7'h2b == rob_alloc_ids_3 ? 4'h0 : _GEN_5932; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6957 = 7'h2c == rob_alloc_ids_3 ? 4'h0 : _GEN_5933; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6958 = 7'h2d == rob_alloc_ids_3 ? 4'h0 : _GEN_5934; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6959 = 7'h2e == rob_alloc_ids_3 ? 4'h0 : _GEN_5935; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6960 = 7'h2f == rob_alloc_ids_3 ? 4'h0 : _GEN_5936; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6961 = 7'h30 == rob_alloc_ids_3 ? 4'h0 : _GEN_5937; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6962 = 7'h31 == rob_alloc_ids_3 ? 4'h0 : _GEN_5938; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6963 = 7'h32 == rob_alloc_ids_3 ? 4'h0 : _GEN_5939; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6964 = 7'h33 == rob_alloc_ids_3 ? 4'h0 : _GEN_5940; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6965 = 7'h34 == rob_alloc_ids_3 ? 4'h0 : _GEN_5941; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6966 = 7'h35 == rob_alloc_ids_3 ? 4'h0 : _GEN_5942; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6967 = 7'h36 == rob_alloc_ids_3 ? 4'h0 : _GEN_5943; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6968 = 7'h37 == rob_alloc_ids_3 ? 4'h0 : _GEN_5944; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6969 = 7'h38 == rob_alloc_ids_3 ? 4'h0 : _GEN_5945; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6970 = 7'h39 == rob_alloc_ids_3 ? 4'h0 : _GEN_5946; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6971 = 7'h3a == rob_alloc_ids_3 ? 4'h0 : _GEN_5947; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6972 = 7'h3b == rob_alloc_ids_3 ? 4'h0 : _GEN_5948; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6973 = 7'h3c == rob_alloc_ids_3 ? 4'h0 : _GEN_5949; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6974 = 7'h3d == rob_alloc_ids_3 ? 4'h0 : _GEN_5950; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6975 = 7'h3e == rob_alloc_ids_3 ? 4'h0 : _GEN_5951; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6976 = 7'h3f == rob_alloc_ids_3 ? 4'h0 : _GEN_5952; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6977 = 7'h40 == rob_alloc_ids_3 ? 4'h0 : _GEN_5953; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6978 = 7'h41 == rob_alloc_ids_3 ? 4'h0 : _GEN_5954; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6979 = 7'h42 == rob_alloc_ids_3 ? 4'h0 : _GEN_5955; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6980 = 7'h43 == rob_alloc_ids_3 ? 4'h0 : _GEN_5956; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6981 = 7'h44 == rob_alloc_ids_3 ? 4'h0 : _GEN_5957; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6982 = 7'h45 == rob_alloc_ids_3 ? 4'h0 : _GEN_5958; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6983 = 7'h46 == rob_alloc_ids_3 ? 4'h0 : _GEN_5959; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6984 = 7'h47 == rob_alloc_ids_3 ? 4'h0 : _GEN_5960; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6985 = 7'h48 == rob_alloc_ids_3 ? 4'h0 : _GEN_5961; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6986 = 7'h49 == rob_alloc_ids_3 ? 4'h0 : _GEN_5962; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6987 = 7'h4a == rob_alloc_ids_3 ? 4'h0 : _GEN_5963; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6988 = 7'h4b == rob_alloc_ids_3 ? 4'h0 : _GEN_5964; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6989 = 7'h4c == rob_alloc_ids_3 ? 4'h0 : _GEN_5965; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6990 = 7'h4d == rob_alloc_ids_3 ? 4'h0 : _GEN_5966; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6991 = 7'h4e == rob_alloc_ids_3 ? 4'h0 : _GEN_5967; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6992 = 7'h4f == rob_alloc_ids_3 ? 4'h0 : _GEN_5968; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6993 = 7'h50 == rob_alloc_ids_3 ? 4'h0 : _GEN_5969; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6994 = 7'h51 == rob_alloc_ids_3 ? 4'h0 : _GEN_5970; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6995 = 7'h52 == rob_alloc_ids_3 ? 4'h0 : _GEN_5971; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6996 = 7'h53 == rob_alloc_ids_3 ? 4'h0 : _GEN_5972; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6997 = 7'h54 == rob_alloc_ids_3 ? 4'h0 : _GEN_5973; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6998 = 7'h55 == rob_alloc_ids_3 ? 4'h0 : _GEN_5974; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_6999 = 7'h56 == rob_alloc_ids_3 ? 4'h0 : _GEN_5975; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_7000 = 7'h57 == rob_alloc_ids_3 ? 4'h0 : _GEN_5976; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_7001 = 7'h58 == rob_alloc_ids_3 ? 4'h0 : _GEN_5977; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_7002 = 7'h59 == rob_alloc_ids_3 ? 4'h0 : _GEN_5978; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_7003 = 7'h5a == rob_alloc_ids_3 ? 4'h0 : _GEN_5979; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_7004 = 7'h5b == rob_alloc_ids_3 ? 4'h0 : _GEN_5980; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_7005 = 7'h5c == rob_alloc_ids_3 ? 4'h0 : _GEN_5981; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_7006 = 7'h5d == rob_alloc_ids_3 ? 4'h0 : _GEN_5982; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_7007 = 7'h5e == rob_alloc_ids_3 ? 4'h0 : _GEN_5983; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_7008 = 7'h5f == rob_alloc_ids_3 ? 4'h0 : _GEN_5984; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_7009 = 7'h60 == rob_alloc_ids_3 ? 4'h0 : _GEN_5985; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_7010 = 7'h61 == rob_alloc_ids_3 ? 4'h0 : _GEN_5986; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_7011 = 7'h62 == rob_alloc_ids_3 ? 4'h0 : _GEN_5987; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_7012 = 7'h63 == rob_alloc_ids_3 ? 4'h0 : _GEN_5988; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_7013 = 7'h64 == rob_alloc_ids_3 ? 4'h0 : _GEN_5989; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_7014 = 7'h65 == rob_alloc_ids_3 ? 4'h0 : _GEN_5990; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_7015 = 7'h66 == rob_alloc_ids_3 ? 4'h0 : _GEN_5991; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_7016 = 7'h67 == rob_alloc_ids_3 ? 4'h0 : _GEN_5992; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_7017 = 7'h68 == rob_alloc_ids_3 ? 4'h0 : _GEN_5993; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_7018 = 7'h69 == rob_alloc_ids_3 ? 4'h0 : _GEN_5994; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_7019 = 7'h6a == rob_alloc_ids_3 ? 4'h0 : _GEN_5995; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_7020 = 7'h6b == rob_alloc_ids_3 ? 4'h0 : _GEN_5996; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_7021 = 7'h6c == rob_alloc_ids_3 ? 4'h0 : _GEN_5997; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_7022 = 7'h6d == rob_alloc_ids_3 ? 4'h0 : _GEN_5998; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_7023 = 7'h6e == rob_alloc_ids_3 ? 4'h0 : _GEN_5999; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_7024 = 7'h6f == rob_alloc_ids_3 ? 4'h0 : _GEN_6000; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_7025 = 7'h70 == rob_alloc_ids_3 ? 4'h0 : _GEN_6001; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_7026 = 7'h71 == rob_alloc_ids_3 ? 4'h0 : _GEN_6002; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_7027 = 7'h72 == rob_alloc_ids_3 ? 4'h0 : _GEN_6003; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_7028 = 7'h73 == rob_alloc_ids_3 ? 4'h0 : _GEN_6004; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_7029 = 7'h74 == rob_alloc_ids_3 ? 4'h0 : _GEN_6005; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_7030 = 7'h75 == rob_alloc_ids_3 ? 4'h0 : _GEN_6006; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_7031 = 7'h76 == rob_alloc_ids_3 ? 4'h0 : _GEN_6007; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_7032 = 7'h77 == rob_alloc_ids_3 ? 4'h0 : _GEN_6008; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_7033 = 7'h78 == rob_alloc_ids_3 ? 4'h0 : _GEN_6009; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_7034 = 7'h79 == rob_alloc_ids_3 ? 4'h0 : _GEN_6010; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_7035 = 7'h7a == rob_alloc_ids_3 ? 4'h0 : _GEN_6011; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_7036 = 7'h7b == rob_alloc_ids_3 ? 4'h0 : _GEN_6012; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_7037 = 7'h7c == rob_alloc_ids_3 ? 4'h0 : _GEN_6013; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_7038 = 7'h7d == rob_alloc_ids_3 ? 4'h0 : _GEN_6014; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_7039 = 7'h7e == rob_alloc_ids_3 ? 4'h0 : _GEN_6015; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_7040 = 7'h7f == rob_alloc_ids_3 ? 4'h0 : _GEN_6016; // @[TestHarness.scala 183:{36,36}]
  wire [15:0] _GEN_7425 = igen_3_io_fire ? _GEN_6401 : _GEN_5377; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7426 = igen_3_io_fire ? _GEN_6402 : _GEN_5378; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7427 = igen_3_io_fire ? _GEN_6403 : _GEN_5379; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7428 = igen_3_io_fire ? _GEN_6404 : _GEN_5380; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7429 = igen_3_io_fire ? _GEN_6405 : _GEN_5381; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7430 = igen_3_io_fire ? _GEN_6406 : _GEN_5382; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7431 = igen_3_io_fire ? _GEN_6407 : _GEN_5383; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7432 = igen_3_io_fire ? _GEN_6408 : _GEN_5384; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7433 = igen_3_io_fire ? _GEN_6409 : _GEN_5385; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7434 = igen_3_io_fire ? _GEN_6410 : _GEN_5386; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7435 = igen_3_io_fire ? _GEN_6411 : _GEN_5387; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7436 = igen_3_io_fire ? _GEN_6412 : _GEN_5388; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7437 = igen_3_io_fire ? _GEN_6413 : _GEN_5389; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7438 = igen_3_io_fire ? _GEN_6414 : _GEN_5390; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7439 = igen_3_io_fire ? _GEN_6415 : _GEN_5391; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7440 = igen_3_io_fire ? _GEN_6416 : _GEN_5392; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7441 = igen_3_io_fire ? _GEN_6417 : _GEN_5393; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7442 = igen_3_io_fire ? _GEN_6418 : _GEN_5394; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7443 = igen_3_io_fire ? _GEN_6419 : _GEN_5395; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7444 = igen_3_io_fire ? _GEN_6420 : _GEN_5396; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7445 = igen_3_io_fire ? _GEN_6421 : _GEN_5397; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7446 = igen_3_io_fire ? _GEN_6422 : _GEN_5398; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7447 = igen_3_io_fire ? _GEN_6423 : _GEN_5399; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7448 = igen_3_io_fire ? _GEN_6424 : _GEN_5400; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7449 = igen_3_io_fire ? _GEN_6425 : _GEN_5401; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7450 = igen_3_io_fire ? _GEN_6426 : _GEN_5402; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7451 = igen_3_io_fire ? _GEN_6427 : _GEN_5403; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7452 = igen_3_io_fire ? _GEN_6428 : _GEN_5404; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7453 = igen_3_io_fire ? _GEN_6429 : _GEN_5405; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7454 = igen_3_io_fire ? _GEN_6430 : _GEN_5406; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7455 = igen_3_io_fire ? _GEN_6431 : _GEN_5407; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7456 = igen_3_io_fire ? _GEN_6432 : _GEN_5408; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7457 = igen_3_io_fire ? _GEN_6433 : _GEN_5409; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7458 = igen_3_io_fire ? _GEN_6434 : _GEN_5410; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7459 = igen_3_io_fire ? _GEN_6435 : _GEN_5411; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7460 = igen_3_io_fire ? _GEN_6436 : _GEN_5412; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7461 = igen_3_io_fire ? _GEN_6437 : _GEN_5413; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7462 = igen_3_io_fire ? _GEN_6438 : _GEN_5414; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7463 = igen_3_io_fire ? _GEN_6439 : _GEN_5415; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7464 = igen_3_io_fire ? _GEN_6440 : _GEN_5416; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7465 = igen_3_io_fire ? _GEN_6441 : _GEN_5417; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7466 = igen_3_io_fire ? _GEN_6442 : _GEN_5418; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7467 = igen_3_io_fire ? _GEN_6443 : _GEN_5419; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7468 = igen_3_io_fire ? _GEN_6444 : _GEN_5420; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7469 = igen_3_io_fire ? _GEN_6445 : _GEN_5421; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7470 = igen_3_io_fire ? _GEN_6446 : _GEN_5422; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7471 = igen_3_io_fire ? _GEN_6447 : _GEN_5423; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7472 = igen_3_io_fire ? _GEN_6448 : _GEN_5424; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7473 = igen_3_io_fire ? _GEN_6449 : _GEN_5425; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7474 = igen_3_io_fire ? _GEN_6450 : _GEN_5426; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7475 = igen_3_io_fire ? _GEN_6451 : _GEN_5427; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7476 = igen_3_io_fire ? _GEN_6452 : _GEN_5428; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7477 = igen_3_io_fire ? _GEN_6453 : _GEN_5429; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7478 = igen_3_io_fire ? _GEN_6454 : _GEN_5430; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7479 = igen_3_io_fire ? _GEN_6455 : _GEN_5431; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7480 = igen_3_io_fire ? _GEN_6456 : _GEN_5432; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7481 = igen_3_io_fire ? _GEN_6457 : _GEN_5433; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7482 = igen_3_io_fire ? _GEN_6458 : _GEN_5434; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7483 = igen_3_io_fire ? _GEN_6459 : _GEN_5435; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7484 = igen_3_io_fire ? _GEN_6460 : _GEN_5436; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7485 = igen_3_io_fire ? _GEN_6461 : _GEN_5437; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7486 = igen_3_io_fire ? _GEN_6462 : _GEN_5438; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7487 = igen_3_io_fire ? _GEN_6463 : _GEN_5439; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7488 = igen_3_io_fire ? _GEN_6464 : _GEN_5440; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7489 = igen_3_io_fire ? _GEN_6465 : _GEN_5441; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7490 = igen_3_io_fire ? _GEN_6466 : _GEN_5442; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7491 = igen_3_io_fire ? _GEN_6467 : _GEN_5443; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7492 = igen_3_io_fire ? _GEN_6468 : _GEN_5444; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7493 = igen_3_io_fire ? _GEN_6469 : _GEN_5445; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7494 = igen_3_io_fire ? _GEN_6470 : _GEN_5446; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7495 = igen_3_io_fire ? _GEN_6471 : _GEN_5447; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7496 = igen_3_io_fire ? _GEN_6472 : _GEN_5448; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7497 = igen_3_io_fire ? _GEN_6473 : _GEN_5449; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7498 = igen_3_io_fire ? _GEN_6474 : _GEN_5450; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7499 = igen_3_io_fire ? _GEN_6475 : _GEN_5451; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7500 = igen_3_io_fire ? _GEN_6476 : _GEN_5452; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7501 = igen_3_io_fire ? _GEN_6477 : _GEN_5453; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7502 = igen_3_io_fire ? _GEN_6478 : _GEN_5454; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7503 = igen_3_io_fire ? _GEN_6479 : _GEN_5455; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7504 = igen_3_io_fire ? _GEN_6480 : _GEN_5456; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7505 = igen_3_io_fire ? _GEN_6481 : _GEN_5457; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7506 = igen_3_io_fire ? _GEN_6482 : _GEN_5458; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7507 = igen_3_io_fire ? _GEN_6483 : _GEN_5459; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7508 = igen_3_io_fire ? _GEN_6484 : _GEN_5460; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7509 = igen_3_io_fire ? _GEN_6485 : _GEN_5461; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7510 = igen_3_io_fire ? _GEN_6486 : _GEN_5462; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7511 = igen_3_io_fire ? _GEN_6487 : _GEN_5463; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7512 = igen_3_io_fire ? _GEN_6488 : _GEN_5464; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7513 = igen_3_io_fire ? _GEN_6489 : _GEN_5465; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7514 = igen_3_io_fire ? _GEN_6490 : _GEN_5466; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7515 = igen_3_io_fire ? _GEN_6491 : _GEN_5467; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7516 = igen_3_io_fire ? _GEN_6492 : _GEN_5468; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7517 = igen_3_io_fire ? _GEN_6493 : _GEN_5469; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7518 = igen_3_io_fire ? _GEN_6494 : _GEN_5470; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7519 = igen_3_io_fire ? _GEN_6495 : _GEN_5471; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7520 = igen_3_io_fire ? _GEN_6496 : _GEN_5472; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7521 = igen_3_io_fire ? _GEN_6497 : _GEN_5473; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7522 = igen_3_io_fire ? _GEN_6498 : _GEN_5474; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7523 = igen_3_io_fire ? _GEN_6499 : _GEN_5475; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7524 = igen_3_io_fire ? _GEN_6500 : _GEN_5476; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7525 = igen_3_io_fire ? _GEN_6501 : _GEN_5477; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7526 = igen_3_io_fire ? _GEN_6502 : _GEN_5478; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7527 = igen_3_io_fire ? _GEN_6503 : _GEN_5479; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7528 = igen_3_io_fire ? _GEN_6504 : _GEN_5480; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7529 = igen_3_io_fire ? _GEN_6505 : _GEN_5481; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7530 = igen_3_io_fire ? _GEN_6506 : _GEN_5482; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7531 = igen_3_io_fire ? _GEN_6507 : _GEN_5483; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7532 = igen_3_io_fire ? _GEN_6508 : _GEN_5484; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7533 = igen_3_io_fire ? _GEN_6509 : _GEN_5485; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7534 = igen_3_io_fire ? _GEN_6510 : _GEN_5486; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7535 = igen_3_io_fire ? _GEN_6511 : _GEN_5487; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7536 = igen_3_io_fire ? _GEN_6512 : _GEN_5488; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7537 = igen_3_io_fire ? _GEN_6513 : _GEN_5489; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7538 = igen_3_io_fire ? _GEN_6514 : _GEN_5490; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7539 = igen_3_io_fire ? _GEN_6515 : _GEN_5491; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7540 = igen_3_io_fire ? _GEN_6516 : _GEN_5492; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7541 = igen_3_io_fire ? _GEN_6517 : _GEN_5493; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7542 = igen_3_io_fire ? _GEN_6518 : _GEN_5494; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7543 = igen_3_io_fire ? _GEN_6519 : _GEN_5495; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7544 = igen_3_io_fire ? _GEN_6520 : _GEN_5496; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7545 = igen_3_io_fire ? _GEN_6521 : _GEN_5497; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7546 = igen_3_io_fire ? _GEN_6522 : _GEN_5498; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7547 = igen_3_io_fire ? _GEN_6523 : _GEN_5499; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7548 = igen_3_io_fire ? _GEN_6524 : _GEN_5500; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7549 = igen_3_io_fire ? _GEN_6525 : _GEN_5501; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7550 = igen_3_io_fire ? _GEN_6526 : _GEN_5502; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7551 = igen_3_io_fire ? _GEN_6527 : _GEN_5503; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_7552 = igen_3_io_fire ? _GEN_6528 : _GEN_5504; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7937 = igen_3_io_fire ? _GEN_6913 : _GEN_5889; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7938 = igen_3_io_fire ? _GEN_6914 : _GEN_5890; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7939 = igen_3_io_fire ? _GEN_6915 : _GEN_5891; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7940 = igen_3_io_fire ? _GEN_6916 : _GEN_5892; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7941 = igen_3_io_fire ? _GEN_6917 : _GEN_5893; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7942 = igen_3_io_fire ? _GEN_6918 : _GEN_5894; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7943 = igen_3_io_fire ? _GEN_6919 : _GEN_5895; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7944 = igen_3_io_fire ? _GEN_6920 : _GEN_5896; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7945 = igen_3_io_fire ? _GEN_6921 : _GEN_5897; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7946 = igen_3_io_fire ? _GEN_6922 : _GEN_5898; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7947 = igen_3_io_fire ? _GEN_6923 : _GEN_5899; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7948 = igen_3_io_fire ? _GEN_6924 : _GEN_5900; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7949 = igen_3_io_fire ? _GEN_6925 : _GEN_5901; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7950 = igen_3_io_fire ? _GEN_6926 : _GEN_5902; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7951 = igen_3_io_fire ? _GEN_6927 : _GEN_5903; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7952 = igen_3_io_fire ? _GEN_6928 : _GEN_5904; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7953 = igen_3_io_fire ? _GEN_6929 : _GEN_5905; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7954 = igen_3_io_fire ? _GEN_6930 : _GEN_5906; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7955 = igen_3_io_fire ? _GEN_6931 : _GEN_5907; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7956 = igen_3_io_fire ? _GEN_6932 : _GEN_5908; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7957 = igen_3_io_fire ? _GEN_6933 : _GEN_5909; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7958 = igen_3_io_fire ? _GEN_6934 : _GEN_5910; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7959 = igen_3_io_fire ? _GEN_6935 : _GEN_5911; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7960 = igen_3_io_fire ? _GEN_6936 : _GEN_5912; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7961 = igen_3_io_fire ? _GEN_6937 : _GEN_5913; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7962 = igen_3_io_fire ? _GEN_6938 : _GEN_5914; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7963 = igen_3_io_fire ? _GEN_6939 : _GEN_5915; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7964 = igen_3_io_fire ? _GEN_6940 : _GEN_5916; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7965 = igen_3_io_fire ? _GEN_6941 : _GEN_5917; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7966 = igen_3_io_fire ? _GEN_6942 : _GEN_5918; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7967 = igen_3_io_fire ? _GEN_6943 : _GEN_5919; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7968 = igen_3_io_fire ? _GEN_6944 : _GEN_5920; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7969 = igen_3_io_fire ? _GEN_6945 : _GEN_5921; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7970 = igen_3_io_fire ? _GEN_6946 : _GEN_5922; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7971 = igen_3_io_fire ? _GEN_6947 : _GEN_5923; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7972 = igen_3_io_fire ? _GEN_6948 : _GEN_5924; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7973 = igen_3_io_fire ? _GEN_6949 : _GEN_5925; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7974 = igen_3_io_fire ? _GEN_6950 : _GEN_5926; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7975 = igen_3_io_fire ? _GEN_6951 : _GEN_5927; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7976 = igen_3_io_fire ? _GEN_6952 : _GEN_5928; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7977 = igen_3_io_fire ? _GEN_6953 : _GEN_5929; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7978 = igen_3_io_fire ? _GEN_6954 : _GEN_5930; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7979 = igen_3_io_fire ? _GEN_6955 : _GEN_5931; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7980 = igen_3_io_fire ? _GEN_6956 : _GEN_5932; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7981 = igen_3_io_fire ? _GEN_6957 : _GEN_5933; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7982 = igen_3_io_fire ? _GEN_6958 : _GEN_5934; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7983 = igen_3_io_fire ? _GEN_6959 : _GEN_5935; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7984 = igen_3_io_fire ? _GEN_6960 : _GEN_5936; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7985 = igen_3_io_fire ? _GEN_6961 : _GEN_5937; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7986 = igen_3_io_fire ? _GEN_6962 : _GEN_5938; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7987 = igen_3_io_fire ? _GEN_6963 : _GEN_5939; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7988 = igen_3_io_fire ? _GEN_6964 : _GEN_5940; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7989 = igen_3_io_fire ? _GEN_6965 : _GEN_5941; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7990 = igen_3_io_fire ? _GEN_6966 : _GEN_5942; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7991 = igen_3_io_fire ? _GEN_6967 : _GEN_5943; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7992 = igen_3_io_fire ? _GEN_6968 : _GEN_5944; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7993 = igen_3_io_fire ? _GEN_6969 : _GEN_5945; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7994 = igen_3_io_fire ? _GEN_6970 : _GEN_5946; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7995 = igen_3_io_fire ? _GEN_6971 : _GEN_5947; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7996 = igen_3_io_fire ? _GEN_6972 : _GEN_5948; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7997 = igen_3_io_fire ? _GEN_6973 : _GEN_5949; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7998 = igen_3_io_fire ? _GEN_6974 : _GEN_5950; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_7999 = igen_3_io_fire ? _GEN_6975 : _GEN_5951; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8000 = igen_3_io_fire ? _GEN_6976 : _GEN_5952; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8001 = igen_3_io_fire ? _GEN_6977 : _GEN_5953; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8002 = igen_3_io_fire ? _GEN_6978 : _GEN_5954; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8003 = igen_3_io_fire ? _GEN_6979 : _GEN_5955; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8004 = igen_3_io_fire ? _GEN_6980 : _GEN_5956; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8005 = igen_3_io_fire ? _GEN_6981 : _GEN_5957; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8006 = igen_3_io_fire ? _GEN_6982 : _GEN_5958; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8007 = igen_3_io_fire ? _GEN_6983 : _GEN_5959; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8008 = igen_3_io_fire ? _GEN_6984 : _GEN_5960; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8009 = igen_3_io_fire ? _GEN_6985 : _GEN_5961; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8010 = igen_3_io_fire ? _GEN_6986 : _GEN_5962; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8011 = igen_3_io_fire ? _GEN_6987 : _GEN_5963; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8012 = igen_3_io_fire ? _GEN_6988 : _GEN_5964; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8013 = igen_3_io_fire ? _GEN_6989 : _GEN_5965; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8014 = igen_3_io_fire ? _GEN_6990 : _GEN_5966; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8015 = igen_3_io_fire ? _GEN_6991 : _GEN_5967; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8016 = igen_3_io_fire ? _GEN_6992 : _GEN_5968; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8017 = igen_3_io_fire ? _GEN_6993 : _GEN_5969; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8018 = igen_3_io_fire ? _GEN_6994 : _GEN_5970; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8019 = igen_3_io_fire ? _GEN_6995 : _GEN_5971; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8020 = igen_3_io_fire ? _GEN_6996 : _GEN_5972; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8021 = igen_3_io_fire ? _GEN_6997 : _GEN_5973; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8022 = igen_3_io_fire ? _GEN_6998 : _GEN_5974; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8023 = igen_3_io_fire ? _GEN_6999 : _GEN_5975; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8024 = igen_3_io_fire ? _GEN_7000 : _GEN_5976; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8025 = igen_3_io_fire ? _GEN_7001 : _GEN_5977; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8026 = igen_3_io_fire ? _GEN_7002 : _GEN_5978; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8027 = igen_3_io_fire ? _GEN_7003 : _GEN_5979; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8028 = igen_3_io_fire ? _GEN_7004 : _GEN_5980; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8029 = igen_3_io_fire ? _GEN_7005 : _GEN_5981; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8030 = igen_3_io_fire ? _GEN_7006 : _GEN_5982; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8031 = igen_3_io_fire ? _GEN_7007 : _GEN_5983; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8032 = igen_3_io_fire ? _GEN_7008 : _GEN_5984; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8033 = igen_3_io_fire ? _GEN_7009 : _GEN_5985; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8034 = igen_3_io_fire ? _GEN_7010 : _GEN_5986; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8035 = igen_3_io_fire ? _GEN_7011 : _GEN_5987; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8036 = igen_3_io_fire ? _GEN_7012 : _GEN_5988; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8037 = igen_3_io_fire ? _GEN_7013 : _GEN_5989; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8038 = igen_3_io_fire ? _GEN_7014 : _GEN_5990; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8039 = igen_3_io_fire ? _GEN_7015 : _GEN_5991; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8040 = igen_3_io_fire ? _GEN_7016 : _GEN_5992; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8041 = igen_3_io_fire ? _GEN_7017 : _GEN_5993; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8042 = igen_3_io_fire ? _GEN_7018 : _GEN_5994; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8043 = igen_3_io_fire ? _GEN_7019 : _GEN_5995; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8044 = igen_3_io_fire ? _GEN_7020 : _GEN_5996; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8045 = igen_3_io_fire ? _GEN_7021 : _GEN_5997; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8046 = igen_3_io_fire ? _GEN_7022 : _GEN_5998; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8047 = igen_3_io_fire ? _GEN_7023 : _GEN_5999; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8048 = igen_3_io_fire ? _GEN_7024 : _GEN_6000; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8049 = igen_3_io_fire ? _GEN_7025 : _GEN_6001; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8050 = igen_3_io_fire ? _GEN_7026 : _GEN_6002; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8051 = igen_3_io_fire ? _GEN_7027 : _GEN_6003; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8052 = igen_3_io_fire ? _GEN_7028 : _GEN_6004; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8053 = igen_3_io_fire ? _GEN_7029 : _GEN_6005; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8054 = igen_3_io_fire ? _GEN_7030 : _GEN_6006; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8055 = igen_3_io_fire ? _GEN_7031 : _GEN_6007; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8056 = igen_3_io_fire ? _GEN_7032 : _GEN_6008; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8057 = igen_3_io_fire ? _GEN_7033 : _GEN_6009; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8058 = igen_3_io_fire ? _GEN_7034 : _GEN_6010; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8059 = igen_3_io_fire ? _GEN_7035 : _GEN_6011; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8060 = igen_3_io_fire ? _GEN_7036 : _GEN_6012; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8061 = igen_3_io_fire ? _GEN_7037 : _GEN_6013; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8062 = igen_3_io_fire ? _GEN_7038 : _GEN_6014; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8063 = igen_3_io_fire ? _GEN_7039 : _GEN_6015; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_8064 = igen_3_io_fire ? _GEN_7040 : _GEN_6016; // @[TestHarness.scala 178:25]
  wire  enable_print_latency = plusarg_reader_out; // @[TestHarness.scala 190:81]
  wire [31:0] out_payload_tsc = io_from_noc_0_flit_bits_payload[63:32]; // @[TestHarness.scala 194:51]
  reg  packet_valid; // @[TestHarness.scala 196:31]
  reg [6:0] packet_rob_idx; // @[TestHarness.scala 197:29]
  wire [127:0] _T_76 = rob_valids >> out_payload_rob_idx; // @[TestHarness.scala 201:24]
  wire [31:0] _GEN_8194 = 7'h1 == out_payload_rob_idx[6:0] ? rob_payload_1_tsc : rob_payload_0_tsc; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8195 = 7'h2 == out_payload_rob_idx[6:0] ? rob_payload_2_tsc : _GEN_8194; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8196 = 7'h3 == out_payload_rob_idx[6:0] ? rob_payload_3_tsc : _GEN_8195; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8197 = 7'h4 == out_payload_rob_idx[6:0] ? rob_payload_4_tsc : _GEN_8196; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8198 = 7'h5 == out_payload_rob_idx[6:0] ? rob_payload_5_tsc : _GEN_8197; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8199 = 7'h6 == out_payload_rob_idx[6:0] ? rob_payload_6_tsc : _GEN_8198; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8200 = 7'h7 == out_payload_rob_idx[6:0] ? rob_payload_7_tsc : _GEN_8199; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8201 = 7'h8 == out_payload_rob_idx[6:0] ? rob_payload_8_tsc : _GEN_8200; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8202 = 7'h9 == out_payload_rob_idx[6:0] ? rob_payload_9_tsc : _GEN_8201; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8203 = 7'ha == out_payload_rob_idx[6:0] ? rob_payload_10_tsc : _GEN_8202; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8204 = 7'hb == out_payload_rob_idx[6:0] ? rob_payload_11_tsc : _GEN_8203; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8205 = 7'hc == out_payload_rob_idx[6:0] ? rob_payload_12_tsc : _GEN_8204; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8206 = 7'hd == out_payload_rob_idx[6:0] ? rob_payload_13_tsc : _GEN_8205; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8207 = 7'he == out_payload_rob_idx[6:0] ? rob_payload_14_tsc : _GEN_8206; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8208 = 7'hf == out_payload_rob_idx[6:0] ? rob_payload_15_tsc : _GEN_8207; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8209 = 7'h10 == out_payload_rob_idx[6:0] ? rob_payload_16_tsc : _GEN_8208; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8210 = 7'h11 == out_payload_rob_idx[6:0] ? rob_payload_17_tsc : _GEN_8209; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8211 = 7'h12 == out_payload_rob_idx[6:0] ? rob_payload_18_tsc : _GEN_8210; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8212 = 7'h13 == out_payload_rob_idx[6:0] ? rob_payload_19_tsc : _GEN_8211; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8213 = 7'h14 == out_payload_rob_idx[6:0] ? rob_payload_20_tsc : _GEN_8212; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8214 = 7'h15 == out_payload_rob_idx[6:0] ? rob_payload_21_tsc : _GEN_8213; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8215 = 7'h16 == out_payload_rob_idx[6:0] ? rob_payload_22_tsc : _GEN_8214; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8216 = 7'h17 == out_payload_rob_idx[6:0] ? rob_payload_23_tsc : _GEN_8215; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8217 = 7'h18 == out_payload_rob_idx[6:0] ? rob_payload_24_tsc : _GEN_8216; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8218 = 7'h19 == out_payload_rob_idx[6:0] ? rob_payload_25_tsc : _GEN_8217; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8219 = 7'h1a == out_payload_rob_idx[6:0] ? rob_payload_26_tsc : _GEN_8218; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8220 = 7'h1b == out_payload_rob_idx[6:0] ? rob_payload_27_tsc : _GEN_8219; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8221 = 7'h1c == out_payload_rob_idx[6:0] ? rob_payload_28_tsc : _GEN_8220; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8222 = 7'h1d == out_payload_rob_idx[6:0] ? rob_payload_29_tsc : _GEN_8221; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8223 = 7'h1e == out_payload_rob_idx[6:0] ? rob_payload_30_tsc : _GEN_8222; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8224 = 7'h1f == out_payload_rob_idx[6:0] ? rob_payload_31_tsc : _GEN_8223; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8225 = 7'h20 == out_payload_rob_idx[6:0] ? rob_payload_32_tsc : _GEN_8224; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8226 = 7'h21 == out_payload_rob_idx[6:0] ? rob_payload_33_tsc : _GEN_8225; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8227 = 7'h22 == out_payload_rob_idx[6:0] ? rob_payload_34_tsc : _GEN_8226; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8228 = 7'h23 == out_payload_rob_idx[6:0] ? rob_payload_35_tsc : _GEN_8227; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8229 = 7'h24 == out_payload_rob_idx[6:0] ? rob_payload_36_tsc : _GEN_8228; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8230 = 7'h25 == out_payload_rob_idx[6:0] ? rob_payload_37_tsc : _GEN_8229; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8231 = 7'h26 == out_payload_rob_idx[6:0] ? rob_payload_38_tsc : _GEN_8230; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8232 = 7'h27 == out_payload_rob_idx[6:0] ? rob_payload_39_tsc : _GEN_8231; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8233 = 7'h28 == out_payload_rob_idx[6:0] ? rob_payload_40_tsc : _GEN_8232; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8234 = 7'h29 == out_payload_rob_idx[6:0] ? rob_payload_41_tsc : _GEN_8233; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8235 = 7'h2a == out_payload_rob_idx[6:0] ? rob_payload_42_tsc : _GEN_8234; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8236 = 7'h2b == out_payload_rob_idx[6:0] ? rob_payload_43_tsc : _GEN_8235; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8237 = 7'h2c == out_payload_rob_idx[6:0] ? rob_payload_44_tsc : _GEN_8236; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8238 = 7'h2d == out_payload_rob_idx[6:0] ? rob_payload_45_tsc : _GEN_8237; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8239 = 7'h2e == out_payload_rob_idx[6:0] ? rob_payload_46_tsc : _GEN_8238; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8240 = 7'h2f == out_payload_rob_idx[6:0] ? rob_payload_47_tsc : _GEN_8239; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8241 = 7'h30 == out_payload_rob_idx[6:0] ? rob_payload_48_tsc : _GEN_8240; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8242 = 7'h31 == out_payload_rob_idx[6:0] ? rob_payload_49_tsc : _GEN_8241; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8243 = 7'h32 == out_payload_rob_idx[6:0] ? rob_payload_50_tsc : _GEN_8242; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8244 = 7'h33 == out_payload_rob_idx[6:0] ? rob_payload_51_tsc : _GEN_8243; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8245 = 7'h34 == out_payload_rob_idx[6:0] ? rob_payload_52_tsc : _GEN_8244; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8246 = 7'h35 == out_payload_rob_idx[6:0] ? rob_payload_53_tsc : _GEN_8245; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8247 = 7'h36 == out_payload_rob_idx[6:0] ? rob_payload_54_tsc : _GEN_8246; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8248 = 7'h37 == out_payload_rob_idx[6:0] ? rob_payload_55_tsc : _GEN_8247; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8249 = 7'h38 == out_payload_rob_idx[6:0] ? rob_payload_56_tsc : _GEN_8248; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8250 = 7'h39 == out_payload_rob_idx[6:0] ? rob_payload_57_tsc : _GEN_8249; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8251 = 7'h3a == out_payload_rob_idx[6:0] ? rob_payload_58_tsc : _GEN_8250; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8252 = 7'h3b == out_payload_rob_idx[6:0] ? rob_payload_59_tsc : _GEN_8251; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8253 = 7'h3c == out_payload_rob_idx[6:0] ? rob_payload_60_tsc : _GEN_8252; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8254 = 7'h3d == out_payload_rob_idx[6:0] ? rob_payload_61_tsc : _GEN_8253; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8255 = 7'h3e == out_payload_rob_idx[6:0] ? rob_payload_62_tsc : _GEN_8254; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8256 = 7'h3f == out_payload_rob_idx[6:0] ? rob_payload_63_tsc : _GEN_8255; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8257 = 7'h40 == out_payload_rob_idx[6:0] ? rob_payload_64_tsc : _GEN_8256; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8258 = 7'h41 == out_payload_rob_idx[6:0] ? rob_payload_65_tsc : _GEN_8257; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8259 = 7'h42 == out_payload_rob_idx[6:0] ? rob_payload_66_tsc : _GEN_8258; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8260 = 7'h43 == out_payload_rob_idx[6:0] ? rob_payload_67_tsc : _GEN_8259; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8261 = 7'h44 == out_payload_rob_idx[6:0] ? rob_payload_68_tsc : _GEN_8260; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8262 = 7'h45 == out_payload_rob_idx[6:0] ? rob_payload_69_tsc : _GEN_8261; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8263 = 7'h46 == out_payload_rob_idx[6:0] ? rob_payload_70_tsc : _GEN_8262; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8264 = 7'h47 == out_payload_rob_idx[6:0] ? rob_payload_71_tsc : _GEN_8263; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8265 = 7'h48 == out_payload_rob_idx[6:0] ? rob_payload_72_tsc : _GEN_8264; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8266 = 7'h49 == out_payload_rob_idx[6:0] ? rob_payload_73_tsc : _GEN_8265; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8267 = 7'h4a == out_payload_rob_idx[6:0] ? rob_payload_74_tsc : _GEN_8266; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8268 = 7'h4b == out_payload_rob_idx[6:0] ? rob_payload_75_tsc : _GEN_8267; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8269 = 7'h4c == out_payload_rob_idx[6:0] ? rob_payload_76_tsc : _GEN_8268; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8270 = 7'h4d == out_payload_rob_idx[6:0] ? rob_payload_77_tsc : _GEN_8269; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8271 = 7'h4e == out_payload_rob_idx[6:0] ? rob_payload_78_tsc : _GEN_8270; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8272 = 7'h4f == out_payload_rob_idx[6:0] ? rob_payload_79_tsc : _GEN_8271; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8273 = 7'h50 == out_payload_rob_idx[6:0] ? rob_payload_80_tsc : _GEN_8272; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8274 = 7'h51 == out_payload_rob_idx[6:0] ? rob_payload_81_tsc : _GEN_8273; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8275 = 7'h52 == out_payload_rob_idx[6:0] ? rob_payload_82_tsc : _GEN_8274; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8276 = 7'h53 == out_payload_rob_idx[6:0] ? rob_payload_83_tsc : _GEN_8275; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8277 = 7'h54 == out_payload_rob_idx[6:0] ? rob_payload_84_tsc : _GEN_8276; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8278 = 7'h55 == out_payload_rob_idx[6:0] ? rob_payload_85_tsc : _GEN_8277; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8279 = 7'h56 == out_payload_rob_idx[6:0] ? rob_payload_86_tsc : _GEN_8278; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8280 = 7'h57 == out_payload_rob_idx[6:0] ? rob_payload_87_tsc : _GEN_8279; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8281 = 7'h58 == out_payload_rob_idx[6:0] ? rob_payload_88_tsc : _GEN_8280; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8282 = 7'h59 == out_payload_rob_idx[6:0] ? rob_payload_89_tsc : _GEN_8281; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8283 = 7'h5a == out_payload_rob_idx[6:0] ? rob_payload_90_tsc : _GEN_8282; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8284 = 7'h5b == out_payload_rob_idx[6:0] ? rob_payload_91_tsc : _GEN_8283; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8285 = 7'h5c == out_payload_rob_idx[6:0] ? rob_payload_92_tsc : _GEN_8284; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8286 = 7'h5d == out_payload_rob_idx[6:0] ? rob_payload_93_tsc : _GEN_8285; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8287 = 7'h5e == out_payload_rob_idx[6:0] ? rob_payload_94_tsc : _GEN_8286; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8288 = 7'h5f == out_payload_rob_idx[6:0] ? rob_payload_95_tsc : _GEN_8287; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8289 = 7'h60 == out_payload_rob_idx[6:0] ? rob_payload_96_tsc : _GEN_8288; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8290 = 7'h61 == out_payload_rob_idx[6:0] ? rob_payload_97_tsc : _GEN_8289; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8291 = 7'h62 == out_payload_rob_idx[6:0] ? rob_payload_98_tsc : _GEN_8290; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8292 = 7'h63 == out_payload_rob_idx[6:0] ? rob_payload_99_tsc : _GEN_8291; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8293 = 7'h64 == out_payload_rob_idx[6:0] ? rob_payload_100_tsc : _GEN_8292; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8294 = 7'h65 == out_payload_rob_idx[6:0] ? rob_payload_101_tsc : _GEN_8293; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8295 = 7'h66 == out_payload_rob_idx[6:0] ? rob_payload_102_tsc : _GEN_8294; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8296 = 7'h67 == out_payload_rob_idx[6:0] ? rob_payload_103_tsc : _GEN_8295; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8297 = 7'h68 == out_payload_rob_idx[6:0] ? rob_payload_104_tsc : _GEN_8296; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8298 = 7'h69 == out_payload_rob_idx[6:0] ? rob_payload_105_tsc : _GEN_8297; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8299 = 7'h6a == out_payload_rob_idx[6:0] ? rob_payload_106_tsc : _GEN_8298; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8300 = 7'h6b == out_payload_rob_idx[6:0] ? rob_payload_107_tsc : _GEN_8299; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8301 = 7'h6c == out_payload_rob_idx[6:0] ? rob_payload_108_tsc : _GEN_8300; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8302 = 7'h6d == out_payload_rob_idx[6:0] ? rob_payload_109_tsc : _GEN_8301; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8303 = 7'h6e == out_payload_rob_idx[6:0] ? rob_payload_110_tsc : _GEN_8302; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8304 = 7'h6f == out_payload_rob_idx[6:0] ? rob_payload_111_tsc : _GEN_8303; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8305 = 7'h70 == out_payload_rob_idx[6:0] ? rob_payload_112_tsc : _GEN_8304; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8306 = 7'h71 == out_payload_rob_idx[6:0] ? rob_payload_113_tsc : _GEN_8305; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8307 = 7'h72 == out_payload_rob_idx[6:0] ? rob_payload_114_tsc : _GEN_8306; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8308 = 7'h73 == out_payload_rob_idx[6:0] ? rob_payload_115_tsc : _GEN_8307; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8309 = 7'h74 == out_payload_rob_idx[6:0] ? rob_payload_116_tsc : _GEN_8308; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8310 = 7'h75 == out_payload_rob_idx[6:0] ? rob_payload_117_tsc : _GEN_8309; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8311 = 7'h76 == out_payload_rob_idx[6:0] ? rob_payload_118_tsc : _GEN_8310; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8312 = 7'h77 == out_payload_rob_idx[6:0] ? rob_payload_119_tsc : _GEN_8311; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8313 = 7'h78 == out_payload_rob_idx[6:0] ? rob_payload_120_tsc : _GEN_8312; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8314 = 7'h79 == out_payload_rob_idx[6:0] ? rob_payload_121_tsc : _GEN_8313; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8315 = 7'h7a == out_payload_rob_idx[6:0] ? rob_payload_122_tsc : _GEN_8314; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8316 = 7'h7b == out_payload_rob_idx[6:0] ? rob_payload_123_tsc : _GEN_8315; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8317 = 7'h7c == out_payload_rob_idx[6:0] ? rob_payload_124_tsc : _GEN_8316; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8318 = 7'h7d == out_payload_rob_idx[6:0] ? rob_payload_125_tsc : _GEN_8317; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8319 = 7'h7e == out_payload_rob_idx[6:0] ? rob_payload_126_tsc : _GEN_8318; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_8320 = 7'h7f == out_payload_rob_idx[6:0] ? rob_payload_127_tsc : _GEN_8319; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8322 = 7'h1 == out_payload_rob_idx[6:0] ? rob_payload_1_rob_idx : rob_payload_0_rob_idx; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8323 = 7'h2 == out_payload_rob_idx[6:0] ? rob_payload_2_rob_idx : _GEN_8322; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8324 = 7'h3 == out_payload_rob_idx[6:0] ? rob_payload_3_rob_idx : _GEN_8323; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8325 = 7'h4 == out_payload_rob_idx[6:0] ? rob_payload_4_rob_idx : _GEN_8324; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8326 = 7'h5 == out_payload_rob_idx[6:0] ? rob_payload_5_rob_idx : _GEN_8325; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8327 = 7'h6 == out_payload_rob_idx[6:0] ? rob_payload_6_rob_idx : _GEN_8326; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8328 = 7'h7 == out_payload_rob_idx[6:0] ? rob_payload_7_rob_idx : _GEN_8327; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8329 = 7'h8 == out_payload_rob_idx[6:0] ? rob_payload_8_rob_idx : _GEN_8328; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8330 = 7'h9 == out_payload_rob_idx[6:0] ? rob_payload_9_rob_idx : _GEN_8329; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8331 = 7'ha == out_payload_rob_idx[6:0] ? rob_payload_10_rob_idx : _GEN_8330; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8332 = 7'hb == out_payload_rob_idx[6:0] ? rob_payload_11_rob_idx : _GEN_8331; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8333 = 7'hc == out_payload_rob_idx[6:0] ? rob_payload_12_rob_idx : _GEN_8332; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8334 = 7'hd == out_payload_rob_idx[6:0] ? rob_payload_13_rob_idx : _GEN_8333; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8335 = 7'he == out_payload_rob_idx[6:0] ? rob_payload_14_rob_idx : _GEN_8334; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8336 = 7'hf == out_payload_rob_idx[6:0] ? rob_payload_15_rob_idx : _GEN_8335; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8337 = 7'h10 == out_payload_rob_idx[6:0] ? rob_payload_16_rob_idx : _GEN_8336; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8338 = 7'h11 == out_payload_rob_idx[6:0] ? rob_payload_17_rob_idx : _GEN_8337; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8339 = 7'h12 == out_payload_rob_idx[6:0] ? rob_payload_18_rob_idx : _GEN_8338; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8340 = 7'h13 == out_payload_rob_idx[6:0] ? rob_payload_19_rob_idx : _GEN_8339; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8341 = 7'h14 == out_payload_rob_idx[6:0] ? rob_payload_20_rob_idx : _GEN_8340; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8342 = 7'h15 == out_payload_rob_idx[6:0] ? rob_payload_21_rob_idx : _GEN_8341; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8343 = 7'h16 == out_payload_rob_idx[6:0] ? rob_payload_22_rob_idx : _GEN_8342; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8344 = 7'h17 == out_payload_rob_idx[6:0] ? rob_payload_23_rob_idx : _GEN_8343; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8345 = 7'h18 == out_payload_rob_idx[6:0] ? rob_payload_24_rob_idx : _GEN_8344; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8346 = 7'h19 == out_payload_rob_idx[6:0] ? rob_payload_25_rob_idx : _GEN_8345; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8347 = 7'h1a == out_payload_rob_idx[6:0] ? rob_payload_26_rob_idx : _GEN_8346; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8348 = 7'h1b == out_payload_rob_idx[6:0] ? rob_payload_27_rob_idx : _GEN_8347; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8349 = 7'h1c == out_payload_rob_idx[6:0] ? rob_payload_28_rob_idx : _GEN_8348; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8350 = 7'h1d == out_payload_rob_idx[6:0] ? rob_payload_29_rob_idx : _GEN_8349; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8351 = 7'h1e == out_payload_rob_idx[6:0] ? rob_payload_30_rob_idx : _GEN_8350; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8352 = 7'h1f == out_payload_rob_idx[6:0] ? rob_payload_31_rob_idx : _GEN_8351; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8353 = 7'h20 == out_payload_rob_idx[6:0] ? rob_payload_32_rob_idx : _GEN_8352; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8354 = 7'h21 == out_payload_rob_idx[6:0] ? rob_payload_33_rob_idx : _GEN_8353; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8355 = 7'h22 == out_payload_rob_idx[6:0] ? rob_payload_34_rob_idx : _GEN_8354; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8356 = 7'h23 == out_payload_rob_idx[6:0] ? rob_payload_35_rob_idx : _GEN_8355; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8357 = 7'h24 == out_payload_rob_idx[6:0] ? rob_payload_36_rob_idx : _GEN_8356; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8358 = 7'h25 == out_payload_rob_idx[6:0] ? rob_payload_37_rob_idx : _GEN_8357; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8359 = 7'h26 == out_payload_rob_idx[6:0] ? rob_payload_38_rob_idx : _GEN_8358; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8360 = 7'h27 == out_payload_rob_idx[6:0] ? rob_payload_39_rob_idx : _GEN_8359; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8361 = 7'h28 == out_payload_rob_idx[6:0] ? rob_payload_40_rob_idx : _GEN_8360; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8362 = 7'h29 == out_payload_rob_idx[6:0] ? rob_payload_41_rob_idx : _GEN_8361; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8363 = 7'h2a == out_payload_rob_idx[6:0] ? rob_payload_42_rob_idx : _GEN_8362; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8364 = 7'h2b == out_payload_rob_idx[6:0] ? rob_payload_43_rob_idx : _GEN_8363; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8365 = 7'h2c == out_payload_rob_idx[6:0] ? rob_payload_44_rob_idx : _GEN_8364; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8366 = 7'h2d == out_payload_rob_idx[6:0] ? rob_payload_45_rob_idx : _GEN_8365; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8367 = 7'h2e == out_payload_rob_idx[6:0] ? rob_payload_46_rob_idx : _GEN_8366; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8368 = 7'h2f == out_payload_rob_idx[6:0] ? rob_payload_47_rob_idx : _GEN_8367; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8369 = 7'h30 == out_payload_rob_idx[6:0] ? rob_payload_48_rob_idx : _GEN_8368; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8370 = 7'h31 == out_payload_rob_idx[6:0] ? rob_payload_49_rob_idx : _GEN_8369; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8371 = 7'h32 == out_payload_rob_idx[6:0] ? rob_payload_50_rob_idx : _GEN_8370; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8372 = 7'h33 == out_payload_rob_idx[6:0] ? rob_payload_51_rob_idx : _GEN_8371; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8373 = 7'h34 == out_payload_rob_idx[6:0] ? rob_payload_52_rob_idx : _GEN_8372; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8374 = 7'h35 == out_payload_rob_idx[6:0] ? rob_payload_53_rob_idx : _GEN_8373; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8375 = 7'h36 == out_payload_rob_idx[6:0] ? rob_payload_54_rob_idx : _GEN_8374; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8376 = 7'h37 == out_payload_rob_idx[6:0] ? rob_payload_55_rob_idx : _GEN_8375; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8377 = 7'h38 == out_payload_rob_idx[6:0] ? rob_payload_56_rob_idx : _GEN_8376; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8378 = 7'h39 == out_payload_rob_idx[6:0] ? rob_payload_57_rob_idx : _GEN_8377; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8379 = 7'h3a == out_payload_rob_idx[6:0] ? rob_payload_58_rob_idx : _GEN_8378; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8380 = 7'h3b == out_payload_rob_idx[6:0] ? rob_payload_59_rob_idx : _GEN_8379; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8381 = 7'h3c == out_payload_rob_idx[6:0] ? rob_payload_60_rob_idx : _GEN_8380; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8382 = 7'h3d == out_payload_rob_idx[6:0] ? rob_payload_61_rob_idx : _GEN_8381; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8383 = 7'h3e == out_payload_rob_idx[6:0] ? rob_payload_62_rob_idx : _GEN_8382; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8384 = 7'h3f == out_payload_rob_idx[6:0] ? rob_payload_63_rob_idx : _GEN_8383; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8385 = 7'h40 == out_payload_rob_idx[6:0] ? rob_payload_64_rob_idx : _GEN_8384; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8386 = 7'h41 == out_payload_rob_idx[6:0] ? rob_payload_65_rob_idx : _GEN_8385; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8387 = 7'h42 == out_payload_rob_idx[6:0] ? rob_payload_66_rob_idx : _GEN_8386; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8388 = 7'h43 == out_payload_rob_idx[6:0] ? rob_payload_67_rob_idx : _GEN_8387; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8389 = 7'h44 == out_payload_rob_idx[6:0] ? rob_payload_68_rob_idx : _GEN_8388; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8390 = 7'h45 == out_payload_rob_idx[6:0] ? rob_payload_69_rob_idx : _GEN_8389; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8391 = 7'h46 == out_payload_rob_idx[6:0] ? rob_payload_70_rob_idx : _GEN_8390; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8392 = 7'h47 == out_payload_rob_idx[6:0] ? rob_payload_71_rob_idx : _GEN_8391; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8393 = 7'h48 == out_payload_rob_idx[6:0] ? rob_payload_72_rob_idx : _GEN_8392; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8394 = 7'h49 == out_payload_rob_idx[6:0] ? rob_payload_73_rob_idx : _GEN_8393; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8395 = 7'h4a == out_payload_rob_idx[6:0] ? rob_payload_74_rob_idx : _GEN_8394; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8396 = 7'h4b == out_payload_rob_idx[6:0] ? rob_payload_75_rob_idx : _GEN_8395; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8397 = 7'h4c == out_payload_rob_idx[6:0] ? rob_payload_76_rob_idx : _GEN_8396; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8398 = 7'h4d == out_payload_rob_idx[6:0] ? rob_payload_77_rob_idx : _GEN_8397; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8399 = 7'h4e == out_payload_rob_idx[6:0] ? rob_payload_78_rob_idx : _GEN_8398; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8400 = 7'h4f == out_payload_rob_idx[6:0] ? rob_payload_79_rob_idx : _GEN_8399; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8401 = 7'h50 == out_payload_rob_idx[6:0] ? rob_payload_80_rob_idx : _GEN_8400; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8402 = 7'h51 == out_payload_rob_idx[6:0] ? rob_payload_81_rob_idx : _GEN_8401; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8403 = 7'h52 == out_payload_rob_idx[6:0] ? rob_payload_82_rob_idx : _GEN_8402; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8404 = 7'h53 == out_payload_rob_idx[6:0] ? rob_payload_83_rob_idx : _GEN_8403; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8405 = 7'h54 == out_payload_rob_idx[6:0] ? rob_payload_84_rob_idx : _GEN_8404; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8406 = 7'h55 == out_payload_rob_idx[6:0] ? rob_payload_85_rob_idx : _GEN_8405; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8407 = 7'h56 == out_payload_rob_idx[6:0] ? rob_payload_86_rob_idx : _GEN_8406; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8408 = 7'h57 == out_payload_rob_idx[6:0] ? rob_payload_87_rob_idx : _GEN_8407; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8409 = 7'h58 == out_payload_rob_idx[6:0] ? rob_payload_88_rob_idx : _GEN_8408; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8410 = 7'h59 == out_payload_rob_idx[6:0] ? rob_payload_89_rob_idx : _GEN_8409; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8411 = 7'h5a == out_payload_rob_idx[6:0] ? rob_payload_90_rob_idx : _GEN_8410; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8412 = 7'h5b == out_payload_rob_idx[6:0] ? rob_payload_91_rob_idx : _GEN_8411; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8413 = 7'h5c == out_payload_rob_idx[6:0] ? rob_payload_92_rob_idx : _GEN_8412; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8414 = 7'h5d == out_payload_rob_idx[6:0] ? rob_payload_93_rob_idx : _GEN_8413; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8415 = 7'h5e == out_payload_rob_idx[6:0] ? rob_payload_94_rob_idx : _GEN_8414; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8416 = 7'h5f == out_payload_rob_idx[6:0] ? rob_payload_95_rob_idx : _GEN_8415; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8417 = 7'h60 == out_payload_rob_idx[6:0] ? rob_payload_96_rob_idx : _GEN_8416; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8418 = 7'h61 == out_payload_rob_idx[6:0] ? rob_payload_97_rob_idx : _GEN_8417; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8419 = 7'h62 == out_payload_rob_idx[6:0] ? rob_payload_98_rob_idx : _GEN_8418; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8420 = 7'h63 == out_payload_rob_idx[6:0] ? rob_payload_99_rob_idx : _GEN_8419; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8421 = 7'h64 == out_payload_rob_idx[6:0] ? rob_payload_100_rob_idx : _GEN_8420; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8422 = 7'h65 == out_payload_rob_idx[6:0] ? rob_payload_101_rob_idx : _GEN_8421; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8423 = 7'h66 == out_payload_rob_idx[6:0] ? rob_payload_102_rob_idx : _GEN_8422; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8424 = 7'h67 == out_payload_rob_idx[6:0] ? rob_payload_103_rob_idx : _GEN_8423; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8425 = 7'h68 == out_payload_rob_idx[6:0] ? rob_payload_104_rob_idx : _GEN_8424; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8426 = 7'h69 == out_payload_rob_idx[6:0] ? rob_payload_105_rob_idx : _GEN_8425; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8427 = 7'h6a == out_payload_rob_idx[6:0] ? rob_payload_106_rob_idx : _GEN_8426; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8428 = 7'h6b == out_payload_rob_idx[6:0] ? rob_payload_107_rob_idx : _GEN_8427; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8429 = 7'h6c == out_payload_rob_idx[6:0] ? rob_payload_108_rob_idx : _GEN_8428; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8430 = 7'h6d == out_payload_rob_idx[6:0] ? rob_payload_109_rob_idx : _GEN_8429; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8431 = 7'h6e == out_payload_rob_idx[6:0] ? rob_payload_110_rob_idx : _GEN_8430; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8432 = 7'h6f == out_payload_rob_idx[6:0] ? rob_payload_111_rob_idx : _GEN_8431; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8433 = 7'h70 == out_payload_rob_idx[6:0] ? rob_payload_112_rob_idx : _GEN_8432; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8434 = 7'h71 == out_payload_rob_idx[6:0] ? rob_payload_113_rob_idx : _GEN_8433; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8435 = 7'h72 == out_payload_rob_idx[6:0] ? rob_payload_114_rob_idx : _GEN_8434; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8436 = 7'h73 == out_payload_rob_idx[6:0] ? rob_payload_115_rob_idx : _GEN_8435; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8437 = 7'h74 == out_payload_rob_idx[6:0] ? rob_payload_116_rob_idx : _GEN_8436; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8438 = 7'h75 == out_payload_rob_idx[6:0] ? rob_payload_117_rob_idx : _GEN_8437; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8439 = 7'h76 == out_payload_rob_idx[6:0] ? rob_payload_118_rob_idx : _GEN_8438; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8440 = 7'h77 == out_payload_rob_idx[6:0] ? rob_payload_119_rob_idx : _GEN_8439; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8441 = 7'h78 == out_payload_rob_idx[6:0] ? rob_payload_120_rob_idx : _GEN_8440; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8442 = 7'h79 == out_payload_rob_idx[6:0] ? rob_payload_121_rob_idx : _GEN_8441; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8443 = 7'h7a == out_payload_rob_idx[6:0] ? rob_payload_122_rob_idx : _GEN_8442; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8444 = 7'h7b == out_payload_rob_idx[6:0] ? rob_payload_123_rob_idx : _GEN_8443; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8445 = 7'h7c == out_payload_rob_idx[6:0] ? rob_payload_124_rob_idx : _GEN_8444; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8446 = 7'h7d == out_payload_rob_idx[6:0] ? rob_payload_125_rob_idx : _GEN_8445; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8447 = 7'h7e == out_payload_rob_idx[6:0] ? rob_payload_126_rob_idx : _GEN_8446; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8448 = 7'h7f == out_payload_rob_idx[6:0] ? rob_payload_127_rob_idx : _GEN_8447; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8450 = 7'h1 == out_payload_rob_idx[6:0] ? rob_payload_1_flits_fired : rob_payload_0_flits_fired; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8451 = 7'h2 == out_payload_rob_idx[6:0] ? rob_payload_2_flits_fired : _GEN_8450; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8452 = 7'h3 == out_payload_rob_idx[6:0] ? rob_payload_3_flits_fired : _GEN_8451; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8453 = 7'h4 == out_payload_rob_idx[6:0] ? rob_payload_4_flits_fired : _GEN_8452; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8454 = 7'h5 == out_payload_rob_idx[6:0] ? rob_payload_5_flits_fired : _GEN_8453; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8455 = 7'h6 == out_payload_rob_idx[6:0] ? rob_payload_6_flits_fired : _GEN_8454; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8456 = 7'h7 == out_payload_rob_idx[6:0] ? rob_payload_7_flits_fired : _GEN_8455; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8457 = 7'h8 == out_payload_rob_idx[6:0] ? rob_payload_8_flits_fired : _GEN_8456; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8458 = 7'h9 == out_payload_rob_idx[6:0] ? rob_payload_9_flits_fired : _GEN_8457; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8459 = 7'ha == out_payload_rob_idx[6:0] ? rob_payload_10_flits_fired : _GEN_8458; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8460 = 7'hb == out_payload_rob_idx[6:0] ? rob_payload_11_flits_fired : _GEN_8459; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8461 = 7'hc == out_payload_rob_idx[6:0] ? rob_payload_12_flits_fired : _GEN_8460; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8462 = 7'hd == out_payload_rob_idx[6:0] ? rob_payload_13_flits_fired : _GEN_8461; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8463 = 7'he == out_payload_rob_idx[6:0] ? rob_payload_14_flits_fired : _GEN_8462; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8464 = 7'hf == out_payload_rob_idx[6:0] ? rob_payload_15_flits_fired : _GEN_8463; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8465 = 7'h10 == out_payload_rob_idx[6:0] ? rob_payload_16_flits_fired : _GEN_8464; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8466 = 7'h11 == out_payload_rob_idx[6:0] ? rob_payload_17_flits_fired : _GEN_8465; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8467 = 7'h12 == out_payload_rob_idx[6:0] ? rob_payload_18_flits_fired : _GEN_8466; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8468 = 7'h13 == out_payload_rob_idx[6:0] ? rob_payload_19_flits_fired : _GEN_8467; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8469 = 7'h14 == out_payload_rob_idx[6:0] ? rob_payload_20_flits_fired : _GEN_8468; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8470 = 7'h15 == out_payload_rob_idx[6:0] ? rob_payload_21_flits_fired : _GEN_8469; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8471 = 7'h16 == out_payload_rob_idx[6:0] ? rob_payload_22_flits_fired : _GEN_8470; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8472 = 7'h17 == out_payload_rob_idx[6:0] ? rob_payload_23_flits_fired : _GEN_8471; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8473 = 7'h18 == out_payload_rob_idx[6:0] ? rob_payload_24_flits_fired : _GEN_8472; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8474 = 7'h19 == out_payload_rob_idx[6:0] ? rob_payload_25_flits_fired : _GEN_8473; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8475 = 7'h1a == out_payload_rob_idx[6:0] ? rob_payload_26_flits_fired : _GEN_8474; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8476 = 7'h1b == out_payload_rob_idx[6:0] ? rob_payload_27_flits_fired : _GEN_8475; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8477 = 7'h1c == out_payload_rob_idx[6:0] ? rob_payload_28_flits_fired : _GEN_8476; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8478 = 7'h1d == out_payload_rob_idx[6:0] ? rob_payload_29_flits_fired : _GEN_8477; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8479 = 7'h1e == out_payload_rob_idx[6:0] ? rob_payload_30_flits_fired : _GEN_8478; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8480 = 7'h1f == out_payload_rob_idx[6:0] ? rob_payload_31_flits_fired : _GEN_8479; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8481 = 7'h20 == out_payload_rob_idx[6:0] ? rob_payload_32_flits_fired : _GEN_8480; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8482 = 7'h21 == out_payload_rob_idx[6:0] ? rob_payload_33_flits_fired : _GEN_8481; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8483 = 7'h22 == out_payload_rob_idx[6:0] ? rob_payload_34_flits_fired : _GEN_8482; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8484 = 7'h23 == out_payload_rob_idx[6:0] ? rob_payload_35_flits_fired : _GEN_8483; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8485 = 7'h24 == out_payload_rob_idx[6:0] ? rob_payload_36_flits_fired : _GEN_8484; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8486 = 7'h25 == out_payload_rob_idx[6:0] ? rob_payload_37_flits_fired : _GEN_8485; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8487 = 7'h26 == out_payload_rob_idx[6:0] ? rob_payload_38_flits_fired : _GEN_8486; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8488 = 7'h27 == out_payload_rob_idx[6:0] ? rob_payload_39_flits_fired : _GEN_8487; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8489 = 7'h28 == out_payload_rob_idx[6:0] ? rob_payload_40_flits_fired : _GEN_8488; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8490 = 7'h29 == out_payload_rob_idx[6:0] ? rob_payload_41_flits_fired : _GEN_8489; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8491 = 7'h2a == out_payload_rob_idx[6:0] ? rob_payload_42_flits_fired : _GEN_8490; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8492 = 7'h2b == out_payload_rob_idx[6:0] ? rob_payload_43_flits_fired : _GEN_8491; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8493 = 7'h2c == out_payload_rob_idx[6:0] ? rob_payload_44_flits_fired : _GEN_8492; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8494 = 7'h2d == out_payload_rob_idx[6:0] ? rob_payload_45_flits_fired : _GEN_8493; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8495 = 7'h2e == out_payload_rob_idx[6:0] ? rob_payload_46_flits_fired : _GEN_8494; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8496 = 7'h2f == out_payload_rob_idx[6:0] ? rob_payload_47_flits_fired : _GEN_8495; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8497 = 7'h30 == out_payload_rob_idx[6:0] ? rob_payload_48_flits_fired : _GEN_8496; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8498 = 7'h31 == out_payload_rob_idx[6:0] ? rob_payload_49_flits_fired : _GEN_8497; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8499 = 7'h32 == out_payload_rob_idx[6:0] ? rob_payload_50_flits_fired : _GEN_8498; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8500 = 7'h33 == out_payload_rob_idx[6:0] ? rob_payload_51_flits_fired : _GEN_8499; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8501 = 7'h34 == out_payload_rob_idx[6:0] ? rob_payload_52_flits_fired : _GEN_8500; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8502 = 7'h35 == out_payload_rob_idx[6:0] ? rob_payload_53_flits_fired : _GEN_8501; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8503 = 7'h36 == out_payload_rob_idx[6:0] ? rob_payload_54_flits_fired : _GEN_8502; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8504 = 7'h37 == out_payload_rob_idx[6:0] ? rob_payload_55_flits_fired : _GEN_8503; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8505 = 7'h38 == out_payload_rob_idx[6:0] ? rob_payload_56_flits_fired : _GEN_8504; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8506 = 7'h39 == out_payload_rob_idx[6:0] ? rob_payload_57_flits_fired : _GEN_8505; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8507 = 7'h3a == out_payload_rob_idx[6:0] ? rob_payload_58_flits_fired : _GEN_8506; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8508 = 7'h3b == out_payload_rob_idx[6:0] ? rob_payload_59_flits_fired : _GEN_8507; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8509 = 7'h3c == out_payload_rob_idx[6:0] ? rob_payload_60_flits_fired : _GEN_8508; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8510 = 7'h3d == out_payload_rob_idx[6:0] ? rob_payload_61_flits_fired : _GEN_8509; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8511 = 7'h3e == out_payload_rob_idx[6:0] ? rob_payload_62_flits_fired : _GEN_8510; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8512 = 7'h3f == out_payload_rob_idx[6:0] ? rob_payload_63_flits_fired : _GEN_8511; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8513 = 7'h40 == out_payload_rob_idx[6:0] ? rob_payload_64_flits_fired : _GEN_8512; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8514 = 7'h41 == out_payload_rob_idx[6:0] ? rob_payload_65_flits_fired : _GEN_8513; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8515 = 7'h42 == out_payload_rob_idx[6:0] ? rob_payload_66_flits_fired : _GEN_8514; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8516 = 7'h43 == out_payload_rob_idx[6:0] ? rob_payload_67_flits_fired : _GEN_8515; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8517 = 7'h44 == out_payload_rob_idx[6:0] ? rob_payload_68_flits_fired : _GEN_8516; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8518 = 7'h45 == out_payload_rob_idx[6:0] ? rob_payload_69_flits_fired : _GEN_8517; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8519 = 7'h46 == out_payload_rob_idx[6:0] ? rob_payload_70_flits_fired : _GEN_8518; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8520 = 7'h47 == out_payload_rob_idx[6:0] ? rob_payload_71_flits_fired : _GEN_8519; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8521 = 7'h48 == out_payload_rob_idx[6:0] ? rob_payload_72_flits_fired : _GEN_8520; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8522 = 7'h49 == out_payload_rob_idx[6:0] ? rob_payload_73_flits_fired : _GEN_8521; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8523 = 7'h4a == out_payload_rob_idx[6:0] ? rob_payload_74_flits_fired : _GEN_8522; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8524 = 7'h4b == out_payload_rob_idx[6:0] ? rob_payload_75_flits_fired : _GEN_8523; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8525 = 7'h4c == out_payload_rob_idx[6:0] ? rob_payload_76_flits_fired : _GEN_8524; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8526 = 7'h4d == out_payload_rob_idx[6:0] ? rob_payload_77_flits_fired : _GEN_8525; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8527 = 7'h4e == out_payload_rob_idx[6:0] ? rob_payload_78_flits_fired : _GEN_8526; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8528 = 7'h4f == out_payload_rob_idx[6:0] ? rob_payload_79_flits_fired : _GEN_8527; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8529 = 7'h50 == out_payload_rob_idx[6:0] ? rob_payload_80_flits_fired : _GEN_8528; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8530 = 7'h51 == out_payload_rob_idx[6:0] ? rob_payload_81_flits_fired : _GEN_8529; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8531 = 7'h52 == out_payload_rob_idx[6:0] ? rob_payload_82_flits_fired : _GEN_8530; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8532 = 7'h53 == out_payload_rob_idx[6:0] ? rob_payload_83_flits_fired : _GEN_8531; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8533 = 7'h54 == out_payload_rob_idx[6:0] ? rob_payload_84_flits_fired : _GEN_8532; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8534 = 7'h55 == out_payload_rob_idx[6:0] ? rob_payload_85_flits_fired : _GEN_8533; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8535 = 7'h56 == out_payload_rob_idx[6:0] ? rob_payload_86_flits_fired : _GEN_8534; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8536 = 7'h57 == out_payload_rob_idx[6:0] ? rob_payload_87_flits_fired : _GEN_8535; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8537 = 7'h58 == out_payload_rob_idx[6:0] ? rob_payload_88_flits_fired : _GEN_8536; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8538 = 7'h59 == out_payload_rob_idx[6:0] ? rob_payload_89_flits_fired : _GEN_8537; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8539 = 7'h5a == out_payload_rob_idx[6:0] ? rob_payload_90_flits_fired : _GEN_8538; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8540 = 7'h5b == out_payload_rob_idx[6:0] ? rob_payload_91_flits_fired : _GEN_8539; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8541 = 7'h5c == out_payload_rob_idx[6:0] ? rob_payload_92_flits_fired : _GEN_8540; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8542 = 7'h5d == out_payload_rob_idx[6:0] ? rob_payload_93_flits_fired : _GEN_8541; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8543 = 7'h5e == out_payload_rob_idx[6:0] ? rob_payload_94_flits_fired : _GEN_8542; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8544 = 7'h5f == out_payload_rob_idx[6:0] ? rob_payload_95_flits_fired : _GEN_8543; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8545 = 7'h60 == out_payload_rob_idx[6:0] ? rob_payload_96_flits_fired : _GEN_8544; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8546 = 7'h61 == out_payload_rob_idx[6:0] ? rob_payload_97_flits_fired : _GEN_8545; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8547 = 7'h62 == out_payload_rob_idx[6:0] ? rob_payload_98_flits_fired : _GEN_8546; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8548 = 7'h63 == out_payload_rob_idx[6:0] ? rob_payload_99_flits_fired : _GEN_8547; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8549 = 7'h64 == out_payload_rob_idx[6:0] ? rob_payload_100_flits_fired : _GEN_8548; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8550 = 7'h65 == out_payload_rob_idx[6:0] ? rob_payload_101_flits_fired : _GEN_8549; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8551 = 7'h66 == out_payload_rob_idx[6:0] ? rob_payload_102_flits_fired : _GEN_8550; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8552 = 7'h67 == out_payload_rob_idx[6:0] ? rob_payload_103_flits_fired : _GEN_8551; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8553 = 7'h68 == out_payload_rob_idx[6:0] ? rob_payload_104_flits_fired : _GEN_8552; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8554 = 7'h69 == out_payload_rob_idx[6:0] ? rob_payload_105_flits_fired : _GEN_8553; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8555 = 7'h6a == out_payload_rob_idx[6:0] ? rob_payload_106_flits_fired : _GEN_8554; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8556 = 7'h6b == out_payload_rob_idx[6:0] ? rob_payload_107_flits_fired : _GEN_8555; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8557 = 7'h6c == out_payload_rob_idx[6:0] ? rob_payload_108_flits_fired : _GEN_8556; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8558 = 7'h6d == out_payload_rob_idx[6:0] ? rob_payload_109_flits_fired : _GEN_8557; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8559 = 7'h6e == out_payload_rob_idx[6:0] ? rob_payload_110_flits_fired : _GEN_8558; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8560 = 7'h6f == out_payload_rob_idx[6:0] ? rob_payload_111_flits_fired : _GEN_8559; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8561 = 7'h70 == out_payload_rob_idx[6:0] ? rob_payload_112_flits_fired : _GEN_8560; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8562 = 7'h71 == out_payload_rob_idx[6:0] ? rob_payload_113_flits_fired : _GEN_8561; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8563 = 7'h72 == out_payload_rob_idx[6:0] ? rob_payload_114_flits_fired : _GEN_8562; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8564 = 7'h73 == out_payload_rob_idx[6:0] ? rob_payload_115_flits_fired : _GEN_8563; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8565 = 7'h74 == out_payload_rob_idx[6:0] ? rob_payload_116_flits_fired : _GEN_8564; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8566 = 7'h75 == out_payload_rob_idx[6:0] ? rob_payload_117_flits_fired : _GEN_8565; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8567 = 7'h76 == out_payload_rob_idx[6:0] ? rob_payload_118_flits_fired : _GEN_8566; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8568 = 7'h77 == out_payload_rob_idx[6:0] ? rob_payload_119_flits_fired : _GEN_8567; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8569 = 7'h78 == out_payload_rob_idx[6:0] ? rob_payload_120_flits_fired : _GEN_8568; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8570 = 7'h79 == out_payload_rob_idx[6:0] ? rob_payload_121_flits_fired : _GEN_8569; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8571 = 7'h7a == out_payload_rob_idx[6:0] ? rob_payload_122_flits_fired : _GEN_8570; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8572 = 7'h7b == out_payload_rob_idx[6:0] ? rob_payload_123_flits_fired : _GEN_8571; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8573 = 7'h7c == out_payload_rob_idx[6:0] ? rob_payload_124_flits_fired : _GEN_8572; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8574 = 7'h7d == out_payload_rob_idx[6:0] ? rob_payload_125_flits_fired : _GEN_8573; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8575 = 7'h7e == out_payload_rob_idx[6:0] ? rob_payload_126_flits_fired : _GEN_8574; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_8576 = 7'h7f == out_payload_rob_idx[6:0] ? rob_payload_127_flits_fired : _GEN_8575; // @[TestHarness.scala 202:{35,35}]
  wire [63:0] _T_82 = {_GEN_8320,_GEN_8448,_GEN_8576}; // @[TestHarness.scala 202:35]
  wire [1:0] _GEN_8578 = 7'h1 == out_payload_rob_idx[6:0] ? rob_ingress_id_1 : rob_ingress_id_0; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8579 = 7'h2 == out_payload_rob_idx[6:0] ? rob_ingress_id_2 : _GEN_8578; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8580 = 7'h3 == out_payload_rob_idx[6:0] ? rob_ingress_id_3 : _GEN_8579; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8581 = 7'h4 == out_payload_rob_idx[6:0] ? rob_ingress_id_4 : _GEN_8580; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8582 = 7'h5 == out_payload_rob_idx[6:0] ? rob_ingress_id_5 : _GEN_8581; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8583 = 7'h6 == out_payload_rob_idx[6:0] ? rob_ingress_id_6 : _GEN_8582; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8584 = 7'h7 == out_payload_rob_idx[6:0] ? rob_ingress_id_7 : _GEN_8583; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8585 = 7'h8 == out_payload_rob_idx[6:0] ? rob_ingress_id_8 : _GEN_8584; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8586 = 7'h9 == out_payload_rob_idx[6:0] ? rob_ingress_id_9 : _GEN_8585; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8587 = 7'ha == out_payload_rob_idx[6:0] ? rob_ingress_id_10 : _GEN_8586; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8588 = 7'hb == out_payload_rob_idx[6:0] ? rob_ingress_id_11 : _GEN_8587; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8589 = 7'hc == out_payload_rob_idx[6:0] ? rob_ingress_id_12 : _GEN_8588; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8590 = 7'hd == out_payload_rob_idx[6:0] ? rob_ingress_id_13 : _GEN_8589; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8591 = 7'he == out_payload_rob_idx[6:0] ? rob_ingress_id_14 : _GEN_8590; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8592 = 7'hf == out_payload_rob_idx[6:0] ? rob_ingress_id_15 : _GEN_8591; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8593 = 7'h10 == out_payload_rob_idx[6:0] ? rob_ingress_id_16 : _GEN_8592; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8594 = 7'h11 == out_payload_rob_idx[6:0] ? rob_ingress_id_17 : _GEN_8593; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8595 = 7'h12 == out_payload_rob_idx[6:0] ? rob_ingress_id_18 : _GEN_8594; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8596 = 7'h13 == out_payload_rob_idx[6:0] ? rob_ingress_id_19 : _GEN_8595; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8597 = 7'h14 == out_payload_rob_idx[6:0] ? rob_ingress_id_20 : _GEN_8596; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8598 = 7'h15 == out_payload_rob_idx[6:0] ? rob_ingress_id_21 : _GEN_8597; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8599 = 7'h16 == out_payload_rob_idx[6:0] ? rob_ingress_id_22 : _GEN_8598; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8600 = 7'h17 == out_payload_rob_idx[6:0] ? rob_ingress_id_23 : _GEN_8599; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8601 = 7'h18 == out_payload_rob_idx[6:0] ? rob_ingress_id_24 : _GEN_8600; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8602 = 7'h19 == out_payload_rob_idx[6:0] ? rob_ingress_id_25 : _GEN_8601; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8603 = 7'h1a == out_payload_rob_idx[6:0] ? rob_ingress_id_26 : _GEN_8602; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8604 = 7'h1b == out_payload_rob_idx[6:0] ? rob_ingress_id_27 : _GEN_8603; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8605 = 7'h1c == out_payload_rob_idx[6:0] ? rob_ingress_id_28 : _GEN_8604; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8606 = 7'h1d == out_payload_rob_idx[6:0] ? rob_ingress_id_29 : _GEN_8605; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8607 = 7'h1e == out_payload_rob_idx[6:0] ? rob_ingress_id_30 : _GEN_8606; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8608 = 7'h1f == out_payload_rob_idx[6:0] ? rob_ingress_id_31 : _GEN_8607; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8609 = 7'h20 == out_payload_rob_idx[6:0] ? rob_ingress_id_32 : _GEN_8608; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8610 = 7'h21 == out_payload_rob_idx[6:0] ? rob_ingress_id_33 : _GEN_8609; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8611 = 7'h22 == out_payload_rob_idx[6:0] ? rob_ingress_id_34 : _GEN_8610; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8612 = 7'h23 == out_payload_rob_idx[6:0] ? rob_ingress_id_35 : _GEN_8611; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8613 = 7'h24 == out_payload_rob_idx[6:0] ? rob_ingress_id_36 : _GEN_8612; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8614 = 7'h25 == out_payload_rob_idx[6:0] ? rob_ingress_id_37 : _GEN_8613; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8615 = 7'h26 == out_payload_rob_idx[6:0] ? rob_ingress_id_38 : _GEN_8614; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8616 = 7'h27 == out_payload_rob_idx[6:0] ? rob_ingress_id_39 : _GEN_8615; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8617 = 7'h28 == out_payload_rob_idx[6:0] ? rob_ingress_id_40 : _GEN_8616; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8618 = 7'h29 == out_payload_rob_idx[6:0] ? rob_ingress_id_41 : _GEN_8617; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8619 = 7'h2a == out_payload_rob_idx[6:0] ? rob_ingress_id_42 : _GEN_8618; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8620 = 7'h2b == out_payload_rob_idx[6:0] ? rob_ingress_id_43 : _GEN_8619; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8621 = 7'h2c == out_payload_rob_idx[6:0] ? rob_ingress_id_44 : _GEN_8620; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8622 = 7'h2d == out_payload_rob_idx[6:0] ? rob_ingress_id_45 : _GEN_8621; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8623 = 7'h2e == out_payload_rob_idx[6:0] ? rob_ingress_id_46 : _GEN_8622; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8624 = 7'h2f == out_payload_rob_idx[6:0] ? rob_ingress_id_47 : _GEN_8623; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8625 = 7'h30 == out_payload_rob_idx[6:0] ? rob_ingress_id_48 : _GEN_8624; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8626 = 7'h31 == out_payload_rob_idx[6:0] ? rob_ingress_id_49 : _GEN_8625; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8627 = 7'h32 == out_payload_rob_idx[6:0] ? rob_ingress_id_50 : _GEN_8626; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8628 = 7'h33 == out_payload_rob_idx[6:0] ? rob_ingress_id_51 : _GEN_8627; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8629 = 7'h34 == out_payload_rob_idx[6:0] ? rob_ingress_id_52 : _GEN_8628; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8630 = 7'h35 == out_payload_rob_idx[6:0] ? rob_ingress_id_53 : _GEN_8629; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8631 = 7'h36 == out_payload_rob_idx[6:0] ? rob_ingress_id_54 : _GEN_8630; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8632 = 7'h37 == out_payload_rob_idx[6:0] ? rob_ingress_id_55 : _GEN_8631; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8633 = 7'h38 == out_payload_rob_idx[6:0] ? rob_ingress_id_56 : _GEN_8632; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8634 = 7'h39 == out_payload_rob_idx[6:0] ? rob_ingress_id_57 : _GEN_8633; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8635 = 7'h3a == out_payload_rob_idx[6:0] ? rob_ingress_id_58 : _GEN_8634; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8636 = 7'h3b == out_payload_rob_idx[6:0] ? rob_ingress_id_59 : _GEN_8635; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8637 = 7'h3c == out_payload_rob_idx[6:0] ? rob_ingress_id_60 : _GEN_8636; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8638 = 7'h3d == out_payload_rob_idx[6:0] ? rob_ingress_id_61 : _GEN_8637; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8639 = 7'h3e == out_payload_rob_idx[6:0] ? rob_ingress_id_62 : _GEN_8638; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8640 = 7'h3f == out_payload_rob_idx[6:0] ? rob_ingress_id_63 : _GEN_8639; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8641 = 7'h40 == out_payload_rob_idx[6:0] ? rob_ingress_id_64 : _GEN_8640; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8642 = 7'h41 == out_payload_rob_idx[6:0] ? rob_ingress_id_65 : _GEN_8641; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8643 = 7'h42 == out_payload_rob_idx[6:0] ? rob_ingress_id_66 : _GEN_8642; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8644 = 7'h43 == out_payload_rob_idx[6:0] ? rob_ingress_id_67 : _GEN_8643; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8645 = 7'h44 == out_payload_rob_idx[6:0] ? rob_ingress_id_68 : _GEN_8644; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8646 = 7'h45 == out_payload_rob_idx[6:0] ? rob_ingress_id_69 : _GEN_8645; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8647 = 7'h46 == out_payload_rob_idx[6:0] ? rob_ingress_id_70 : _GEN_8646; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8648 = 7'h47 == out_payload_rob_idx[6:0] ? rob_ingress_id_71 : _GEN_8647; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8649 = 7'h48 == out_payload_rob_idx[6:0] ? rob_ingress_id_72 : _GEN_8648; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8650 = 7'h49 == out_payload_rob_idx[6:0] ? rob_ingress_id_73 : _GEN_8649; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8651 = 7'h4a == out_payload_rob_idx[6:0] ? rob_ingress_id_74 : _GEN_8650; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8652 = 7'h4b == out_payload_rob_idx[6:0] ? rob_ingress_id_75 : _GEN_8651; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8653 = 7'h4c == out_payload_rob_idx[6:0] ? rob_ingress_id_76 : _GEN_8652; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8654 = 7'h4d == out_payload_rob_idx[6:0] ? rob_ingress_id_77 : _GEN_8653; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8655 = 7'h4e == out_payload_rob_idx[6:0] ? rob_ingress_id_78 : _GEN_8654; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8656 = 7'h4f == out_payload_rob_idx[6:0] ? rob_ingress_id_79 : _GEN_8655; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8657 = 7'h50 == out_payload_rob_idx[6:0] ? rob_ingress_id_80 : _GEN_8656; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8658 = 7'h51 == out_payload_rob_idx[6:0] ? rob_ingress_id_81 : _GEN_8657; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8659 = 7'h52 == out_payload_rob_idx[6:0] ? rob_ingress_id_82 : _GEN_8658; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8660 = 7'h53 == out_payload_rob_idx[6:0] ? rob_ingress_id_83 : _GEN_8659; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8661 = 7'h54 == out_payload_rob_idx[6:0] ? rob_ingress_id_84 : _GEN_8660; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8662 = 7'h55 == out_payload_rob_idx[6:0] ? rob_ingress_id_85 : _GEN_8661; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8663 = 7'h56 == out_payload_rob_idx[6:0] ? rob_ingress_id_86 : _GEN_8662; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8664 = 7'h57 == out_payload_rob_idx[6:0] ? rob_ingress_id_87 : _GEN_8663; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8665 = 7'h58 == out_payload_rob_idx[6:0] ? rob_ingress_id_88 : _GEN_8664; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8666 = 7'h59 == out_payload_rob_idx[6:0] ? rob_ingress_id_89 : _GEN_8665; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8667 = 7'h5a == out_payload_rob_idx[6:0] ? rob_ingress_id_90 : _GEN_8666; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8668 = 7'h5b == out_payload_rob_idx[6:0] ? rob_ingress_id_91 : _GEN_8667; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8669 = 7'h5c == out_payload_rob_idx[6:0] ? rob_ingress_id_92 : _GEN_8668; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8670 = 7'h5d == out_payload_rob_idx[6:0] ? rob_ingress_id_93 : _GEN_8669; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8671 = 7'h5e == out_payload_rob_idx[6:0] ? rob_ingress_id_94 : _GEN_8670; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8672 = 7'h5f == out_payload_rob_idx[6:0] ? rob_ingress_id_95 : _GEN_8671; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8673 = 7'h60 == out_payload_rob_idx[6:0] ? rob_ingress_id_96 : _GEN_8672; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8674 = 7'h61 == out_payload_rob_idx[6:0] ? rob_ingress_id_97 : _GEN_8673; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8675 = 7'h62 == out_payload_rob_idx[6:0] ? rob_ingress_id_98 : _GEN_8674; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8676 = 7'h63 == out_payload_rob_idx[6:0] ? rob_ingress_id_99 : _GEN_8675; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8677 = 7'h64 == out_payload_rob_idx[6:0] ? rob_ingress_id_100 : _GEN_8676; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8678 = 7'h65 == out_payload_rob_idx[6:0] ? rob_ingress_id_101 : _GEN_8677; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8679 = 7'h66 == out_payload_rob_idx[6:0] ? rob_ingress_id_102 : _GEN_8678; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8680 = 7'h67 == out_payload_rob_idx[6:0] ? rob_ingress_id_103 : _GEN_8679; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8681 = 7'h68 == out_payload_rob_idx[6:0] ? rob_ingress_id_104 : _GEN_8680; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8682 = 7'h69 == out_payload_rob_idx[6:0] ? rob_ingress_id_105 : _GEN_8681; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8683 = 7'h6a == out_payload_rob_idx[6:0] ? rob_ingress_id_106 : _GEN_8682; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8684 = 7'h6b == out_payload_rob_idx[6:0] ? rob_ingress_id_107 : _GEN_8683; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8685 = 7'h6c == out_payload_rob_idx[6:0] ? rob_ingress_id_108 : _GEN_8684; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8686 = 7'h6d == out_payload_rob_idx[6:0] ? rob_ingress_id_109 : _GEN_8685; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8687 = 7'h6e == out_payload_rob_idx[6:0] ? rob_ingress_id_110 : _GEN_8686; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8688 = 7'h6f == out_payload_rob_idx[6:0] ? rob_ingress_id_111 : _GEN_8687; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8689 = 7'h70 == out_payload_rob_idx[6:0] ? rob_ingress_id_112 : _GEN_8688; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8690 = 7'h71 == out_payload_rob_idx[6:0] ? rob_ingress_id_113 : _GEN_8689; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8691 = 7'h72 == out_payload_rob_idx[6:0] ? rob_ingress_id_114 : _GEN_8690; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8692 = 7'h73 == out_payload_rob_idx[6:0] ? rob_ingress_id_115 : _GEN_8691; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8693 = 7'h74 == out_payload_rob_idx[6:0] ? rob_ingress_id_116 : _GEN_8692; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8694 = 7'h75 == out_payload_rob_idx[6:0] ? rob_ingress_id_117 : _GEN_8693; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8695 = 7'h76 == out_payload_rob_idx[6:0] ? rob_ingress_id_118 : _GEN_8694; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8696 = 7'h77 == out_payload_rob_idx[6:0] ? rob_ingress_id_119 : _GEN_8695; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8697 = 7'h78 == out_payload_rob_idx[6:0] ? rob_ingress_id_120 : _GEN_8696; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8698 = 7'h79 == out_payload_rob_idx[6:0] ? rob_ingress_id_121 : _GEN_8697; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8699 = 7'h7a == out_payload_rob_idx[6:0] ? rob_ingress_id_122 : _GEN_8698; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8700 = 7'h7b == out_payload_rob_idx[6:0] ? rob_ingress_id_123 : _GEN_8699; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8701 = 7'h7c == out_payload_rob_idx[6:0] ? rob_ingress_id_124 : _GEN_8700; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8702 = 7'h7d == out_payload_rob_idx[6:0] ? rob_ingress_id_125 : _GEN_8701; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8703 = 7'h7e == out_payload_rob_idx[6:0] ? rob_ingress_id_126 : _GEN_8702; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8704 = 7'h7f == out_payload_rob_idx[6:0] ? rob_ingress_id_127 : _GEN_8703; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_8706 = 7'h1 == out_payload_rob_idx[6:0] ? rob_egress_id_1 : rob_egress_id_0; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8707 = 7'h2 == out_payload_rob_idx[6:0] ? rob_egress_id_2 : _GEN_8706; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8708 = 7'h3 == out_payload_rob_idx[6:0] ? rob_egress_id_3 : _GEN_8707; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8709 = 7'h4 == out_payload_rob_idx[6:0] ? rob_egress_id_4 : _GEN_8708; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8710 = 7'h5 == out_payload_rob_idx[6:0] ? rob_egress_id_5 : _GEN_8709; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8711 = 7'h6 == out_payload_rob_idx[6:0] ? rob_egress_id_6 : _GEN_8710; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8712 = 7'h7 == out_payload_rob_idx[6:0] ? rob_egress_id_7 : _GEN_8711; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8713 = 7'h8 == out_payload_rob_idx[6:0] ? rob_egress_id_8 : _GEN_8712; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8714 = 7'h9 == out_payload_rob_idx[6:0] ? rob_egress_id_9 : _GEN_8713; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8715 = 7'ha == out_payload_rob_idx[6:0] ? rob_egress_id_10 : _GEN_8714; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8716 = 7'hb == out_payload_rob_idx[6:0] ? rob_egress_id_11 : _GEN_8715; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8717 = 7'hc == out_payload_rob_idx[6:0] ? rob_egress_id_12 : _GEN_8716; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8718 = 7'hd == out_payload_rob_idx[6:0] ? rob_egress_id_13 : _GEN_8717; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8719 = 7'he == out_payload_rob_idx[6:0] ? rob_egress_id_14 : _GEN_8718; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8720 = 7'hf == out_payload_rob_idx[6:0] ? rob_egress_id_15 : _GEN_8719; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8721 = 7'h10 == out_payload_rob_idx[6:0] ? rob_egress_id_16 : _GEN_8720; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8722 = 7'h11 == out_payload_rob_idx[6:0] ? rob_egress_id_17 : _GEN_8721; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8723 = 7'h12 == out_payload_rob_idx[6:0] ? rob_egress_id_18 : _GEN_8722; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8724 = 7'h13 == out_payload_rob_idx[6:0] ? rob_egress_id_19 : _GEN_8723; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8725 = 7'h14 == out_payload_rob_idx[6:0] ? rob_egress_id_20 : _GEN_8724; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8726 = 7'h15 == out_payload_rob_idx[6:0] ? rob_egress_id_21 : _GEN_8725; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8727 = 7'h16 == out_payload_rob_idx[6:0] ? rob_egress_id_22 : _GEN_8726; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8728 = 7'h17 == out_payload_rob_idx[6:0] ? rob_egress_id_23 : _GEN_8727; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8729 = 7'h18 == out_payload_rob_idx[6:0] ? rob_egress_id_24 : _GEN_8728; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8730 = 7'h19 == out_payload_rob_idx[6:0] ? rob_egress_id_25 : _GEN_8729; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8731 = 7'h1a == out_payload_rob_idx[6:0] ? rob_egress_id_26 : _GEN_8730; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8732 = 7'h1b == out_payload_rob_idx[6:0] ? rob_egress_id_27 : _GEN_8731; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8733 = 7'h1c == out_payload_rob_idx[6:0] ? rob_egress_id_28 : _GEN_8732; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8734 = 7'h1d == out_payload_rob_idx[6:0] ? rob_egress_id_29 : _GEN_8733; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8735 = 7'h1e == out_payload_rob_idx[6:0] ? rob_egress_id_30 : _GEN_8734; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8736 = 7'h1f == out_payload_rob_idx[6:0] ? rob_egress_id_31 : _GEN_8735; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8737 = 7'h20 == out_payload_rob_idx[6:0] ? rob_egress_id_32 : _GEN_8736; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8738 = 7'h21 == out_payload_rob_idx[6:0] ? rob_egress_id_33 : _GEN_8737; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8739 = 7'h22 == out_payload_rob_idx[6:0] ? rob_egress_id_34 : _GEN_8738; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8740 = 7'h23 == out_payload_rob_idx[6:0] ? rob_egress_id_35 : _GEN_8739; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8741 = 7'h24 == out_payload_rob_idx[6:0] ? rob_egress_id_36 : _GEN_8740; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8742 = 7'h25 == out_payload_rob_idx[6:0] ? rob_egress_id_37 : _GEN_8741; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8743 = 7'h26 == out_payload_rob_idx[6:0] ? rob_egress_id_38 : _GEN_8742; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8744 = 7'h27 == out_payload_rob_idx[6:0] ? rob_egress_id_39 : _GEN_8743; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8745 = 7'h28 == out_payload_rob_idx[6:0] ? rob_egress_id_40 : _GEN_8744; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8746 = 7'h29 == out_payload_rob_idx[6:0] ? rob_egress_id_41 : _GEN_8745; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8747 = 7'h2a == out_payload_rob_idx[6:0] ? rob_egress_id_42 : _GEN_8746; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8748 = 7'h2b == out_payload_rob_idx[6:0] ? rob_egress_id_43 : _GEN_8747; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8749 = 7'h2c == out_payload_rob_idx[6:0] ? rob_egress_id_44 : _GEN_8748; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8750 = 7'h2d == out_payload_rob_idx[6:0] ? rob_egress_id_45 : _GEN_8749; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8751 = 7'h2e == out_payload_rob_idx[6:0] ? rob_egress_id_46 : _GEN_8750; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8752 = 7'h2f == out_payload_rob_idx[6:0] ? rob_egress_id_47 : _GEN_8751; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8753 = 7'h30 == out_payload_rob_idx[6:0] ? rob_egress_id_48 : _GEN_8752; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8754 = 7'h31 == out_payload_rob_idx[6:0] ? rob_egress_id_49 : _GEN_8753; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8755 = 7'h32 == out_payload_rob_idx[6:0] ? rob_egress_id_50 : _GEN_8754; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8756 = 7'h33 == out_payload_rob_idx[6:0] ? rob_egress_id_51 : _GEN_8755; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8757 = 7'h34 == out_payload_rob_idx[6:0] ? rob_egress_id_52 : _GEN_8756; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8758 = 7'h35 == out_payload_rob_idx[6:0] ? rob_egress_id_53 : _GEN_8757; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8759 = 7'h36 == out_payload_rob_idx[6:0] ? rob_egress_id_54 : _GEN_8758; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8760 = 7'h37 == out_payload_rob_idx[6:0] ? rob_egress_id_55 : _GEN_8759; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8761 = 7'h38 == out_payload_rob_idx[6:0] ? rob_egress_id_56 : _GEN_8760; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8762 = 7'h39 == out_payload_rob_idx[6:0] ? rob_egress_id_57 : _GEN_8761; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8763 = 7'h3a == out_payload_rob_idx[6:0] ? rob_egress_id_58 : _GEN_8762; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8764 = 7'h3b == out_payload_rob_idx[6:0] ? rob_egress_id_59 : _GEN_8763; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8765 = 7'h3c == out_payload_rob_idx[6:0] ? rob_egress_id_60 : _GEN_8764; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8766 = 7'h3d == out_payload_rob_idx[6:0] ? rob_egress_id_61 : _GEN_8765; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8767 = 7'h3e == out_payload_rob_idx[6:0] ? rob_egress_id_62 : _GEN_8766; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8768 = 7'h3f == out_payload_rob_idx[6:0] ? rob_egress_id_63 : _GEN_8767; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8769 = 7'h40 == out_payload_rob_idx[6:0] ? rob_egress_id_64 : _GEN_8768; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8770 = 7'h41 == out_payload_rob_idx[6:0] ? rob_egress_id_65 : _GEN_8769; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8771 = 7'h42 == out_payload_rob_idx[6:0] ? rob_egress_id_66 : _GEN_8770; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8772 = 7'h43 == out_payload_rob_idx[6:0] ? rob_egress_id_67 : _GEN_8771; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8773 = 7'h44 == out_payload_rob_idx[6:0] ? rob_egress_id_68 : _GEN_8772; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8774 = 7'h45 == out_payload_rob_idx[6:0] ? rob_egress_id_69 : _GEN_8773; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8775 = 7'h46 == out_payload_rob_idx[6:0] ? rob_egress_id_70 : _GEN_8774; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8776 = 7'h47 == out_payload_rob_idx[6:0] ? rob_egress_id_71 : _GEN_8775; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8777 = 7'h48 == out_payload_rob_idx[6:0] ? rob_egress_id_72 : _GEN_8776; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8778 = 7'h49 == out_payload_rob_idx[6:0] ? rob_egress_id_73 : _GEN_8777; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8779 = 7'h4a == out_payload_rob_idx[6:0] ? rob_egress_id_74 : _GEN_8778; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8780 = 7'h4b == out_payload_rob_idx[6:0] ? rob_egress_id_75 : _GEN_8779; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8781 = 7'h4c == out_payload_rob_idx[6:0] ? rob_egress_id_76 : _GEN_8780; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8782 = 7'h4d == out_payload_rob_idx[6:0] ? rob_egress_id_77 : _GEN_8781; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8783 = 7'h4e == out_payload_rob_idx[6:0] ? rob_egress_id_78 : _GEN_8782; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8784 = 7'h4f == out_payload_rob_idx[6:0] ? rob_egress_id_79 : _GEN_8783; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8785 = 7'h50 == out_payload_rob_idx[6:0] ? rob_egress_id_80 : _GEN_8784; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8786 = 7'h51 == out_payload_rob_idx[6:0] ? rob_egress_id_81 : _GEN_8785; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8787 = 7'h52 == out_payload_rob_idx[6:0] ? rob_egress_id_82 : _GEN_8786; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8788 = 7'h53 == out_payload_rob_idx[6:0] ? rob_egress_id_83 : _GEN_8787; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8789 = 7'h54 == out_payload_rob_idx[6:0] ? rob_egress_id_84 : _GEN_8788; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8790 = 7'h55 == out_payload_rob_idx[6:0] ? rob_egress_id_85 : _GEN_8789; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8791 = 7'h56 == out_payload_rob_idx[6:0] ? rob_egress_id_86 : _GEN_8790; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8792 = 7'h57 == out_payload_rob_idx[6:0] ? rob_egress_id_87 : _GEN_8791; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8793 = 7'h58 == out_payload_rob_idx[6:0] ? rob_egress_id_88 : _GEN_8792; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8794 = 7'h59 == out_payload_rob_idx[6:0] ? rob_egress_id_89 : _GEN_8793; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8795 = 7'h5a == out_payload_rob_idx[6:0] ? rob_egress_id_90 : _GEN_8794; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8796 = 7'h5b == out_payload_rob_idx[6:0] ? rob_egress_id_91 : _GEN_8795; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8797 = 7'h5c == out_payload_rob_idx[6:0] ? rob_egress_id_92 : _GEN_8796; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8798 = 7'h5d == out_payload_rob_idx[6:0] ? rob_egress_id_93 : _GEN_8797; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8799 = 7'h5e == out_payload_rob_idx[6:0] ? rob_egress_id_94 : _GEN_8798; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8800 = 7'h5f == out_payload_rob_idx[6:0] ? rob_egress_id_95 : _GEN_8799; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8801 = 7'h60 == out_payload_rob_idx[6:0] ? rob_egress_id_96 : _GEN_8800; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8802 = 7'h61 == out_payload_rob_idx[6:0] ? rob_egress_id_97 : _GEN_8801; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8803 = 7'h62 == out_payload_rob_idx[6:0] ? rob_egress_id_98 : _GEN_8802; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8804 = 7'h63 == out_payload_rob_idx[6:0] ? rob_egress_id_99 : _GEN_8803; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8805 = 7'h64 == out_payload_rob_idx[6:0] ? rob_egress_id_100 : _GEN_8804; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8806 = 7'h65 == out_payload_rob_idx[6:0] ? rob_egress_id_101 : _GEN_8805; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8807 = 7'h66 == out_payload_rob_idx[6:0] ? rob_egress_id_102 : _GEN_8806; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8808 = 7'h67 == out_payload_rob_idx[6:0] ? rob_egress_id_103 : _GEN_8807; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8809 = 7'h68 == out_payload_rob_idx[6:0] ? rob_egress_id_104 : _GEN_8808; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8810 = 7'h69 == out_payload_rob_idx[6:0] ? rob_egress_id_105 : _GEN_8809; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8811 = 7'h6a == out_payload_rob_idx[6:0] ? rob_egress_id_106 : _GEN_8810; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8812 = 7'h6b == out_payload_rob_idx[6:0] ? rob_egress_id_107 : _GEN_8811; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8813 = 7'h6c == out_payload_rob_idx[6:0] ? rob_egress_id_108 : _GEN_8812; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8814 = 7'h6d == out_payload_rob_idx[6:0] ? rob_egress_id_109 : _GEN_8813; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8815 = 7'h6e == out_payload_rob_idx[6:0] ? rob_egress_id_110 : _GEN_8814; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8816 = 7'h6f == out_payload_rob_idx[6:0] ? rob_egress_id_111 : _GEN_8815; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8817 = 7'h70 == out_payload_rob_idx[6:0] ? rob_egress_id_112 : _GEN_8816; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8818 = 7'h71 == out_payload_rob_idx[6:0] ? rob_egress_id_113 : _GEN_8817; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8819 = 7'h72 == out_payload_rob_idx[6:0] ? rob_egress_id_114 : _GEN_8818; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8820 = 7'h73 == out_payload_rob_idx[6:0] ? rob_egress_id_115 : _GEN_8819; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8821 = 7'h74 == out_payload_rob_idx[6:0] ? rob_egress_id_116 : _GEN_8820; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8822 = 7'h75 == out_payload_rob_idx[6:0] ? rob_egress_id_117 : _GEN_8821; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8823 = 7'h76 == out_payload_rob_idx[6:0] ? rob_egress_id_118 : _GEN_8822; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8824 = 7'h77 == out_payload_rob_idx[6:0] ? rob_egress_id_119 : _GEN_8823; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8825 = 7'h78 == out_payload_rob_idx[6:0] ? rob_egress_id_120 : _GEN_8824; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8826 = 7'h79 == out_payload_rob_idx[6:0] ? rob_egress_id_121 : _GEN_8825; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8827 = 7'h7a == out_payload_rob_idx[6:0] ? rob_egress_id_122 : _GEN_8826; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8828 = 7'h7b == out_payload_rob_idx[6:0] ? rob_egress_id_123 : _GEN_8827; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8829 = 7'h7c == out_payload_rob_idx[6:0] ? rob_egress_id_124 : _GEN_8828; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8830 = 7'h7d == out_payload_rob_idx[6:0] ? rob_egress_id_125 : _GEN_8829; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8831 = 7'h7e == out_payload_rob_idx[6:0] ? rob_egress_id_126 : _GEN_8830; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_8832 = 7'h7f == out_payload_rob_idx[6:0] ? rob_egress_id_127 : _GEN_8831; // @[TestHarness.scala 204:{18,18}]
  wire [3:0] _GEN_8834 = 7'h1 == out_payload_rob_idx[6:0] ? rob_flits_returned_1 : rob_flits_returned_0; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8835 = 7'h2 == out_payload_rob_idx[6:0] ? rob_flits_returned_2 : _GEN_8834; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8836 = 7'h3 == out_payload_rob_idx[6:0] ? rob_flits_returned_3 : _GEN_8835; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8837 = 7'h4 == out_payload_rob_idx[6:0] ? rob_flits_returned_4 : _GEN_8836; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8838 = 7'h5 == out_payload_rob_idx[6:0] ? rob_flits_returned_5 : _GEN_8837; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8839 = 7'h6 == out_payload_rob_idx[6:0] ? rob_flits_returned_6 : _GEN_8838; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8840 = 7'h7 == out_payload_rob_idx[6:0] ? rob_flits_returned_7 : _GEN_8839; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8841 = 7'h8 == out_payload_rob_idx[6:0] ? rob_flits_returned_8 : _GEN_8840; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8842 = 7'h9 == out_payload_rob_idx[6:0] ? rob_flits_returned_9 : _GEN_8841; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8843 = 7'ha == out_payload_rob_idx[6:0] ? rob_flits_returned_10 : _GEN_8842; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8844 = 7'hb == out_payload_rob_idx[6:0] ? rob_flits_returned_11 : _GEN_8843; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8845 = 7'hc == out_payload_rob_idx[6:0] ? rob_flits_returned_12 : _GEN_8844; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8846 = 7'hd == out_payload_rob_idx[6:0] ? rob_flits_returned_13 : _GEN_8845; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8847 = 7'he == out_payload_rob_idx[6:0] ? rob_flits_returned_14 : _GEN_8846; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8848 = 7'hf == out_payload_rob_idx[6:0] ? rob_flits_returned_15 : _GEN_8847; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8849 = 7'h10 == out_payload_rob_idx[6:0] ? rob_flits_returned_16 : _GEN_8848; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8850 = 7'h11 == out_payload_rob_idx[6:0] ? rob_flits_returned_17 : _GEN_8849; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8851 = 7'h12 == out_payload_rob_idx[6:0] ? rob_flits_returned_18 : _GEN_8850; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8852 = 7'h13 == out_payload_rob_idx[6:0] ? rob_flits_returned_19 : _GEN_8851; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8853 = 7'h14 == out_payload_rob_idx[6:0] ? rob_flits_returned_20 : _GEN_8852; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8854 = 7'h15 == out_payload_rob_idx[6:0] ? rob_flits_returned_21 : _GEN_8853; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8855 = 7'h16 == out_payload_rob_idx[6:0] ? rob_flits_returned_22 : _GEN_8854; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8856 = 7'h17 == out_payload_rob_idx[6:0] ? rob_flits_returned_23 : _GEN_8855; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8857 = 7'h18 == out_payload_rob_idx[6:0] ? rob_flits_returned_24 : _GEN_8856; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8858 = 7'h19 == out_payload_rob_idx[6:0] ? rob_flits_returned_25 : _GEN_8857; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8859 = 7'h1a == out_payload_rob_idx[6:0] ? rob_flits_returned_26 : _GEN_8858; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8860 = 7'h1b == out_payload_rob_idx[6:0] ? rob_flits_returned_27 : _GEN_8859; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8861 = 7'h1c == out_payload_rob_idx[6:0] ? rob_flits_returned_28 : _GEN_8860; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8862 = 7'h1d == out_payload_rob_idx[6:0] ? rob_flits_returned_29 : _GEN_8861; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8863 = 7'h1e == out_payload_rob_idx[6:0] ? rob_flits_returned_30 : _GEN_8862; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8864 = 7'h1f == out_payload_rob_idx[6:0] ? rob_flits_returned_31 : _GEN_8863; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8865 = 7'h20 == out_payload_rob_idx[6:0] ? rob_flits_returned_32 : _GEN_8864; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8866 = 7'h21 == out_payload_rob_idx[6:0] ? rob_flits_returned_33 : _GEN_8865; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8867 = 7'h22 == out_payload_rob_idx[6:0] ? rob_flits_returned_34 : _GEN_8866; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8868 = 7'h23 == out_payload_rob_idx[6:0] ? rob_flits_returned_35 : _GEN_8867; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8869 = 7'h24 == out_payload_rob_idx[6:0] ? rob_flits_returned_36 : _GEN_8868; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8870 = 7'h25 == out_payload_rob_idx[6:0] ? rob_flits_returned_37 : _GEN_8869; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8871 = 7'h26 == out_payload_rob_idx[6:0] ? rob_flits_returned_38 : _GEN_8870; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8872 = 7'h27 == out_payload_rob_idx[6:0] ? rob_flits_returned_39 : _GEN_8871; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8873 = 7'h28 == out_payload_rob_idx[6:0] ? rob_flits_returned_40 : _GEN_8872; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8874 = 7'h29 == out_payload_rob_idx[6:0] ? rob_flits_returned_41 : _GEN_8873; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8875 = 7'h2a == out_payload_rob_idx[6:0] ? rob_flits_returned_42 : _GEN_8874; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8876 = 7'h2b == out_payload_rob_idx[6:0] ? rob_flits_returned_43 : _GEN_8875; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8877 = 7'h2c == out_payload_rob_idx[6:0] ? rob_flits_returned_44 : _GEN_8876; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8878 = 7'h2d == out_payload_rob_idx[6:0] ? rob_flits_returned_45 : _GEN_8877; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8879 = 7'h2e == out_payload_rob_idx[6:0] ? rob_flits_returned_46 : _GEN_8878; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8880 = 7'h2f == out_payload_rob_idx[6:0] ? rob_flits_returned_47 : _GEN_8879; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8881 = 7'h30 == out_payload_rob_idx[6:0] ? rob_flits_returned_48 : _GEN_8880; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8882 = 7'h31 == out_payload_rob_idx[6:0] ? rob_flits_returned_49 : _GEN_8881; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8883 = 7'h32 == out_payload_rob_idx[6:0] ? rob_flits_returned_50 : _GEN_8882; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8884 = 7'h33 == out_payload_rob_idx[6:0] ? rob_flits_returned_51 : _GEN_8883; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8885 = 7'h34 == out_payload_rob_idx[6:0] ? rob_flits_returned_52 : _GEN_8884; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8886 = 7'h35 == out_payload_rob_idx[6:0] ? rob_flits_returned_53 : _GEN_8885; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8887 = 7'h36 == out_payload_rob_idx[6:0] ? rob_flits_returned_54 : _GEN_8886; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8888 = 7'h37 == out_payload_rob_idx[6:0] ? rob_flits_returned_55 : _GEN_8887; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8889 = 7'h38 == out_payload_rob_idx[6:0] ? rob_flits_returned_56 : _GEN_8888; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8890 = 7'h39 == out_payload_rob_idx[6:0] ? rob_flits_returned_57 : _GEN_8889; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8891 = 7'h3a == out_payload_rob_idx[6:0] ? rob_flits_returned_58 : _GEN_8890; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8892 = 7'h3b == out_payload_rob_idx[6:0] ? rob_flits_returned_59 : _GEN_8891; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8893 = 7'h3c == out_payload_rob_idx[6:0] ? rob_flits_returned_60 : _GEN_8892; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8894 = 7'h3d == out_payload_rob_idx[6:0] ? rob_flits_returned_61 : _GEN_8893; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8895 = 7'h3e == out_payload_rob_idx[6:0] ? rob_flits_returned_62 : _GEN_8894; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8896 = 7'h3f == out_payload_rob_idx[6:0] ? rob_flits_returned_63 : _GEN_8895; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8897 = 7'h40 == out_payload_rob_idx[6:0] ? rob_flits_returned_64 : _GEN_8896; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8898 = 7'h41 == out_payload_rob_idx[6:0] ? rob_flits_returned_65 : _GEN_8897; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8899 = 7'h42 == out_payload_rob_idx[6:0] ? rob_flits_returned_66 : _GEN_8898; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8900 = 7'h43 == out_payload_rob_idx[6:0] ? rob_flits_returned_67 : _GEN_8899; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8901 = 7'h44 == out_payload_rob_idx[6:0] ? rob_flits_returned_68 : _GEN_8900; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8902 = 7'h45 == out_payload_rob_idx[6:0] ? rob_flits_returned_69 : _GEN_8901; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8903 = 7'h46 == out_payload_rob_idx[6:0] ? rob_flits_returned_70 : _GEN_8902; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8904 = 7'h47 == out_payload_rob_idx[6:0] ? rob_flits_returned_71 : _GEN_8903; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8905 = 7'h48 == out_payload_rob_idx[6:0] ? rob_flits_returned_72 : _GEN_8904; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8906 = 7'h49 == out_payload_rob_idx[6:0] ? rob_flits_returned_73 : _GEN_8905; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8907 = 7'h4a == out_payload_rob_idx[6:0] ? rob_flits_returned_74 : _GEN_8906; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8908 = 7'h4b == out_payload_rob_idx[6:0] ? rob_flits_returned_75 : _GEN_8907; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8909 = 7'h4c == out_payload_rob_idx[6:0] ? rob_flits_returned_76 : _GEN_8908; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8910 = 7'h4d == out_payload_rob_idx[6:0] ? rob_flits_returned_77 : _GEN_8909; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8911 = 7'h4e == out_payload_rob_idx[6:0] ? rob_flits_returned_78 : _GEN_8910; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8912 = 7'h4f == out_payload_rob_idx[6:0] ? rob_flits_returned_79 : _GEN_8911; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8913 = 7'h50 == out_payload_rob_idx[6:0] ? rob_flits_returned_80 : _GEN_8912; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8914 = 7'h51 == out_payload_rob_idx[6:0] ? rob_flits_returned_81 : _GEN_8913; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8915 = 7'h52 == out_payload_rob_idx[6:0] ? rob_flits_returned_82 : _GEN_8914; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8916 = 7'h53 == out_payload_rob_idx[6:0] ? rob_flits_returned_83 : _GEN_8915; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8917 = 7'h54 == out_payload_rob_idx[6:0] ? rob_flits_returned_84 : _GEN_8916; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8918 = 7'h55 == out_payload_rob_idx[6:0] ? rob_flits_returned_85 : _GEN_8917; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8919 = 7'h56 == out_payload_rob_idx[6:0] ? rob_flits_returned_86 : _GEN_8918; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8920 = 7'h57 == out_payload_rob_idx[6:0] ? rob_flits_returned_87 : _GEN_8919; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8921 = 7'h58 == out_payload_rob_idx[6:0] ? rob_flits_returned_88 : _GEN_8920; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8922 = 7'h59 == out_payload_rob_idx[6:0] ? rob_flits_returned_89 : _GEN_8921; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8923 = 7'h5a == out_payload_rob_idx[6:0] ? rob_flits_returned_90 : _GEN_8922; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8924 = 7'h5b == out_payload_rob_idx[6:0] ? rob_flits_returned_91 : _GEN_8923; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8925 = 7'h5c == out_payload_rob_idx[6:0] ? rob_flits_returned_92 : _GEN_8924; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8926 = 7'h5d == out_payload_rob_idx[6:0] ? rob_flits_returned_93 : _GEN_8925; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8927 = 7'h5e == out_payload_rob_idx[6:0] ? rob_flits_returned_94 : _GEN_8926; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8928 = 7'h5f == out_payload_rob_idx[6:0] ? rob_flits_returned_95 : _GEN_8927; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8929 = 7'h60 == out_payload_rob_idx[6:0] ? rob_flits_returned_96 : _GEN_8928; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8930 = 7'h61 == out_payload_rob_idx[6:0] ? rob_flits_returned_97 : _GEN_8929; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8931 = 7'h62 == out_payload_rob_idx[6:0] ? rob_flits_returned_98 : _GEN_8930; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8932 = 7'h63 == out_payload_rob_idx[6:0] ? rob_flits_returned_99 : _GEN_8931; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8933 = 7'h64 == out_payload_rob_idx[6:0] ? rob_flits_returned_100 : _GEN_8932; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8934 = 7'h65 == out_payload_rob_idx[6:0] ? rob_flits_returned_101 : _GEN_8933; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8935 = 7'h66 == out_payload_rob_idx[6:0] ? rob_flits_returned_102 : _GEN_8934; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8936 = 7'h67 == out_payload_rob_idx[6:0] ? rob_flits_returned_103 : _GEN_8935; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8937 = 7'h68 == out_payload_rob_idx[6:0] ? rob_flits_returned_104 : _GEN_8936; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8938 = 7'h69 == out_payload_rob_idx[6:0] ? rob_flits_returned_105 : _GEN_8937; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8939 = 7'h6a == out_payload_rob_idx[6:0] ? rob_flits_returned_106 : _GEN_8938; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8940 = 7'h6b == out_payload_rob_idx[6:0] ? rob_flits_returned_107 : _GEN_8939; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8941 = 7'h6c == out_payload_rob_idx[6:0] ? rob_flits_returned_108 : _GEN_8940; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8942 = 7'h6d == out_payload_rob_idx[6:0] ? rob_flits_returned_109 : _GEN_8941; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8943 = 7'h6e == out_payload_rob_idx[6:0] ? rob_flits_returned_110 : _GEN_8942; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8944 = 7'h6f == out_payload_rob_idx[6:0] ? rob_flits_returned_111 : _GEN_8943; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8945 = 7'h70 == out_payload_rob_idx[6:0] ? rob_flits_returned_112 : _GEN_8944; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8946 = 7'h71 == out_payload_rob_idx[6:0] ? rob_flits_returned_113 : _GEN_8945; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8947 = 7'h72 == out_payload_rob_idx[6:0] ? rob_flits_returned_114 : _GEN_8946; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8948 = 7'h73 == out_payload_rob_idx[6:0] ? rob_flits_returned_115 : _GEN_8947; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8949 = 7'h74 == out_payload_rob_idx[6:0] ? rob_flits_returned_116 : _GEN_8948; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8950 = 7'h75 == out_payload_rob_idx[6:0] ? rob_flits_returned_117 : _GEN_8949; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8951 = 7'h76 == out_payload_rob_idx[6:0] ? rob_flits_returned_118 : _GEN_8950; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8952 = 7'h77 == out_payload_rob_idx[6:0] ? rob_flits_returned_119 : _GEN_8951; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8953 = 7'h78 == out_payload_rob_idx[6:0] ? rob_flits_returned_120 : _GEN_8952; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8954 = 7'h79 == out_payload_rob_idx[6:0] ? rob_flits_returned_121 : _GEN_8953; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8955 = 7'h7a == out_payload_rob_idx[6:0] ? rob_flits_returned_122 : _GEN_8954; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8956 = 7'h7b == out_payload_rob_idx[6:0] ? rob_flits_returned_123 : _GEN_8955; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8957 = 7'h7c == out_payload_rob_idx[6:0] ? rob_flits_returned_124 : _GEN_8956; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8958 = 7'h7d == out_payload_rob_idx[6:0] ? rob_flits_returned_125 : _GEN_8957; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8959 = 7'h7e == out_payload_rob_idx[6:0] ? rob_flits_returned_126 : _GEN_8958; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8960 = 7'h7f == out_payload_rob_idx[6:0] ? rob_flits_returned_127 : _GEN_8959; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8962 = 7'h1 == out_payload_rob_idx[6:0] ? rob_n_flits_1 : rob_n_flits_0; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8963 = 7'h2 == out_payload_rob_idx[6:0] ? rob_n_flits_2 : _GEN_8962; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8964 = 7'h3 == out_payload_rob_idx[6:0] ? rob_n_flits_3 : _GEN_8963; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8965 = 7'h4 == out_payload_rob_idx[6:0] ? rob_n_flits_4 : _GEN_8964; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8966 = 7'h5 == out_payload_rob_idx[6:0] ? rob_n_flits_5 : _GEN_8965; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8967 = 7'h6 == out_payload_rob_idx[6:0] ? rob_n_flits_6 : _GEN_8966; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8968 = 7'h7 == out_payload_rob_idx[6:0] ? rob_n_flits_7 : _GEN_8967; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8969 = 7'h8 == out_payload_rob_idx[6:0] ? rob_n_flits_8 : _GEN_8968; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8970 = 7'h9 == out_payload_rob_idx[6:0] ? rob_n_flits_9 : _GEN_8969; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8971 = 7'ha == out_payload_rob_idx[6:0] ? rob_n_flits_10 : _GEN_8970; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8972 = 7'hb == out_payload_rob_idx[6:0] ? rob_n_flits_11 : _GEN_8971; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8973 = 7'hc == out_payload_rob_idx[6:0] ? rob_n_flits_12 : _GEN_8972; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8974 = 7'hd == out_payload_rob_idx[6:0] ? rob_n_flits_13 : _GEN_8973; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8975 = 7'he == out_payload_rob_idx[6:0] ? rob_n_flits_14 : _GEN_8974; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8976 = 7'hf == out_payload_rob_idx[6:0] ? rob_n_flits_15 : _GEN_8975; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8977 = 7'h10 == out_payload_rob_idx[6:0] ? rob_n_flits_16 : _GEN_8976; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8978 = 7'h11 == out_payload_rob_idx[6:0] ? rob_n_flits_17 : _GEN_8977; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8979 = 7'h12 == out_payload_rob_idx[6:0] ? rob_n_flits_18 : _GEN_8978; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8980 = 7'h13 == out_payload_rob_idx[6:0] ? rob_n_flits_19 : _GEN_8979; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8981 = 7'h14 == out_payload_rob_idx[6:0] ? rob_n_flits_20 : _GEN_8980; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8982 = 7'h15 == out_payload_rob_idx[6:0] ? rob_n_flits_21 : _GEN_8981; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8983 = 7'h16 == out_payload_rob_idx[6:0] ? rob_n_flits_22 : _GEN_8982; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8984 = 7'h17 == out_payload_rob_idx[6:0] ? rob_n_flits_23 : _GEN_8983; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8985 = 7'h18 == out_payload_rob_idx[6:0] ? rob_n_flits_24 : _GEN_8984; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8986 = 7'h19 == out_payload_rob_idx[6:0] ? rob_n_flits_25 : _GEN_8985; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8987 = 7'h1a == out_payload_rob_idx[6:0] ? rob_n_flits_26 : _GEN_8986; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8988 = 7'h1b == out_payload_rob_idx[6:0] ? rob_n_flits_27 : _GEN_8987; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8989 = 7'h1c == out_payload_rob_idx[6:0] ? rob_n_flits_28 : _GEN_8988; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8990 = 7'h1d == out_payload_rob_idx[6:0] ? rob_n_flits_29 : _GEN_8989; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8991 = 7'h1e == out_payload_rob_idx[6:0] ? rob_n_flits_30 : _GEN_8990; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8992 = 7'h1f == out_payload_rob_idx[6:0] ? rob_n_flits_31 : _GEN_8991; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8993 = 7'h20 == out_payload_rob_idx[6:0] ? rob_n_flits_32 : _GEN_8992; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8994 = 7'h21 == out_payload_rob_idx[6:0] ? rob_n_flits_33 : _GEN_8993; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8995 = 7'h22 == out_payload_rob_idx[6:0] ? rob_n_flits_34 : _GEN_8994; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8996 = 7'h23 == out_payload_rob_idx[6:0] ? rob_n_flits_35 : _GEN_8995; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8997 = 7'h24 == out_payload_rob_idx[6:0] ? rob_n_flits_36 : _GEN_8996; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8998 = 7'h25 == out_payload_rob_idx[6:0] ? rob_n_flits_37 : _GEN_8997; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_8999 = 7'h26 == out_payload_rob_idx[6:0] ? rob_n_flits_38 : _GEN_8998; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9000 = 7'h27 == out_payload_rob_idx[6:0] ? rob_n_flits_39 : _GEN_8999; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9001 = 7'h28 == out_payload_rob_idx[6:0] ? rob_n_flits_40 : _GEN_9000; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9002 = 7'h29 == out_payload_rob_idx[6:0] ? rob_n_flits_41 : _GEN_9001; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9003 = 7'h2a == out_payload_rob_idx[6:0] ? rob_n_flits_42 : _GEN_9002; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9004 = 7'h2b == out_payload_rob_idx[6:0] ? rob_n_flits_43 : _GEN_9003; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9005 = 7'h2c == out_payload_rob_idx[6:0] ? rob_n_flits_44 : _GEN_9004; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9006 = 7'h2d == out_payload_rob_idx[6:0] ? rob_n_flits_45 : _GEN_9005; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9007 = 7'h2e == out_payload_rob_idx[6:0] ? rob_n_flits_46 : _GEN_9006; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9008 = 7'h2f == out_payload_rob_idx[6:0] ? rob_n_flits_47 : _GEN_9007; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9009 = 7'h30 == out_payload_rob_idx[6:0] ? rob_n_flits_48 : _GEN_9008; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9010 = 7'h31 == out_payload_rob_idx[6:0] ? rob_n_flits_49 : _GEN_9009; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9011 = 7'h32 == out_payload_rob_idx[6:0] ? rob_n_flits_50 : _GEN_9010; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9012 = 7'h33 == out_payload_rob_idx[6:0] ? rob_n_flits_51 : _GEN_9011; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9013 = 7'h34 == out_payload_rob_idx[6:0] ? rob_n_flits_52 : _GEN_9012; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9014 = 7'h35 == out_payload_rob_idx[6:0] ? rob_n_flits_53 : _GEN_9013; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9015 = 7'h36 == out_payload_rob_idx[6:0] ? rob_n_flits_54 : _GEN_9014; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9016 = 7'h37 == out_payload_rob_idx[6:0] ? rob_n_flits_55 : _GEN_9015; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9017 = 7'h38 == out_payload_rob_idx[6:0] ? rob_n_flits_56 : _GEN_9016; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9018 = 7'h39 == out_payload_rob_idx[6:0] ? rob_n_flits_57 : _GEN_9017; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9019 = 7'h3a == out_payload_rob_idx[6:0] ? rob_n_flits_58 : _GEN_9018; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9020 = 7'h3b == out_payload_rob_idx[6:0] ? rob_n_flits_59 : _GEN_9019; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9021 = 7'h3c == out_payload_rob_idx[6:0] ? rob_n_flits_60 : _GEN_9020; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9022 = 7'h3d == out_payload_rob_idx[6:0] ? rob_n_flits_61 : _GEN_9021; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9023 = 7'h3e == out_payload_rob_idx[6:0] ? rob_n_flits_62 : _GEN_9022; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9024 = 7'h3f == out_payload_rob_idx[6:0] ? rob_n_flits_63 : _GEN_9023; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9025 = 7'h40 == out_payload_rob_idx[6:0] ? rob_n_flits_64 : _GEN_9024; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9026 = 7'h41 == out_payload_rob_idx[6:0] ? rob_n_flits_65 : _GEN_9025; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9027 = 7'h42 == out_payload_rob_idx[6:0] ? rob_n_flits_66 : _GEN_9026; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9028 = 7'h43 == out_payload_rob_idx[6:0] ? rob_n_flits_67 : _GEN_9027; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9029 = 7'h44 == out_payload_rob_idx[6:0] ? rob_n_flits_68 : _GEN_9028; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9030 = 7'h45 == out_payload_rob_idx[6:0] ? rob_n_flits_69 : _GEN_9029; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9031 = 7'h46 == out_payload_rob_idx[6:0] ? rob_n_flits_70 : _GEN_9030; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9032 = 7'h47 == out_payload_rob_idx[6:0] ? rob_n_flits_71 : _GEN_9031; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9033 = 7'h48 == out_payload_rob_idx[6:0] ? rob_n_flits_72 : _GEN_9032; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9034 = 7'h49 == out_payload_rob_idx[6:0] ? rob_n_flits_73 : _GEN_9033; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9035 = 7'h4a == out_payload_rob_idx[6:0] ? rob_n_flits_74 : _GEN_9034; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9036 = 7'h4b == out_payload_rob_idx[6:0] ? rob_n_flits_75 : _GEN_9035; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9037 = 7'h4c == out_payload_rob_idx[6:0] ? rob_n_flits_76 : _GEN_9036; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9038 = 7'h4d == out_payload_rob_idx[6:0] ? rob_n_flits_77 : _GEN_9037; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9039 = 7'h4e == out_payload_rob_idx[6:0] ? rob_n_flits_78 : _GEN_9038; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9040 = 7'h4f == out_payload_rob_idx[6:0] ? rob_n_flits_79 : _GEN_9039; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9041 = 7'h50 == out_payload_rob_idx[6:0] ? rob_n_flits_80 : _GEN_9040; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9042 = 7'h51 == out_payload_rob_idx[6:0] ? rob_n_flits_81 : _GEN_9041; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9043 = 7'h52 == out_payload_rob_idx[6:0] ? rob_n_flits_82 : _GEN_9042; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9044 = 7'h53 == out_payload_rob_idx[6:0] ? rob_n_flits_83 : _GEN_9043; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9045 = 7'h54 == out_payload_rob_idx[6:0] ? rob_n_flits_84 : _GEN_9044; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9046 = 7'h55 == out_payload_rob_idx[6:0] ? rob_n_flits_85 : _GEN_9045; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9047 = 7'h56 == out_payload_rob_idx[6:0] ? rob_n_flits_86 : _GEN_9046; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9048 = 7'h57 == out_payload_rob_idx[6:0] ? rob_n_flits_87 : _GEN_9047; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9049 = 7'h58 == out_payload_rob_idx[6:0] ? rob_n_flits_88 : _GEN_9048; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9050 = 7'h59 == out_payload_rob_idx[6:0] ? rob_n_flits_89 : _GEN_9049; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9051 = 7'h5a == out_payload_rob_idx[6:0] ? rob_n_flits_90 : _GEN_9050; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9052 = 7'h5b == out_payload_rob_idx[6:0] ? rob_n_flits_91 : _GEN_9051; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9053 = 7'h5c == out_payload_rob_idx[6:0] ? rob_n_flits_92 : _GEN_9052; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9054 = 7'h5d == out_payload_rob_idx[6:0] ? rob_n_flits_93 : _GEN_9053; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9055 = 7'h5e == out_payload_rob_idx[6:0] ? rob_n_flits_94 : _GEN_9054; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9056 = 7'h5f == out_payload_rob_idx[6:0] ? rob_n_flits_95 : _GEN_9055; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9057 = 7'h60 == out_payload_rob_idx[6:0] ? rob_n_flits_96 : _GEN_9056; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9058 = 7'h61 == out_payload_rob_idx[6:0] ? rob_n_flits_97 : _GEN_9057; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9059 = 7'h62 == out_payload_rob_idx[6:0] ? rob_n_flits_98 : _GEN_9058; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9060 = 7'h63 == out_payload_rob_idx[6:0] ? rob_n_flits_99 : _GEN_9059; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9061 = 7'h64 == out_payload_rob_idx[6:0] ? rob_n_flits_100 : _GEN_9060; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9062 = 7'h65 == out_payload_rob_idx[6:0] ? rob_n_flits_101 : _GEN_9061; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9063 = 7'h66 == out_payload_rob_idx[6:0] ? rob_n_flits_102 : _GEN_9062; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9064 = 7'h67 == out_payload_rob_idx[6:0] ? rob_n_flits_103 : _GEN_9063; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9065 = 7'h68 == out_payload_rob_idx[6:0] ? rob_n_flits_104 : _GEN_9064; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9066 = 7'h69 == out_payload_rob_idx[6:0] ? rob_n_flits_105 : _GEN_9065; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9067 = 7'h6a == out_payload_rob_idx[6:0] ? rob_n_flits_106 : _GEN_9066; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9068 = 7'h6b == out_payload_rob_idx[6:0] ? rob_n_flits_107 : _GEN_9067; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9069 = 7'h6c == out_payload_rob_idx[6:0] ? rob_n_flits_108 : _GEN_9068; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9070 = 7'h6d == out_payload_rob_idx[6:0] ? rob_n_flits_109 : _GEN_9069; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9071 = 7'h6e == out_payload_rob_idx[6:0] ? rob_n_flits_110 : _GEN_9070; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9072 = 7'h6f == out_payload_rob_idx[6:0] ? rob_n_flits_111 : _GEN_9071; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9073 = 7'h70 == out_payload_rob_idx[6:0] ? rob_n_flits_112 : _GEN_9072; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9074 = 7'h71 == out_payload_rob_idx[6:0] ? rob_n_flits_113 : _GEN_9073; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9075 = 7'h72 == out_payload_rob_idx[6:0] ? rob_n_flits_114 : _GEN_9074; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9076 = 7'h73 == out_payload_rob_idx[6:0] ? rob_n_flits_115 : _GEN_9075; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9077 = 7'h74 == out_payload_rob_idx[6:0] ? rob_n_flits_116 : _GEN_9076; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9078 = 7'h75 == out_payload_rob_idx[6:0] ? rob_n_flits_117 : _GEN_9077; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9079 = 7'h76 == out_payload_rob_idx[6:0] ? rob_n_flits_118 : _GEN_9078; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9080 = 7'h77 == out_payload_rob_idx[6:0] ? rob_n_flits_119 : _GEN_9079; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9081 = 7'h78 == out_payload_rob_idx[6:0] ? rob_n_flits_120 : _GEN_9080; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9082 = 7'h79 == out_payload_rob_idx[6:0] ? rob_n_flits_121 : _GEN_9081; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9083 = 7'h7a == out_payload_rob_idx[6:0] ? rob_n_flits_122 : _GEN_9082; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9084 = 7'h7b == out_payload_rob_idx[6:0] ? rob_n_flits_123 : _GEN_9083; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9085 = 7'h7c == out_payload_rob_idx[6:0] ? rob_n_flits_124 : _GEN_9084; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9086 = 7'h7d == out_payload_rob_idx[6:0] ? rob_n_flits_125 : _GEN_9085; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9087 = 7'h7e == out_payload_rob_idx[6:0] ? rob_n_flits_126 : _GEN_9086; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_9088 = 7'h7f == out_payload_rob_idx[6:0] ? rob_n_flits_127 : _GEN_9087; // @[TestHarness.scala 205:{42,42}]
  wire [15:0] _GEN_15381 = {{9'd0}, packet_rob_idx}; // @[TestHarness.scala 206:61]
  wire  _T_110 = io_from_noc_0_flit_bits_head & enable_print_latency; // @[TestHarness.scala 208:30]
  wire [3:0] _rob_flits_returned_T_2 = _GEN_8960 + 4'h1; // @[TestHarness.scala 213:66]
  wire [3:0] _GEN_9345 = 7'h0 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7937; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9346 = 7'h1 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7938; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9347 = 7'h2 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7939; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9348 = 7'h3 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7940; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9349 = 7'h4 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7941; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9350 = 7'h5 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7942; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9351 = 7'h6 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7943; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9352 = 7'h7 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7944; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9353 = 7'h8 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7945; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9354 = 7'h9 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7946; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9355 = 7'ha == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7947; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9356 = 7'hb == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7948; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9357 = 7'hc == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7949; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9358 = 7'hd == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7950; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9359 = 7'he == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7951; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9360 = 7'hf == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7952; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9361 = 7'h10 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7953; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9362 = 7'h11 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7954; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9363 = 7'h12 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7955; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9364 = 7'h13 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7956; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9365 = 7'h14 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7957; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9366 = 7'h15 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7958; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9367 = 7'h16 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7959; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9368 = 7'h17 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7960; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9369 = 7'h18 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7961; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9370 = 7'h19 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7962; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9371 = 7'h1a == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7963; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9372 = 7'h1b == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7964; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9373 = 7'h1c == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7965; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9374 = 7'h1d == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7966; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9375 = 7'h1e == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7967; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9376 = 7'h1f == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7968; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9377 = 7'h20 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7969; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9378 = 7'h21 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7970; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9379 = 7'h22 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7971; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9380 = 7'h23 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7972; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9381 = 7'h24 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7973; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9382 = 7'h25 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7974; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9383 = 7'h26 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7975; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9384 = 7'h27 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7976; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9385 = 7'h28 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7977; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9386 = 7'h29 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7978; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9387 = 7'h2a == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7979; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9388 = 7'h2b == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7980; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9389 = 7'h2c == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7981; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9390 = 7'h2d == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7982; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9391 = 7'h2e == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7983; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9392 = 7'h2f == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7984; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9393 = 7'h30 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7985; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9394 = 7'h31 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7986; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9395 = 7'h32 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7987; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9396 = 7'h33 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7988; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9397 = 7'h34 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7989; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9398 = 7'h35 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7990; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9399 = 7'h36 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7991; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9400 = 7'h37 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7992; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9401 = 7'h38 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7993; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9402 = 7'h39 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7994; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9403 = 7'h3a == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7995; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9404 = 7'h3b == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7996; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9405 = 7'h3c == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7997; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9406 = 7'h3d == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7998; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9407 = 7'h3e == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_7999; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9408 = 7'h3f == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8000; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9409 = 7'h40 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8001; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9410 = 7'h41 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8002; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9411 = 7'h42 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8003; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9412 = 7'h43 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8004; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9413 = 7'h44 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8005; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9414 = 7'h45 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8006; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9415 = 7'h46 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8007; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9416 = 7'h47 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8008; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9417 = 7'h48 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8009; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9418 = 7'h49 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8010; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9419 = 7'h4a == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8011; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9420 = 7'h4b == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8012; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9421 = 7'h4c == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8013; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9422 = 7'h4d == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8014; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9423 = 7'h4e == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8015; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9424 = 7'h4f == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8016; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9425 = 7'h50 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8017; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9426 = 7'h51 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8018; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9427 = 7'h52 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8019; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9428 = 7'h53 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8020; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9429 = 7'h54 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8021; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9430 = 7'h55 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8022; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9431 = 7'h56 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8023; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9432 = 7'h57 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8024; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9433 = 7'h58 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8025; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9434 = 7'h59 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8026; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9435 = 7'h5a == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8027; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9436 = 7'h5b == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8028; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9437 = 7'h5c == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8029; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9438 = 7'h5d == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8030; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9439 = 7'h5e == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8031; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9440 = 7'h5f == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8032; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9441 = 7'h60 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8033; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9442 = 7'h61 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8034; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9443 = 7'h62 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8035; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9444 = 7'h63 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8036; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9445 = 7'h64 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8037; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9446 = 7'h65 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8038; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9447 = 7'h66 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8039; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9448 = 7'h67 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8040; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9449 = 7'h68 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8041; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9450 = 7'h69 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8042; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9451 = 7'h6a == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8043; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9452 = 7'h6b == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8044; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9453 = 7'h6c == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8045; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9454 = 7'h6d == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8046; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9455 = 7'h6e == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8047; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9456 = 7'h6f == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8048; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9457 = 7'h70 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8049; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9458 = 7'h71 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8050; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9459 = 7'h72 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8051; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9460 = 7'h73 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8052; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9461 = 7'h74 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8053; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9462 = 7'h75 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8054; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9463 = 7'h76 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8055; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9464 = 7'h77 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8056; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9465 = 7'h78 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8057; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9466 = 7'h79 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8058; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9467 = 7'h7a == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8059; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9468 = 7'h7b == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8060; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9469 = 7'h7c == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8061; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9470 = 7'h7d == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8062; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9471 = 7'h7e == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8063; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_9472 = 7'h7f == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_8064; // @[TestHarness.scala 213:{35,35}]
  wire [15:0] _rob_payload_flits_fired_T_2 = _GEN_8576 + 16'h1; // @[TestHarness.scala 214:76]
  wire [15:0] _GEN_9601 = 7'h0 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7425; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9602 = 7'h1 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7426; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9603 = 7'h2 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7427; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9604 = 7'h3 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7428; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9605 = 7'h4 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7429; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9606 = 7'h5 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7430; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9607 = 7'h6 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7431; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9608 = 7'h7 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7432; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9609 = 7'h8 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7433; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9610 = 7'h9 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7434; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9611 = 7'ha == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7435; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9612 = 7'hb == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7436; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9613 = 7'hc == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7437; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9614 = 7'hd == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7438; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9615 = 7'he == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7439; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9616 = 7'hf == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7440; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9617 = 7'h10 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7441; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9618 = 7'h11 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7442; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9619 = 7'h12 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7443; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9620 = 7'h13 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7444; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9621 = 7'h14 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7445; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9622 = 7'h15 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7446; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9623 = 7'h16 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7447; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9624 = 7'h17 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7448; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9625 = 7'h18 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7449; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9626 = 7'h19 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7450; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9627 = 7'h1a == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7451; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9628 = 7'h1b == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7452; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9629 = 7'h1c == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7453; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9630 = 7'h1d == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7454; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9631 = 7'h1e == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7455; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9632 = 7'h1f == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7456; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9633 = 7'h20 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7457; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9634 = 7'h21 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7458; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9635 = 7'h22 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7459; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9636 = 7'h23 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7460; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9637 = 7'h24 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7461; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9638 = 7'h25 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7462; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9639 = 7'h26 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7463; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9640 = 7'h27 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7464; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9641 = 7'h28 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7465; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9642 = 7'h29 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7466; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9643 = 7'h2a == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7467; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9644 = 7'h2b == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7468; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9645 = 7'h2c == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7469; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9646 = 7'h2d == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7470; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9647 = 7'h2e == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7471; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9648 = 7'h2f == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7472; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9649 = 7'h30 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7473; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9650 = 7'h31 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7474; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9651 = 7'h32 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7475; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9652 = 7'h33 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7476; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9653 = 7'h34 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7477; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9654 = 7'h35 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7478; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9655 = 7'h36 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7479; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9656 = 7'h37 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7480; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9657 = 7'h38 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7481; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9658 = 7'h39 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7482; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9659 = 7'h3a == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7483; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9660 = 7'h3b == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7484; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9661 = 7'h3c == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7485; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9662 = 7'h3d == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7486; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9663 = 7'h3e == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7487; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9664 = 7'h3f == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7488; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9665 = 7'h40 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7489; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9666 = 7'h41 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7490; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9667 = 7'h42 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7491; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9668 = 7'h43 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7492; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9669 = 7'h44 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7493; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9670 = 7'h45 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7494; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9671 = 7'h46 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7495; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9672 = 7'h47 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7496; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9673 = 7'h48 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7497; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9674 = 7'h49 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7498; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9675 = 7'h4a == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7499; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9676 = 7'h4b == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7500; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9677 = 7'h4c == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7501; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9678 = 7'h4d == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7502; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9679 = 7'h4e == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7503; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9680 = 7'h4f == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7504; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9681 = 7'h50 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7505; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9682 = 7'h51 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7506; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9683 = 7'h52 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7507; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9684 = 7'h53 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7508; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9685 = 7'h54 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7509; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9686 = 7'h55 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7510; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9687 = 7'h56 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7511; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9688 = 7'h57 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7512; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9689 = 7'h58 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7513; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9690 = 7'h59 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7514; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9691 = 7'h5a == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7515; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9692 = 7'h5b == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7516; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9693 = 7'h5c == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7517; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9694 = 7'h5d == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7518; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9695 = 7'h5e == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7519; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9696 = 7'h5f == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7520; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9697 = 7'h60 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7521; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9698 = 7'h61 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7522; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9699 = 7'h62 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7523; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9700 = 7'h63 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7524; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9701 = 7'h64 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7525; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9702 = 7'h65 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7526; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9703 = 7'h66 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7527; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9704 = 7'h67 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7528; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9705 = 7'h68 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7529; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9706 = 7'h69 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7530; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9707 = 7'h6a == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7531; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9708 = 7'h6b == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7532; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9709 = 7'h6c == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7533; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9710 = 7'h6d == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7534; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9711 = 7'h6e == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7535; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9712 = 7'h6f == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7536; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9713 = 7'h70 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7537; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9714 = 7'h71 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7538; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9715 = 7'h72 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7539; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9716 = 7'h73 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7540; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9717 = 7'h74 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7541; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9718 = 7'h75 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7542; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9719 = 7'h76 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7543; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9720 = 7'h77 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7544; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9721 = 7'h78 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7545; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9722 = 7'h79 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7546; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9723 = 7'h7a == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7547; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9724 = 7'h7b == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7548; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9725 = 7'h7c == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7549; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9726 = 7'h7d == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7550; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9727 = 7'h7e == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7551; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_9728 = 7'h7f == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_7552; // @[TestHarness.scala 214:{40,40}]
  wire  _GEN_9729 = io_from_noc_0_flit_bits_head | packet_valid; // @[TestHarness.scala 196:31 215:{31,46}]
  wire [15:0] _GEN_9730 = io_from_noc_0_flit_bits_head ? out_payload_rob_idx : {{9'd0}, packet_rob_idx}; // @[TestHarness.scala 197:29 215:{31,72}]
  wire [3:0] _GEN_9732 = _T_118 ? _GEN_9345 : _GEN_7937; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9733 = _T_118 ? _GEN_9346 : _GEN_7938; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9734 = _T_118 ? _GEN_9347 : _GEN_7939; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9735 = _T_118 ? _GEN_9348 : _GEN_7940; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9736 = _T_118 ? _GEN_9349 : _GEN_7941; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9737 = _T_118 ? _GEN_9350 : _GEN_7942; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9738 = _T_118 ? _GEN_9351 : _GEN_7943; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9739 = _T_118 ? _GEN_9352 : _GEN_7944; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9740 = _T_118 ? _GEN_9353 : _GEN_7945; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9741 = _T_118 ? _GEN_9354 : _GEN_7946; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9742 = _T_118 ? _GEN_9355 : _GEN_7947; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9743 = _T_118 ? _GEN_9356 : _GEN_7948; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9744 = _T_118 ? _GEN_9357 : _GEN_7949; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9745 = _T_118 ? _GEN_9358 : _GEN_7950; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9746 = _T_118 ? _GEN_9359 : _GEN_7951; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9747 = _T_118 ? _GEN_9360 : _GEN_7952; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9748 = _T_118 ? _GEN_9361 : _GEN_7953; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9749 = _T_118 ? _GEN_9362 : _GEN_7954; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9750 = _T_118 ? _GEN_9363 : _GEN_7955; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9751 = _T_118 ? _GEN_9364 : _GEN_7956; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9752 = _T_118 ? _GEN_9365 : _GEN_7957; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9753 = _T_118 ? _GEN_9366 : _GEN_7958; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9754 = _T_118 ? _GEN_9367 : _GEN_7959; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9755 = _T_118 ? _GEN_9368 : _GEN_7960; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9756 = _T_118 ? _GEN_9369 : _GEN_7961; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9757 = _T_118 ? _GEN_9370 : _GEN_7962; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9758 = _T_118 ? _GEN_9371 : _GEN_7963; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9759 = _T_118 ? _GEN_9372 : _GEN_7964; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9760 = _T_118 ? _GEN_9373 : _GEN_7965; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9761 = _T_118 ? _GEN_9374 : _GEN_7966; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9762 = _T_118 ? _GEN_9375 : _GEN_7967; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9763 = _T_118 ? _GEN_9376 : _GEN_7968; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9764 = _T_118 ? _GEN_9377 : _GEN_7969; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9765 = _T_118 ? _GEN_9378 : _GEN_7970; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9766 = _T_118 ? _GEN_9379 : _GEN_7971; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9767 = _T_118 ? _GEN_9380 : _GEN_7972; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9768 = _T_118 ? _GEN_9381 : _GEN_7973; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9769 = _T_118 ? _GEN_9382 : _GEN_7974; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9770 = _T_118 ? _GEN_9383 : _GEN_7975; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9771 = _T_118 ? _GEN_9384 : _GEN_7976; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9772 = _T_118 ? _GEN_9385 : _GEN_7977; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9773 = _T_118 ? _GEN_9386 : _GEN_7978; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9774 = _T_118 ? _GEN_9387 : _GEN_7979; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9775 = _T_118 ? _GEN_9388 : _GEN_7980; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9776 = _T_118 ? _GEN_9389 : _GEN_7981; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9777 = _T_118 ? _GEN_9390 : _GEN_7982; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9778 = _T_118 ? _GEN_9391 : _GEN_7983; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9779 = _T_118 ? _GEN_9392 : _GEN_7984; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9780 = _T_118 ? _GEN_9393 : _GEN_7985; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9781 = _T_118 ? _GEN_9394 : _GEN_7986; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9782 = _T_118 ? _GEN_9395 : _GEN_7987; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9783 = _T_118 ? _GEN_9396 : _GEN_7988; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9784 = _T_118 ? _GEN_9397 : _GEN_7989; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9785 = _T_118 ? _GEN_9398 : _GEN_7990; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9786 = _T_118 ? _GEN_9399 : _GEN_7991; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9787 = _T_118 ? _GEN_9400 : _GEN_7992; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9788 = _T_118 ? _GEN_9401 : _GEN_7993; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9789 = _T_118 ? _GEN_9402 : _GEN_7994; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9790 = _T_118 ? _GEN_9403 : _GEN_7995; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9791 = _T_118 ? _GEN_9404 : _GEN_7996; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9792 = _T_118 ? _GEN_9405 : _GEN_7997; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9793 = _T_118 ? _GEN_9406 : _GEN_7998; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9794 = _T_118 ? _GEN_9407 : _GEN_7999; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9795 = _T_118 ? _GEN_9408 : _GEN_8000; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9796 = _T_118 ? _GEN_9409 : _GEN_8001; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9797 = _T_118 ? _GEN_9410 : _GEN_8002; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9798 = _T_118 ? _GEN_9411 : _GEN_8003; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9799 = _T_118 ? _GEN_9412 : _GEN_8004; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9800 = _T_118 ? _GEN_9413 : _GEN_8005; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9801 = _T_118 ? _GEN_9414 : _GEN_8006; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9802 = _T_118 ? _GEN_9415 : _GEN_8007; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9803 = _T_118 ? _GEN_9416 : _GEN_8008; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9804 = _T_118 ? _GEN_9417 : _GEN_8009; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9805 = _T_118 ? _GEN_9418 : _GEN_8010; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9806 = _T_118 ? _GEN_9419 : _GEN_8011; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9807 = _T_118 ? _GEN_9420 : _GEN_8012; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9808 = _T_118 ? _GEN_9421 : _GEN_8013; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9809 = _T_118 ? _GEN_9422 : _GEN_8014; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9810 = _T_118 ? _GEN_9423 : _GEN_8015; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9811 = _T_118 ? _GEN_9424 : _GEN_8016; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9812 = _T_118 ? _GEN_9425 : _GEN_8017; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9813 = _T_118 ? _GEN_9426 : _GEN_8018; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9814 = _T_118 ? _GEN_9427 : _GEN_8019; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9815 = _T_118 ? _GEN_9428 : _GEN_8020; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9816 = _T_118 ? _GEN_9429 : _GEN_8021; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9817 = _T_118 ? _GEN_9430 : _GEN_8022; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9818 = _T_118 ? _GEN_9431 : _GEN_8023; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9819 = _T_118 ? _GEN_9432 : _GEN_8024; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9820 = _T_118 ? _GEN_9433 : _GEN_8025; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9821 = _T_118 ? _GEN_9434 : _GEN_8026; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9822 = _T_118 ? _GEN_9435 : _GEN_8027; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9823 = _T_118 ? _GEN_9436 : _GEN_8028; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9824 = _T_118 ? _GEN_9437 : _GEN_8029; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9825 = _T_118 ? _GEN_9438 : _GEN_8030; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9826 = _T_118 ? _GEN_9439 : _GEN_8031; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9827 = _T_118 ? _GEN_9440 : _GEN_8032; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9828 = _T_118 ? _GEN_9441 : _GEN_8033; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9829 = _T_118 ? _GEN_9442 : _GEN_8034; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9830 = _T_118 ? _GEN_9443 : _GEN_8035; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9831 = _T_118 ? _GEN_9444 : _GEN_8036; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9832 = _T_118 ? _GEN_9445 : _GEN_8037; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9833 = _T_118 ? _GEN_9446 : _GEN_8038; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9834 = _T_118 ? _GEN_9447 : _GEN_8039; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9835 = _T_118 ? _GEN_9448 : _GEN_8040; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9836 = _T_118 ? _GEN_9449 : _GEN_8041; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9837 = _T_118 ? _GEN_9450 : _GEN_8042; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9838 = _T_118 ? _GEN_9451 : _GEN_8043; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9839 = _T_118 ? _GEN_9452 : _GEN_8044; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9840 = _T_118 ? _GEN_9453 : _GEN_8045; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9841 = _T_118 ? _GEN_9454 : _GEN_8046; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9842 = _T_118 ? _GEN_9455 : _GEN_8047; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9843 = _T_118 ? _GEN_9456 : _GEN_8048; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9844 = _T_118 ? _GEN_9457 : _GEN_8049; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9845 = _T_118 ? _GEN_9458 : _GEN_8050; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9846 = _T_118 ? _GEN_9459 : _GEN_8051; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9847 = _T_118 ? _GEN_9460 : _GEN_8052; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9848 = _T_118 ? _GEN_9461 : _GEN_8053; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9849 = _T_118 ? _GEN_9462 : _GEN_8054; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9850 = _T_118 ? _GEN_9463 : _GEN_8055; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9851 = _T_118 ? _GEN_9464 : _GEN_8056; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9852 = _T_118 ? _GEN_9465 : _GEN_8057; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9853 = _T_118 ? _GEN_9466 : _GEN_8058; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9854 = _T_118 ? _GEN_9467 : _GEN_8059; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9855 = _T_118 ? _GEN_9468 : _GEN_8060; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9856 = _T_118 ? _GEN_9469 : _GEN_8061; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9857 = _T_118 ? _GEN_9470 : _GEN_8062; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9858 = _T_118 ? _GEN_9471 : _GEN_8063; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_9859 = _T_118 ? _GEN_9472 : _GEN_8064; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9860 = _T_118 ? _GEN_9601 : _GEN_7425; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9861 = _T_118 ? _GEN_9602 : _GEN_7426; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9862 = _T_118 ? _GEN_9603 : _GEN_7427; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9863 = _T_118 ? _GEN_9604 : _GEN_7428; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9864 = _T_118 ? _GEN_9605 : _GEN_7429; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9865 = _T_118 ? _GEN_9606 : _GEN_7430; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9866 = _T_118 ? _GEN_9607 : _GEN_7431; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9867 = _T_118 ? _GEN_9608 : _GEN_7432; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9868 = _T_118 ? _GEN_9609 : _GEN_7433; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9869 = _T_118 ? _GEN_9610 : _GEN_7434; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9870 = _T_118 ? _GEN_9611 : _GEN_7435; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9871 = _T_118 ? _GEN_9612 : _GEN_7436; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9872 = _T_118 ? _GEN_9613 : _GEN_7437; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9873 = _T_118 ? _GEN_9614 : _GEN_7438; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9874 = _T_118 ? _GEN_9615 : _GEN_7439; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9875 = _T_118 ? _GEN_9616 : _GEN_7440; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9876 = _T_118 ? _GEN_9617 : _GEN_7441; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9877 = _T_118 ? _GEN_9618 : _GEN_7442; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9878 = _T_118 ? _GEN_9619 : _GEN_7443; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9879 = _T_118 ? _GEN_9620 : _GEN_7444; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9880 = _T_118 ? _GEN_9621 : _GEN_7445; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9881 = _T_118 ? _GEN_9622 : _GEN_7446; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9882 = _T_118 ? _GEN_9623 : _GEN_7447; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9883 = _T_118 ? _GEN_9624 : _GEN_7448; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9884 = _T_118 ? _GEN_9625 : _GEN_7449; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9885 = _T_118 ? _GEN_9626 : _GEN_7450; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9886 = _T_118 ? _GEN_9627 : _GEN_7451; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9887 = _T_118 ? _GEN_9628 : _GEN_7452; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9888 = _T_118 ? _GEN_9629 : _GEN_7453; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9889 = _T_118 ? _GEN_9630 : _GEN_7454; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9890 = _T_118 ? _GEN_9631 : _GEN_7455; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9891 = _T_118 ? _GEN_9632 : _GEN_7456; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9892 = _T_118 ? _GEN_9633 : _GEN_7457; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9893 = _T_118 ? _GEN_9634 : _GEN_7458; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9894 = _T_118 ? _GEN_9635 : _GEN_7459; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9895 = _T_118 ? _GEN_9636 : _GEN_7460; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9896 = _T_118 ? _GEN_9637 : _GEN_7461; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9897 = _T_118 ? _GEN_9638 : _GEN_7462; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9898 = _T_118 ? _GEN_9639 : _GEN_7463; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9899 = _T_118 ? _GEN_9640 : _GEN_7464; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9900 = _T_118 ? _GEN_9641 : _GEN_7465; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9901 = _T_118 ? _GEN_9642 : _GEN_7466; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9902 = _T_118 ? _GEN_9643 : _GEN_7467; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9903 = _T_118 ? _GEN_9644 : _GEN_7468; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9904 = _T_118 ? _GEN_9645 : _GEN_7469; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9905 = _T_118 ? _GEN_9646 : _GEN_7470; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9906 = _T_118 ? _GEN_9647 : _GEN_7471; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9907 = _T_118 ? _GEN_9648 : _GEN_7472; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9908 = _T_118 ? _GEN_9649 : _GEN_7473; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9909 = _T_118 ? _GEN_9650 : _GEN_7474; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9910 = _T_118 ? _GEN_9651 : _GEN_7475; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9911 = _T_118 ? _GEN_9652 : _GEN_7476; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9912 = _T_118 ? _GEN_9653 : _GEN_7477; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9913 = _T_118 ? _GEN_9654 : _GEN_7478; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9914 = _T_118 ? _GEN_9655 : _GEN_7479; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9915 = _T_118 ? _GEN_9656 : _GEN_7480; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9916 = _T_118 ? _GEN_9657 : _GEN_7481; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9917 = _T_118 ? _GEN_9658 : _GEN_7482; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9918 = _T_118 ? _GEN_9659 : _GEN_7483; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9919 = _T_118 ? _GEN_9660 : _GEN_7484; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9920 = _T_118 ? _GEN_9661 : _GEN_7485; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9921 = _T_118 ? _GEN_9662 : _GEN_7486; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9922 = _T_118 ? _GEN_9663 : _GEN_7487; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9923 = _T_118 ? _GEN_9664 : _GEN_7488; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9924 = _T_118 ? _GEN_9665 : _GEN_7489; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9925 = _T_118 ? _GEN_9666 : _GEN_7490; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9926 = _T_118 ? _GEN_9667 : _GEN_7491; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9927 = _T_118 ? _GEN_9668 : _GEN_7492; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9928 = _T_118 ? _GEN_9669 : _GEN_7493; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9929 = _T_118 ? _GEN_9670 : _GEN_7494; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9930 = _T_118 ? _GEN_9671 : _GEN_7495; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9931 = _T_118 ? _GEN_9672 : _GEN_7496; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9932 = _T_118 ? _GEN_9673 : _GEN_7497; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9933 = _T_118 ? _GEN_9674 : _GEN_7498; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9934 = _T_118 ? _GEN_9675 : _GEN_7499; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9935 = _T_118 ? _GEN_9676 : _GEN_7500; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9936 = _T_118 ? _GEN_9677 : _GEN_7501; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9937 = _T_118 ? _GEN_9678 : _GEN_7502; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9938 = _T_118 ? _GEN_9679 : _GEN_7503; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9939 = _T_118 ? _GEN_9680 : _GEN_7504; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9940 = _T_118 ? _GEN_9681 : _GEN_7505; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9941 = _T_118 ? _GEN_9682 : _GEN_7506; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9942 = _T_118 ? _GEN_9683 : _GEN_7507; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9943 = _T_118 ? _GEN_9684 : _GEN_7508; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9944 = _T_118 ? _GEN_9685 : _GEN_7509; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9945 = _T_118 ? _GEN_9686 : _GEN_7510; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9946 = _T_118 ? _GEN_9687 : _GEN_7511; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9947 = _T_118 ? _GEN_9688 : _GEN_7512; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9948 = _T_118 ? _GEN_9689 : _GEN_7513; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9949 = _T_118 ? _GEN_9690 : _GEN_7514; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9950 = _T_118 ? _GEN_9691 : _GEN_7515; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9951 = _T_118 ? _GEN_9692 : _GEN_7516; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9952 = _T_118 ? _GEN_9693 : _GEN_7517; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9953 = _T_118 ? _GEN_9694 : _GEN_7518; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9954 = _T_118 ? _GEN_9695 : _GEN_7519; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9955 = _T_118 ? _GEN_9696 : _GEN_7520; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9956 = _T_118 ? _GEN_9697 : _GEN_7521; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9957 = _T_118 ? _GEN_9698 : _GEN_7522; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9958 = _T_118 ? _GEN_9699 : _GEN_7523; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9959 = _T_118 ? _GEN_9700 : _GEN_7524; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9960 = _T_118 ? _GEN_9701 : _GEN_7525; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9961 = _T_118 ? _GEN_9702 : _GEN_7526; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9962 = _T_118 ? _GEN_9703 : _GEN_7527; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9963 = _T_118 ? _GEN_9704 : _GEN_7528; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9964 = _T_118 ? _GEN_9705 : _GEN_7529; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9965 = _T_118 ? _GEN_9706 : _GEN_7530; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9966 = _T_118 ? _GEN_9707 : _GEN_7531; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9967 = _T_118 ? _GEN_9708 : _GEN_7532; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9968 = _T_118 ? _GEN_9709 : _GEN_7533; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9969 = _T_118 ? _GEN_9710 : _GEN_7534; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9970 = _T_118 ? _GEN_9711 : _GEN_7535; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9971 = _T_118 ? _GEN_9712 : _GEN_7536; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9972 = _T_118 ? _GEN_9713 : _GEN_7537; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9973 = _T_118 ? _GEN_9714 : _GEN_7538; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9974 = _T_118 ? _GEN_9715 : _GEN_7539; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9975 = _T_118 ? _GEN_9716 : _GEN_7540; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9976 = _T_118 ? _GEN_9717 : _GEN_7541; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9977 = _T_118 ? _GEN_9718 : _GEN_7542; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9978 = _T_118 ? _GEN_9719 : _GEN_7543; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9979 = _T_118 ? _GEN_9720 : _GEN_7544; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9980 = _T_118 ? _GEN_9721 : _GEN_7545; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9981 = _T_118 ? _GEN_9722 : _GEN_7546; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9982 = _T_118 ? _GEN_9723 : _GEN_7547; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9983 = _T_118 ? _GEN_9724 : _GEN_7548; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9984 = _T_118 ? _GEN_9725 : _GEN_7549; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9985 = _T_118 ? _GEN_9726 : _GEN_7550; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9986 = _T_118 ? _GEN_9727 : _GEN_7551; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9987 = _T_118 ? _GEN_9728 : _GEN_7552; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_9989 = _T_118 ? _GEN_9730 : {{9'd0}, packet_rob_idx}; // @[TestHarness.scala 199:26 197:29]
  wire [31:0] out_payload_1_tsc = io_from_noc_1_flit_bits_payload[63:32]; // @[TestHarness.scala 194:51]
  reg  packet_valid_1; // @[TestHarness.scala 196:31]
  reg [6:0] packet_rob_idx_1; // @[TestHarness.scala 197:29]
  wire [127:0] _T_123 = rob_valids >> out_payload_1_rob_idx; // @[TestHarness.scala 201:24]
  wire [31:0] _GEN_9991 = 7'h1 == out_payload_1_rob_idx[6:0] ? rob_payload_1_tsc : rob_payload_0_tsc; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_9992 = 7'h2 == out_payload_1_rob_idx[6:0] ? rob_payload_2_tsc : _GEN_9991; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_9993 = 7'h3 == out_payload_1_rob_idx[6:0] ? rob_payload_3_tsc : _GEN_9992; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_9994 = 7'h4 == out_payload_1_rob_idx[6:0] ? rob_payload_4_tsc : _GEN_9993; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_9995 = 7'h5 == out_payload_1_rob_idx[6:0] ? rob_payload_5_tsc : _GEN_9994; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_9996 = 7'h6 == out_payload_1_rob_idx[6:0] ? rob_payload_6_tsc : _GEN_9995; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_9997 = 7'h7 == out_payload_1_rob_idx[6:0] ? rob_payload_7_tsc : _GEN_9996; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_9998 = 7'h8 == out_payload_1_rob_idx[6:0] ? rob_payload_8_tsc : _GEN_9997; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_9999 = 7'h9 == out_payload_1_rob_idx[6:0] ? rob_payload_9_tsc : _GEN_9998; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10000 = 7'ha == out_payload_1_rob_idx[6:0] ? rob_payload_10_tsc : _GEN_9999; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10001 = 7'hb == out_payload_1_rob_idx[6:0] ? rob_payload_11_tsc : _GEN_10000; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10002 = 7'hc == out_payload_1_rob_idx[6:0] ? rob_payload_12_tsc : _GEN_10001; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10003 = 7'hd == out_payload_1_rob_idx[6:0] ? rob_payload_13_tsc : _GEN_10002; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10004 = 7'he == out_payload_1_rob_idx[6:0] ? rob_payload_14_tsc : _GEN_10003; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10005 = 7'hf == out_payload_1_rob_idx[6:0] ? rob_payload_15_tsc : _GEN_10004; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10006 = 7'h10 == out_payload_1_rob_idx[6:0] ? rob_payload_16_tsc : _GEN_10005; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10007 = 7'h11 == out_payload_1_rob_idx[6:0] ? rob_payload_17_tsc : _GEN_10006; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10008 = 7'h12 == out_payload_1_rob_idx[6:0] ? rob_payload_18_tsc : _GEN_10007; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10009 = 7'h13 == out_payload_1_rob_idx[6:0] ? rob_payload_19_tsc : _GEN_10008; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10010 = 7'h14 == out_payload_1_rob_idx[6:0] ? rob_payload_20_tsc : _GEN_10009; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10011 = 7'h15 == out_payload_1_rob_idx[6:0] ? rob_payload_21_tsc : _GEN_10010; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10012 = 7'h16 == out_payload_1_rob_idx[6:0] ? rob_payload_22_tsc : _GEN_10011; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10013 = 7'h17 == out_payload_1_rob_idx[6:0] ? rob_payload_23_tsc : _GEN_10012; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10014 = 7'h18 == out_payload_1_rob_idx[6:0] ? rob_payload_24_tsc : _GEN_10013; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10015 = 7'h19 == out_payload_1_rob_idx[6:0] ? rob_payload_25_tsc : _GEN_10014; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10016 = 7'h1a == out_payload_1_rob_idx[6:0] ? rob_payload_26_tsc : _GEN_10015; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10017 = 7'h1b == out_payload_1_rob_idx[6:0] ? rob_payload_27_tsc : _GEN_10016; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10018 = 7'h1c == out_payload_1_rob_idx[6:0] ? rob_payload_28_tsc : _GEN_10017; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10019 = 7'h1d == out_payload_1_rob_idx[6:0] ? rob_payload_29_tsc : _GEN_10018; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10020 = 7'h1e == out_payload_1_rob_idx[6:0] ? rob_payload_30_tsc : _GEN_10019; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10021 = 7'h1f == out_payload_1_rob_idx[6:0] ? rob_payload_31_tsc : _GEN_10020; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10022 = 7'h20 == out_payload_1_rob_idx[6:0] ? rob_payload_32_tsc : _GEN_10021; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10023 = 7'h21 == out_payload_1_rob_idx[6:0] ? rob_payload_33_tsc : _GEN_10022; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10024 = 7'h22 == out_payload_1_rob_idx[6:0] ? rob_payload_34_tsc : _GEN_10023; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10025 = 7'h23 == out_payload_1_rob_idx[6:0] ? rob_payload_35_tsc : _GEN_10024; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10026 = 7'h24 == out_payload_1_rob_idx[6:0] ? rob_payload_36_tsc : _GEN_10025; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10027 = 7'h25 == out_payload_1_rob_idx[6:0] ? rob_payload_37_tsc : _GEN_10026; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10028 = 7'h26 == out_payload_1_rob_idx[6:0] ? rob_payload_38_tsc : _GEN_10027; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10029 = 7'h27 == out_payload_1_rob_idx[6:0] ? rob_payload_39_tsc : _GEN_10028; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10030 = 7'h28 == out_payload_1_rob_idx[6:0] ? rob_payload_40_tsc : _GEN_10029; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10031 = 7'h29 == out_payload_1_rob_idx[6:0] ? rob_payload_41_tsc : _GEN_10030; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10032 = 7'h2a == out_payload_1_rob_idx[6:0] ? rob_payload_42_tsc : _GEN_10031; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10033 = 7'h2b == out_payload_1_rob_idx[6:0] ? rob_payload_43_tsc : _GEN_10032; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10034 = 7'h2c == out_payload_1_rob_idx[6:0] ? rob_payload_44_tsc : _GEN_10033; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10035 = 7'h2d == out_payload_1_rob_idx[6:0] ? rob_payload_45_tsc : _GEN_10034; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10036 = 7'h2e == out_payload_1_rob_idx[6:0] ? rob_payload_46_tsc : _GEN_10035; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10037 = 7'h2f == out_payload_1_rob_idx[6:0] ? rob_payload_47_tsc : _GEN_10036; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10038 = 7'h30 == out_payload_1_rob_idx[6:0] ? rob_payload_48_tsc : _GEN_10037; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10039 = 7'h31 == out_payload_1_rob_idx[6:0] ? rob_payload_49_tsc : _GEN_10038; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10040 = 7'h32 == out_payload_1_rob_idx[6:0] ? rob_payload_50_tsc : _GEN_10039; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10041 = 7'h33 == out_payload_1_rob_idx[6:0] ? rob_payload_51_tsc : _GEN_10040; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10042 = 7'h34 == out_payload_1_rob_idx[6:0] ? rob_payload_52_tsc : _GEN_10041; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10043 = 7'h35 == out_payload_1_rob_idx[6:0] ? rob_payload_53_tsc : _GEN_10042; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10044 = 7'h36 == out_payload_1_rob_idx[6:0] ? rob_payload_54_tsc : _GEN_10043; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10045 = 7'h37 == out_payload_1_rob_idx[6:0] ? rob_payload_55_tsc : _GEN_10044; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10046 = 7'h38 == out_payload_1_rob_idx[6:0] ? rob_payload_56_tsc : _GEN_10045; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10047 = 7'h39 == out_payload_1_rob_idx[6:0] ? rob_payload_57_tsc : _GEN_10046; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10048 = 7'h3a == out_payload_1_rob_idx[6:0] ? rob_payload_58_tsc : _GEN_10047; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10049 = 7'h3b == out_payload_1_rob_idx[6:0] ? rob_payload_59_tsc : _GEN_10048; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10050 = 7'h3c == out_payload_1_rob_idx[6:0] ? rob_payload_60_tsc : _GEN_10049; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10051 = 7'h3d == out_payload_1_rob_idx[6:0] ? rob_payload_61_tsc : _GEN_10050; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10052 = 7'h3e == out_payload_1_rob_idx[6:0] ? rob_payload_62_tsc : _GEN_10051; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10053 = 7'h3f == out_payload_1_rob_idx[6:0] ? rob_payload_63_tsc : _GEN_10052; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10054 = 7'h40 == out_payload_1_rob_idx[6:0] ? rob_payload_64_tsc : _GEN_10053; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10055 = 7'h41 == out_payload_1_rob_idx[6:0] ? rob_payload_65_tsc : _GEN_10054; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10056 = 7'h42 == out_payload_1_rob_idx[6:0] ? rob_payload_66_tsc : _GEN_10055; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10057 = 7'h43 == out_payload_1_rob_idx[6:0] ? rob_payload_67_tsc : _GEN_10056; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10058 = 7'h44 == out_payload_1_rob_idx[6:0] ? rob_payload_68_tsc : _GEN_10057; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10059 = 7'h45 == out_payload_1_rob_idx[6:0] ? rob_payload_69_tsc : _GEN_10058; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10060 = 7'h46 == out_payload_1_rob_idx[6:0] ? rob_payload_70_tsc : _GEN_10059; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10061 = 7'h47 == out_payload_1_rob_idx[6:0] ? rob_payload_71_tsc : _GEN_10060; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10062 = 7'h48 == out_payload_1_rob_idx[6:0] ? rob_payload_72_tsc : _GEN_10061; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10063 = 7'h49 == out_payload_1_rob_idx[6:0] ? rob_payload_73_tsc : _GEN_10062; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10064 = 7'h4a == out_payload_1_rob_idx[6:0] ? rob_payload_74_tsc : _GEN_10063; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10065 = 7'h4b == out_payload_1_rob_idx[6:0] ? rob_payload_75_tsc : _GEN_10064; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10066 = 7'h4c == out_payload_1_rob_idx[6:0] ? rob_payload_76_tsc : _GEN_10065; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10067 = 7'h4d == out_payload_1_rob_idx[6:0] ? rob_payload_77_tsc : _GEN_10066; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10068 = 7'h4e == out_payload_1_rob_idx[6:0] ? rob_payload_78_tsc : _GEN_10067; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10069 = 7'h4f == out_payload_1_rob_idx[6:0] ? rob_payload_79_tsc : _GEN_10068; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10070 = 7'h50 == out_payload_1_rob_idx[6:0] ? rob_payload_80_tsc : _GEN_10069; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10071 = 7'h51 == out_payload_1_rob_idx[6:0] ? rob_payload_81_tsc : _GEN_10070; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10072 = 7'h52 == out_payload_1_rob_idx[6:0] ? rob_payload_82_tsc : _GEN_10071; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10073 = 7'h53 == out_payload_1_rob_idx[6:0] ? rob_payload_83_tsc : _GEN_10072; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10074 = 7'h54 == out_payload_1_rob_idx[6:0] ? rob_payload_84_tsc : _GEN_10073; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10075 = 7'h55 == out_payload_1_rob_idx[6:0] ? rob_payload_85_tsc : _GEN_10074; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10076 = 7'h56 == out_payload_1_rob_idx[6:0] ? rob_payload_86_tsc : _GEN_10075; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10077 = 7'h57 == out_payload_1_rob_idx[6:0] ? rob_payload_87_tsc : _GEN_10076; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10078 = 7'h58 == out_payload_1_rob_idx[6:0] ? rob_payload_88_tsc : _GEN_10077; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10079 = 7'h59 == out_payload_1_rob_idx[6:0] ? rob_payload_89_tsc : _GEN_10078; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10080 = 7'h5a == out_payload_1_rob_idx[6:0] ? rob_payload_90_tsc : _GEN_10079; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10081 = 7'h5b == out_payload_1_rob_idx[6:0] ? rob_payload_91_tsc : _GEN_10080; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10082 = 7'h5c == out_payload_1_rob_idx[6:0] ? rob_payload_92_tsc : _GEN_10081; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10083 = 7'h5d == out_payload_1_rob_idx[6:0] ? rob_payload_93_tsc : _GEN_10082; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10084 = 7'h5e == out_payload_1_rob_idx[6:0] ? rob_payload_94_tsc : _GEN_10083; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10085 = 7'h5f == out_payload_1_rob_idx[6:0] ? rob_payload_95_tsc : _GEN_10084; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10086 = 7'h60 == out_payload_1_rob_idx[6:0] ? rob_payload_96_tsc : _GEN_10085; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10087 = 7'h61 == out_payload_1_rob_idx[6:0] ? rob_payload_97_tsc : _GEN_10086; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10088 = 7'h62 == out_payload_1_rob_idx[6:0] ? rob_payload_98_tsc : _GEN_10087; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10089 = 7'h63 == out_payload_1_rob_idx[6:0] ? rob_payload_99_tsc : _GEN_10088; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10090 = 7'h64 == out_payload_1_rob_idx[6:0] ? rob_payload_100_tsc : _GEN_10089; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10091 = 7'h65 == out_payload_1_rob_idx[6:0] ? rob_payload_101_tsc : _GEN_10090; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10092 = 7'h66 == out_payload_1_rob_idx[6:0] ? rob_payload_102_tsc : _GEN_10091; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10093 = 7'h67 == out_payload_1_rob_idx[6:0] ? rob_payload_103_tsc : _GEN_10092; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10094 = 7'h68 == out_payload_1_rob_idx[6:0] ? rob_payload_104_tsc : _GEN_10093; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10095 = 7'h69 == out_payload_1_rob_idx[6:0] ? rob_payload_105_tsc : _GEN_10094; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10096 = 7'h6a == out_payload_1_rob_idx[6:0] ? rob_payload_106_tsc : _GEN_10095; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10097 = 7'h6b == out_payload_1_rob_idx[6:0] ? rob_payload_107_tsc : _GEN_10096; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10098 = 7'h6c == out_payload_1_rob_idx[6:0] ? rob_payload_108_tsc : _GEN_10097; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10099 = 7'h6d == out_payload_1_rob_idx[6:0] ? rob_payload_109_tsc : _GEN_10098; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10100 = 7'h6e == out_payload_1_rob_idx[6:0] ? rob_payload_110_tsc : _GEN_10099; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10101 = 7'h6f == out_payload_1_rob_idx[6:0] ? rob_payload_111_tsc : _GEN_10100; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10102 = 7'h70 == out_payload_1_rob_idx[6:0] ? rob_payload_112_tsc : _GEN_10101; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10103 = 7'h71 == out_payload_1_rob_idx[6:0] ? rob_payload_113_tsc : _GEN_10102; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10104 = 7'h72 == out_payload_1_rob_idx[6:0] ? rob_payload_114_tsc : _GEN_10103; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10105 = 7'h73 == out_payload_1_rob_idx[6:0] ? rob_payload_115_tsc : _GEN_10104; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10106 = 7'h74 == out_payload_1_rob_idx[6:0] ? rob_payload_116_tsc : _GEN_10105; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10107 = 7'h75 == out_payload_1_rob_idx[6:0] ? rob_payload_117_tsc : _GEN_10106; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10108 = 7'h76 == out_payload_1_rob_idx[6:0] ? rob_payload_118_tsc : _GEN_10107; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10109 = 7'h77 == out_payload_1_rob_idx[6:0] ? rob_payload_119_tsc : _GEN_10108; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10110 = 7'h78 == out_payload_1_rob_idx[6:0] ? rob_payload_120_tsc : _GEN_10109; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10111 = 7'h79 == out_payload_1_rob_idx[6:0] ? rob_payload_121_tsc : _GEN_10110; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10112 = 7'h7a == out_payload_1_rob_idx[6:0] ? rob_payload_122_tsc : _GEN_10111; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10113 = 7'h7b == out_payload_1_rob_idx[6:0] ? rob_payload_123_tsc : _GEN_10112; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10114 = 7'h7c == out_payload_1_rob_idx[6:0] ? rob_payload_124_tsc : _GEN_10113; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10115 = 7'h7d == out_payload_1_rob_idx[6:0] ? rob_payload_125_tsc : _GEN_10114; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10116 = 7'h7e == out_payload_1_rob_idx[6:0] ? rob_payload_126_tsc : _GEN_10115; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_10117 = 7'h7f == out_payload_1_rob_idx[6:0] ? rob_payload_127_tsc : _GEN_10116; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10119 = 7'h1 == out_payload_1_rob_idx[6:0] ? rob_payload_1_rob_idx : rob_payload_0_rob_idx; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10120 = 7'h2 == out_payload_1_rob_idx[6:0] ? rob_payload_2_rob_idx : _GEN_10119; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10121 = 7'h3 == out_payload_1_rob_idx[6:0] ? rob_payload_3_rob_idx : _GEN_10120; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10122 = 7'h4 == out_payload_1_rob_idx[6:0] ? rob_payload_4_rob_idx : _GEN_10121; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10123 = 7'h5 == out_payload_1_rob_idx[6:0] ? rob_payload_5_rob_idx : _GEN_10122; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10124 = 7'h6 == out_payload_1_rob_idx[6:0] ? rob_payload_6_rob_idx : _GEN_10123; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10125 = 7'h7 == out_payload_1_rob_idx[6:0] ? rob_payload_7_rob_idx : _GEN_10124; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10126 = 7'h8 == out_payload_1_rob_idx[6:0] ? rob_payload_8_rob_idx : _GEN_10125; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10127 = 7'h9 == out_payload_1_rob_idx[6:0] ? rob_payload_9_rob_idx : _GEN_10126; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10128 = 7'ha == out_payload_1_rob_idx[6:0] ? rob_payload_10_rob_idx : _GEN_10127; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10129 = 7'hb == out_payload_1_rob_idx[6:0] ? rob_payload_11_rob_idx : _GEN_10128; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10130 = 7'hc == out_payload_1_rob_idx[6:0] ? rob_payload_12_rob_idx : _GEN_10129; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10131 = 7'hd == out_payload_1_rob_idx[6:0] ? rob_payload_13_rob_idx : _GEN_10130; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10132 = 7'he == out_payload_1_rob_idx[6:0] ? rob_payload_14_rob_idx : _GEN_10131; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10133 = 7'hf == out_payload_1_rob_idx[6:0] ? rob_payload_15_rob_idx : _GEN_10132; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10134 = 7'h10 == out_payload_1_rob_idx[6:0] ? rob_payload_16_rob_idx : _GEN_10133; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10135 = 7'h11 == out_payload_1_rob_idx[6:0] ? rob_payload_17_rob_idx : _GEN_10134; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10136 = 7'h12 == out_payload_1_rob_idx[6:0] ? rob_payload_18_rob_idx : _GEN_10135; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10137 = 7'h13 == out_payload_1_rob_idx[6:0] ? rob_payload_19_rob_idx : _GEN_10136; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10138 = 7'h14 == out_payload_1_rob_idx[6:0] ? rob_payload_20_rob_idx : _GEN_10137; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10139 = 7'h15 == out_payload_1_rob_idx[6:0] ? rob_payload_21_rob_idx : _GEN_10138; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10140 = 7'h16 == out_payload_1_rob_idx[6:0] ? rob_payload_22_rob_idx : _GEN_10139; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10141 = 7'h17 == out_payload_1_rob_idx[6:0] ? rob_payload_23_rob_idx : _GEN_10140; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10142 = 7'h18 == out_payload_1_rob_idx[6:0] ? rob_payload_24_rob_idx : _GEN_10141; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10143 = 7'h19 == out_payload_1_rob_idx[6:0] ? rob_payload_25_rob_idx : _GEN_10142; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10144 = 7'h1a == out_payload_1_rob_idx[6:0] ? rob_payload_26_rob_idx : _GEN_10143; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10145 = 7'h1b == out_payload_1_rob_idx[6:0] ? rob_payload_27_rob_idx : _GEN_10144; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10146 = 7'h1c == out_payload_1_rob_idx[6:0] ? rob_payload_28_rob_idx : _GEN_10145; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10147 = 7'h1d == out_payload_1_rob_idx[6:0] ? rob_payload_29_rob_idx : _GEN_10146; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10148 = 7'h1e == out_payload_1_rob_idx[6:0] ? rob_payload_30_rob_idx : _GEN_10147; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10149 = 7'h1f == out_payload_1_rob_idx[6:0] ? rob_payload_31_rob_idx : _GEN_10148; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10150 = 7'h20 == out_payload_1_rob_idx[6:0] ? rob_payload_32_rob_idx : _GEN_10149; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10151 = 7'h21 == out_payload_1_rob_idx[6:0] ? rob_payload_33_rob_idx : _GEN_10150; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10152 = 7'h22 == out_payload_1_rob_idx[6:0] ? rob_payload_34_rob_idx : _GEN_10151; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10153 = 7'h23 == out_payload_1_rob_idx[6:0] ? rob_payload_35_rob_idx : _GEN_10152; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10154 = 7'h24 == out_payload_1_rob_idx[6:0] ? rob_payload_36_rob_idx : _GEN_10153; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10155 = 7'h25 == out_payload_1_rob_idx[6:0] ? rob_payload_37_rob_idx : _GEN_10154; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10156 = 7'h26 == out_payload_1_rob_idx[6:0] ? rob_payload_38_rob_idx : _GEN_10155; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10157 = 7'h27 == out_payload_1_rob_idx[6:0] ? rob_payload_39_rob_idx : _GEN_10156; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10158 = 7'h28 == out_payload_1_rob_idx[6:0] ? rob_payload_40_rob_idx : _GEN_10157; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10159 = 7'h29 == out_payload_1_rob_idx[6:0] ? rob_payload_41_rob_idx : _GEN_10158; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10160 = 7'h2a == out_payload_1_rob_idx[6:0] ? rob_payload_42_rob_idx : _GEN_10159; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10161 = 7'h2b == out_payload_1_rob_idx[6:0] ? rob_payload_43_rob_idx : _GEN_10160; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10162 = 7'h2c == out_payload_1_rob_idx[6:0] ? rob_payload_44_rob_idx : _GEN_10161; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10163 = 7'h2d == out_payload_1_rob_idx[6:0] ? rob_payload_45_rob_idx : _GEN_10162; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10164 = 7'h2e == out_payload_1_rob_idx[6:0] ? rob_payload_46_rob_idx : _GEN_10163; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10165 = 7'h2f == out_payload_1_rob_idx[6:0] ? rob_payload_47_rob_idx : _GEN_10164; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10166 = 7'h30 == out_payload_1_rob_idx[6:0] ? rob_payload_48_rob_idx : _GEN_10165; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10167 = 7'h31 == out_payload_1_rob_idx[6:0] ? rob_payload_49_rob_idx : _GEN_10166; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10168 = 7'h32 == out_payload_1_rob_idx[6:0] ? rob_payload_50_rob_idx : _GEN_10167; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10169 = 7'h33 == out_payload_1_rob_idx[6:0] ? rob_payload_51_rob_idx : _GEN_10168; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10170 = 7'h34 == out_payload_1_rob_idx[6:0] ? rob_payload_52_rob_idx : _GEN_10169; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10171 = 7'h35 == out_payload_1_rob_idx[6:0] ? rob_payload_53_rob_idx : _GEN_10170; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10172 = 7'h36 == out_payload_1_rob_idx[6:0] ? rob_payload_54_rob_idx : _GEN_10171; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10173 = 7'h37 == out_payload_1_rob_idx[6:0] ? rob_payload_55_rob_idx : _GEN_10172; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10174 = 7'h38 == out_payload_1_rob_idx[6:0] ? rob_payload_56_rob_idx : _GEN_10173; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10175 = 7'h39 == out_payload_1_rob_idx[6:0] ? rob_payload_57_rob_idx : _GEN_10174; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10176 = 7'h3a == out_payload_1_rob_idx[6:0] ? rob_payload_58_rob_idx : _GEN_10175; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10177 = 7'h3b == out_payload_1_rob_idx[6:0] ? rob_payload_59_rob_idx : _GEN_10176; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10178 = 7'h3c == out_payload_1_rob_idx[6:0] ? rob_payload_60_rob_idx : _GEN_10177; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10179 = 7'h3d == out_payload_1_rob_idx[6:0] ? rob_payload_61_rob_idx : _GEN_10178; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10180 = 7'h3e == out_payload_1_rob_idx[6:0] ? rob_payload_62_rob_idx : _GEN_10179; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10181 = 7'h3f == out_payload_1_rob_idx[6:0] ? rob_payload_63_rob_idx : _GEN_10180; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10182 = 7'h40 == out_payload_1_rob_idx[6:0] ? rob_payload_64_rob_idx : _GEN_10181; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10183 = 7'h41 == out_payload_1_rob_idx[6:0] ? rob_payload_65_rob_idx : _GEN_10182; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10184 = 7'h42 == out_payload_1_rob_idx[6:0] ? rob_payload_66_rob_idx : _GEN_10183; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10185 = 7'h43 == out_payload_1_rob_idx[6:0] ? rob_payload_67_rob_idx : _GEN_10184; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10186 = 7'h44 == out_payload_1_rob_idx[6:0] ? rob_payload_68_rob_idx : _GEN_10185; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10187 = 7'h45 == out_payload_1_rob_idx[6:0] ? rob_payload_69_rob_idx : _GEN_10186; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10188 = 7'h46 == out_payload_1_rob_idx[6:0] ? rob_payload_70_rob_idx : _GEN_10187; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10189 = 7'h47 == out_payload_1_rob_idx[6:0] ? rob_payload_71_rob_idx : _GEN_10188; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10190 = 7'h48 == out_payload_1_rob_idx[6:0] ? rob_payload_72_rob_idx : _GEN_10189; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10191 = 7'h49 == out_payload_1_rob_idx[6:0] ? rob_payload_73_rob_idx : _GEN_10190; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10192 = 7'h4a == out_payload_1_rob_idx[6:0] ? rob_payload_74_rob_idx : _GEN_10191; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10193 = 7'h4b == out_payload_1_rob_idx[6:0] ? rob_payload_75_rob_idx : _GEN_10192; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10194 = 7'h4c == out_payload_1_rob_idx[6:0] ? rob_payload_76_rob_idx : _GEN_10193; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10195 = 7'h4d == out_payload_1_rob_idx[6:0] ? rob_payload_77_rob_idx : _GEN_10194; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10196 = 7'h4e == out_payload_1_rob_idx[6:0] ? rob_payload_78_rob_idx : _GEN_10195; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10197 = 7'h4f == out_payload_1_rob_idx[6:0] ? rob_payload_79_rob_idx : _GEN_10196; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10198 = 7'h50 == out_payload_1_rob_idx[6:0] ? rob_payload_80_rob_idx : _GEN_10197; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10199 = 7'h51 == out_payload_1_rob_idx[6:0] ? rob_payload_81_rob_idx : _GEN_10198; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10200 = 7'h52 == out_payload_1_rob_idx[6:0] ? rob_payload_82_rob_idx : _GEN_10199; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10201 = 7'h53 == out_payload_1_rob_idx[6:0] ? rob_payload_83_rob_idx : _GEN_10200; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10202 = 7'h54 == out_payload_1_rob_idx[6:0] ? rob_payload_84_rob_idx : _GEN_10201; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10203 = 7'h55 == out_payload_1_rob_idx[6:0] ? rob_payload_85_rob_idx : _GEN_10202; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10204 = 7'h56 == out_payload_1_rob_idx[6:0] ? rob_payload_86_rob_idx : _GEN_10203; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10205 = 7'h57 == out_payload_1_rob_idx[6:0] ? rob_payload_87_rob_idx : _GEN_10204; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10206 = 7'h58 == out_payload_1_rob_idx[6:0] ? rob_payload_88_rob_idx : _GEN_10205; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10207 = 7'h59 == out_payload_1_rob_idx[6:0] ? rob_payload_89_rob_idx : _GEN_10206; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10208 = 7'h5a == out_payload_1_rob_idx[6:0] ? rob_payload_90_rob_idx : _GEN_10207; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10209 = 7'h5b == out_payload_1_rob_idx[6:0] ? rob_payload_91_rob_idx : _GEN_10208; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10210 = 7'h5c == out_payload_1_rob_idx[6:0] ? rob_payload_92_rob_idx : _GEN_10209; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10211 = 7'h5d == out_payload_1_rob_idx[6:0] ? rob_payload_93_rob_idx : _GEN_10210; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10212 = 7'h5e == out_payload_1_rob_idx[6:0] ? rob_payload_94_rob_idx : _GEN_10211; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10213 = 7'h5f == out_payload_1_rob_idx[6:0] ? rob_payload_95_rob_idx : _GEN_10212; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10214 = 7'h60 == out_payload_1_rob_idx[6:0] ? rob_payload_96_rob_idx : _GEN_10213; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10215 = 7'h61 == out_payload_1_rob_idx[6:0] ? rob_payload_97_rob_idx : _GEN_10214; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10216 = 7'h62 == out_payload_1_rob_idx[6:0] ? rob_payload_98_rob_idx : _GEN_10215; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10217 = 7'h63 == out_payload_1_rob_idx[6:0] ? rob_payload_99_rob_idx : _GEN_10216; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10218 = 7'h64 == out_payload_1_rob_idx[6:0] ? rob_payload_100_rob_idx : _GEN_10217; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10219 = 7'h65 == out_payload_1_rob_idx[6:0] ? rob_payload_101_rob_idx : _GEN_10218; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10220 = 7'h66 == out_payload_1_rob_idx[6:0] ? rob_payload_102_rob_idx : _GEN_10219; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10221 = 7'h67 == out_payload_1_rob_idx[6:0] ? rob_payload_103_rob_idx : _GEN_10220; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10222 = 7'h68 == out_payload_1_rob_idx[6:0] ? rob_payload_104_rob_idx : _GEN_10221; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10223 = 7'h69 == out_payload_1_rob_idx[6:0] ? rob_payload_105_rob_idx : _GEN_10222; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10224 = 7'h6a == out_payload_1_rob_idx[6:0] ? rob_payload_106_rob_idx : _GEN_10223; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10225 = 7'h6b == out_payload_1_rob_idx[6:0] ? rob_payload_107_rob_idx : _GEN_10224; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10226 = 7'h6c == out_payload_1_rob_idx[6:0] ? rob_payload_108_rob_idx : _GEN_10225; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10227 = 7'h6d == out_payload_1_rob_idx[6:0] ? rob_payload_109_rob_idx : _GEN_10226; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10228 = 7'h6e == out_payload_1_rob_idx[6:0] ? rob_payload_110_rob_idx : _GEN_10227; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10229 = 7'h6f == out_payload_1_rob_idx[6:0] ? rob_payload_111_rob_idx : _GEN_10228; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10230 = 7'h70 == out_payload_1_rob_idx[6:0] ? rob_payload_112_rob_idx : _GEN_10229; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10231 = 7'h71 == out_payload_1_rob_idx[6:0] ? rob_payload_113_rob_idx : _GEN_10230; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10232 = 7'h72 == out_payload_1_rob_idx[6:0] ? rob_payload_114_rob_idx : _GEN_10231; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10233 = 7'h73 == out_payload_1_rob_idx[6:0] ? rob_payload_115_rob_idx : _GEN_10232; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10234 = 7'h74 == out_payload_1_rob_idx[6:0] ? rob_payload_116_rob_idx : _GEN_10233; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10235 = 7'h75 == out_payload_1_rob_idx[6:0] ? rob_payload_117_rob_idx : _GEN_10234; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10236 = 7'h76 == out_payload_1_rob_idx[6:0] ? rob_payload_118_rob_idx : _GEN_10235; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10237 = 7'h77 == out_payload_1_rob_idx[6:0] ? rob_payload_119_rob_idx : _GEN_10236; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10238 = 7'h78 == out_payload_1_rob_idx[6:0] ? rob_payload_120_rob_idx : _GEN_10237; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10239 = 7'h79 == out_payload_1_rob_idx[6:0] ? rob_payload_121_rob_idx : _GEN_10238; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10240 = 7'h7a == out_payload_1_rob_idx[6:0] ? rob_payload_122_rob_idx : _GEN_10239; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10241 = 7'h7b == out_payload_1_rob_idx[6:0] ? rob_payload_123_rob_idx : _GEN_10240; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10242 = 7'h7c == out_payload_1_rob_idx[6:0] ? rob_payload_124_rob_idx : _GEN_10241; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10243 = 7'h7d == out_payload_1_rob_idx[6:0] ? rob_payload_125_rob_idx : _GEN_10242; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10244 = 7'h7e == out_payload_1_rob_idx[6:0] ? rob_payload_126_rob_idx : _GEN_10243; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10245 = 7'h7f == out_payload_1_rob_idx[6:0] ? rob_payload_127_rob_idx : _GEN_10244; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10247 = 7'h1 == out_payload_1_rob_idx[6:0] ? rob_payload_1_flits_fired : rob_payload_0_flits_fired; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10248 = 7'h2 == out_payload_1_rob_idx[6:0] ? rob_payload_2_flits_fired : _GEN_10247; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10249 = 7'h3 == out_payload_1_rob_idx[6:0] ? rob_payload_3_flits_fired : _GEN_10248; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10250 = 7'h4 == out_payload_1_rob_idx[6:0] ? rob_payload_4_flits_fired : _GEN_10249; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10251 = 7'h5 == out_payload_1_rob_idx[6:0] ? rob_payload_5_flits_fired : _GEN_10250; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10252 = 7'h6 == out_payload_1_rob_idx[6:0] ? rob_payload_6_flits_fired : _GEN_10251; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10253 = 7'h7 == out_payload_1_rob_idx[6:0] ? rob_payload_7_flits_fired : _GEN_10252; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10254 = 7'h8 == out_payload_1_rob_idx[6:0] ? rob_payload_8_flits_fired : _GEN_10253; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10255 = 7'h9 == out_payload_1_rob_idx[6:0] ? rob_payload_9_flits_fired : _GEN_10254; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10256 = 7'ha == out_payload_1_rob_idx[6:0] ? rob_payload_10_flits_fired : _GEN_10255; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10257 = 7'hb == out_payload_1_rob_idx[6:0] ? rob_payload_11_flits_fired : _GEN_10256; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10258 = 7'hc == out_payload_1_rob_idx[6:0] ? rob_payload_12_flits_fired : _GEN_10257; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10259 = 7'hd == out_payload_1_rob_idx[6:0] ? rob_payload_13_flits_fired : _GEN_10258; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10260 = 7'he == out_payload_1_rob_idx[6:0] ? rob_payload_14_flits_fired : _GEN_10259; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10261 = 7'hf == out_payload_1_rob_idx[6:0] ? rob_payload_15_flits_fired : _GEN_10260; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10262 = 7'h10 == out_payload_1_rob_idx[6:0] ? rob_payload_16_flits_fired : _GEN_10261; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10263 = 7'h11 == out_payload_1_rob_idx[6:0] ? rob_payload_17_flits_fired : _GEN_10262; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10264 = 7'h12 == out_payload_1_rob_idx[6:0] ? rob_payload_18_flits_fired : _GEN_10263; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10265 = 7'h13 == out_payload_1_rob_idx[6:0] ? rob_payload_19_flits_fired : _GEN_10264; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10266 = 7'h14 == out_payload_1_rob_idx[6:0] ? rob_payload_20_flits_fired : _GEN_10265; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10267 = 7'h15 == out_payload_1_rob_idx[6:0] ? rob_payload_21_flits_fired : _GEN_10266; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10268 = 7'h16 == out_payload_1_rob_idx[6:0] ? rob_payload_22_flits_fired : _GEN_10267; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10269 = 7'h17 == out_payload_1_rob_idx[6:0] ? rob_payload_23_flits_fired : _GEN_10268; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10270 = 7'h18 == out_payload_1_rob_idx[6:0] ? rob_payload_24_flits_fired : _GEN_10269; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10271 = 7'h19 == out_payload_1_rob_idx[6:0] ? rob_payload_25_flits_fired : _GEN_10270; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10272 = 7'h1a == out_payload_1_rob_idx[6:0] ? rob_payload_26_flits_fired : _GEN_10271; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10273 = 7'h1b == out_payload_1_rob_idx[6:0] ? rob_payload_27_flits_fired : _GEN_10272; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10274 = 7'h1c == out_payload_1_rob_idx[6:0] ? rob_payload_28_flits_fired : _GEN_10273; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10275 = 7'h1d == out_payload_1_rob_idx[6:0] ? rob_payload_29_flits_fired : _GEN_10274; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10276 = 7'h1e == out_payload_1_rob_idx[6:0] ? rob_payload_30_flits_fired : _GEN_10275; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10277 = 7'h1f == out_payload_1_rob_idx[6:0] ? rob_payload_31_flits_fired : _GEN_10276; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10278 = 7'h20 == out_payload_1_rob_idx[6:0] ? rob_payload_32_flits_fired : _GEN_10277; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10279 = 7'h21 == out_payload_1_rob_idx[6:0] ? rob_payload_33_flits_fired : _GEN_10278; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10280 = 7'h22 == out_payload_1_rob_idx[6:0] ? rob_payload_34_flits_fired : _GEN_10279; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10281 = 7'h23 == out_payload_1_rob_idx[6:0] ? rob_payload_35_flits_fired : _GEN_10280; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10282 = 7'h24 == out_payload_1_rob_idx[6:0] ? rob_payload_36_flits_fired : _GEN_10281; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10283 = 7'h25 == out_payload_1_rob_idx[6:0] ? rob_payload_37_flits_fired : _GEN_10282; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10284 = 7'h26 == out_payload_1_rob_idx[6:0] ? rob_payload_38_flits_fired : _GEN_10283; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10285 = 7'h27 == out_payload_1_rob_idx[6:0] ? rob_payload_39_flits_fired : _GEN_10284; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10286 = 7'h28 == out_payload_1_rob_idx[6:0] ? rob_payload_40_flits_fired : _GEN_10285; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10287 = 7'h29 == out_payload_1_rob_idx[6:0] ? rob_payload_41_flits_fired : _GEN_10286; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10288 = 7'h2a == out_payload_1_rob_idx[6:0] ? rob_payload_42_flits_fired : _GEN_10287; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10289 = 7'h2b == out_payload_1_rob_idx[6:0] ? rob_payload_43_flits_fired : _GEN_10288; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10290 = 7'h2c == out_payload_1_rob_idx[6:0] ? rob_payload_44_flits_fired : _GEN_10289; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10291 = 7'h2d == out_payload_1_rob_idx[6:0] ? rob_payload_45_flits_fired : _GEN_10290; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10292 = 7'h2e == out_payload_1_rob_idx[6:0] ? rob_payload_46_flits_fired : _GEN_10291; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10293 = 7'h2f == out_payload_1_rob_idx[6:0] ? rob_payload_47_flits_fired : _GEN_10292; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10294 = 7'h30 == out_payload_1_rob_idx[6:0] ? rob_payload_48_flits_fired : _GEN_10293; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10295 = 7'h31 == out_payload_1_rob_idx[6:0] ? rob_payload_49_flits_fired : _GEN_10294; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10296 = 7'h32 == out_payload_1_rob_idx[6:0] ? rob_payload_50_flits_fired : _GEN_10295; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10297 = 7'h33 == out_payload_1_rob_idx[6:0] ? rob_payload_51_flits_fired : _GEN_10296; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10298 = 7'h34 == out_payload_1_rob_idx[6:0] ? rob_payload_52_flits_fired : _GEN_10297; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10299 = 7'h35 == out_payload_1_rob_idx[6:0] ? rob_payload_53_flits_fired : _GEN_10298; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10300 = 7'h36 == out_payload_1_rob_idx[6:0] ? rob_payload_54_flits_fired : _GEN_10299; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10301 = 7'h37 == out_payload_1_rob_idx[6:0] ? rob_payload_55_flits_fired : _GEN_10300; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10302 = 7'h38 == out_payload_1_rob_idx[6:0] ? rob_payload_56_flits_fired : _GEN_10301; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10303 = 7'h39 == out_payload_1_rob_idx[6:0] ? rob_payload_57_flits_fired : _GEN_10302; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10304 = 7'h3a == out_payload_1_rob_idx[6:0] ? rob_payload_58_flits_fired : _GEN_10303; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10305 = 7'h3b == out_payload_1_rob_idx[6:0] ? rob_payload_59_flits_fired : _GEN_10304; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10306 = 7'h3c == out_payload_1_rob_idx[6:0] ? rob_payload_60_flits_fired : _GEN_10305; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10307 = 7'h3d == out_payload_1_rob_idx[6:0] ? rob_payload_61_flits_fired : _GEN_10306; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10308 = 7'h3e == out_payload_1_rob_idx[6:0] ? rob_payload_62_flits_fired : _GEN_10307; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10309 = 7'h3f == out_payload_1_rob_idx[6:0] ? rob_payload_63_flits_fired : _GEN_10308; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10310 = 7'h40 == out_payload_1_rob_idx[6:0] ? rob_payload_64_flits_fired : _GEN_10309; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10311 = 7'h41 == out_payload_1_rob_idx[6:0] ? rob_payload_65_flits_fired : _GEN_10310; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10312 = 7'h42 == out_payload_1_rob_idx[6:0] ? rob_payload_66_flits_fired : _GEN_10311; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10313 = 7'h43 == out_payload_1_rob_idx[6:0] ? rob_payload_67_flits_fired : _GEN_10312; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10314 = 7'h44 == out_payload_1_rob_idx[6:0] ? rob_payload_68_flits_fired : _GEN_10313; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10315 = 7'h45 == out_payload_1_rob_idx[6:0] ? rob_payload_69_flits_fired : _GEN_10314; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10316 = 7'h46 == out_payload_1_rob_idx[6:0] ? rob_payload_70_flits_fired : _GEN_10315; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10317 = 7'h47 == out_payload_1_rob_idx[6:0] ? rob_payload_71_flits_fired : _GEN_10316; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10318 = 7'h48 == out_payload_1_rob_idx[6:0] ? rob_payload_72_flits_fired : _GEN_10317; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10319 = 7'h49 == out_payload_1_rob_idx[6:0] ? rob_payload_73_flits_fired : _GEN_10318; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10320 = 7'h4a == out_payload_1_rob_idx[6:0] ? rob_payload_74_flits_fired : _GEN_10319; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10321 = 7'h4b == out_payload_1_rob_idx[6:0] ? rob_payload_75_flits_fired : _GEN_10320; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10322 = 7'h4c == out_payload_1_rob_idx[6:0] ? rob_payload_76_flits_fired : _GEN_10321; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10323 = 7'h4d == out_payload_1_rob_idx[6:0] ? rob_payload_77_flits_fired : _GEN_10322; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10324 = 7'h4e == out_payload_1_rob_idx[6:0] ? rob_payload_78_flits_fired : _GEN_10323; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10325 = 7'h4f == out_payload_1_rob_idx[6:0] ? rob_payload_79_flits_fired : _GEN_10324; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10326 = 7'h50 == out_payload_1_rob_idx[6:0] ? rob_payload_80_flits_fired : _GEN_10325; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10327 = 7'h51 == out_payload_1_rob_idx[6:0] ? rob_payload_81_flits_fired : _GEN_10326; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10328 = 7'h52 == out_payload_1_rob_idx[6:0] ? rob_payload_82_flits_fired : _GEN_10327; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10329 = 7'h53 == out_payload_1_rob_idx[6:0] ? rob_payload_83_flits_fired : _GEN_10328; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10330 = 7'h54 == out_payload_1_rob_idx[6:0] ? rob_payload_84_flits_fired : _GEN_10329; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10331 = 7'h55 == out_payload_1_rob_idx[6:0] ? rob_payload_85_flits_fired : _GEN_10330; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10332 = 7'h56 == out_payload_1_rob_idx[6:0] ? rob_payload_86_flits_fired : _GEN_10331; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10333 = 7'h57 == out_payload_1_rob_idx[6:0] ? rob_payload_87_flits_fired : _GEN_10332; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10334 = 7'h58 == out_payload_1_rob_idx[6:0] ? rob_payload_88_flits_fired : _GEN_10333; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10335 = 7'h59 == out_payload_1_rob_idx[6:0] ? rob_payload_89_flits_fired : _GEN_10334; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10336 = 7'h5a == out_payload_1_rob_idx[6:0] ? rob_payload_90_flits_fired : _GEN_10335; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10337 = 7'h5b == out_payload_1_rob_idx[6:0] ? rob_payload_91_flits_fired : _GEN_10336; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10338 = 7'h5c == out_payload_1_rob_idx[6:0] ? rob_payload_92_flits_fired : _GEN_10337; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10339 = 7'h5d == out_payload_1_rob_idx[6:0] ? rob_payload_93_flits_fired : _GEN_10338; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10340 = 7'h5e == out_payload_1_rob_idx[6:0] ? rob_payload_94_flits_fired : _GEN_10339; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10341 = 7'h5f == out_payload_1_rob_idx[6:0] ? rob_payload_95_flits_fired : _GEN_10340; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10342 = 7'h60 == out_payload_1_rob_idx[6:0] ? rob_payload_96_flits_fired : _GEN_10341; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10343 = 7'h61 == out_payload_1_rob_idx[6:0] ? rob_payload_97_flits_fired : _GEN_10342; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10344 = 7'h62 == out_payload_1_rob_idx[6:0] ? rob_payload_98_flits_fired : _GEN_10343; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10345 = 7'h63 == out_payload_1_rob_idx[6:0] ? rob_payload_99_flits_fired : _GEN_10344; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10346 = 7'h64 == out_payload_1_rob_idx[6:0] ? rob_payload_100_flits_fired : _GEN_10345; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10347 = 7'h65 == out_payload_1_rob_idx[6:0] ? rob_payload_101_flits_fired : _GEN_10346; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10348 = 7'h66 == out_payload_1_rob_idx[6:0] ? rob_payload_102_flits_fired : _GEN_10347; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10349 = 7'h67 == out_payload_1_rob_idx[6:0] ? rob_payload_103_flits_fired : _GEN_10348; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10350 = 7'h68 == out_payload_1_rob_idx[6:0] ? rob_payload_104_flits_fired : _GEN_10349; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10351 = 7'h69 == out_payload_1_rob_idx[6:0] ? rob_payload_105_flits_fired : _GEN_10350; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10352 = 7'h6a == out_payload_1_rob_idx[6:0] ? rob_payload_106_flits_fired : _GEN_10351; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10353 = 7'h6b == out_payload_1_rob_idx[6:0] ? rob_payload_107_flits_fired : _GEN_10352; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10354 = 7'h6c == out_payload_1_rob_idx[6:0] ? rob_payload_108_flits_fired : _GEN_10353; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10355 = 7'h6d == out_payload_1_rob_idx[6:0] ? rob_payload_109_flits_fired : _GEN_10354; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10356 = 7'h6e == out_payload_1_rob_idx[6:0] ? rob_payload_110_flits_fired : _GEN_10355; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10357 = 7'h6f == out_payload_1_rob_idx[6:0] ? rob_payload_111_flits_fired : _GEN_10356; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10358 = 7'h70 == out_payload_1_rob_idx[6:0] ? rob_payload_112_flits_fired : _GEN_10357; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10359 = 7'h71 == out_payload_1_rob_idx[6:0] ? rob_payload_113_flits_fired : _GEN_10358; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10360 = 7'h72 == out_payload_1_rob_idx[6:0] ? rob_payload_114_flits_fired : _GEN_10359; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10361 = 7'h73 == out_payload_1_rob_idx[6:0] ? rob_payload_115_flits_fired : _GEN_10360; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10362 = 7'h74 == out_payload_1_rob_idx[6:0] ? rob_payload_116_flits_fired : _GEN_10361; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10363 = 7'h75 == out_payload_1_rob_idx[6:0] ? rob_payload_117_flits_fired : _GEN_10362; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10364 = 7'h76 == out_payload_1_rob_idx[6:0] ? rob_payload_118_flits_fired : _GEN_10363; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10365 = 7'h77 == out_payload_1_rob_idx[6:0] ? rob_payload_119_flits_fired : _GEN_10364; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10366 = 7'h78 == out_payload_1_rob_idx[6:0] ? rob_payload_120_flits_fired : _GEN_10365; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10367 = 7'h79 == out_payload_1_rob_idx[6:0] ? rob_payload_121_flits_fired : _GEN_10366; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10368 = 7'h7a == out_payload_1_rob_idx[6:0] ? rob_payload_122_flits_fired : _GEN_10367; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10369 = 7'h7b == out_payload_1_rob_idx[6:0] ? rob_payload_123_flits_fired : _GEN_10368; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10370 = 7'h7c == out_payload_1_rob_idx[6:0] ? rob_payload_124_flits_fired : _GEN_10369; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10371 = 7'h7d == out_payload_1_rob_idx[6:0] ? rob_payload_125_flits_fired : _GEN_10370; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10372 = 7'h7e == out_payload_1_rob_idx[6:0] ? rob_payload_126_flits_fired : _GEN_10371; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_10373 = 7'h7f == out_payload_1_rob_idx[6:0] ? rob_payload_127_flits_fired : _GEN_10372; // @[TestHarness.scala 202:{35,35}]
  wire [63:0] _T_129 = {_GEN_10117,_GEN_10245,_GEN_10373}; // @[TestHarness.scala 202:35]
  wire [1:0] _GEN_10375 = 7'h1 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_1 : rob_ingress_id_0; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10376 = 7'h2 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_2 : _GEN_10375; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10377 = 7'h3 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_3 : _GEN_10376; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10378 = 7'h4 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_4 : _GEN_10377; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10379 = 7'h5 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_5 : _GEN_10378; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10380 = 7'h6 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_6 : _GEN_10379; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10381 = 7'h7 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_7 : _GEN_10380; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10382 = 7'h8 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_8 : _GEN_10381; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10383 = 7'h9 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_9 : _GEN_10382; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10384 = 7'ha == out_payload_1_rob_idx[6:0] ? rob_ingress_id_10 : _GEN_10383; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10385 = 7'hb == out_payload_1_rob_idx[6:0] ? rob_ingress_id_11 : _GEN_10384; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10386 = 7'hc == out_payload_1_rob_idx[6:0] ? rob_ingress_id_12 : _GEN_10385; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10387 = 7'hd == out_payload_1_rob_idx[6:0] ? rob_ingress_id_13 : _GEN_10386; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10388 = 7'he == out_payload_1_rob_idx[6:0] ? rob_ingress_id_14 : _GEN_10387; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10389 = 7'hf == out_payload_1_rob_idx[6:0] ? rob_ingress_id_15 : _GEN_10388; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10390 = 7'h10 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_16 : _GEN_10389; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10391 = 7'h11 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_17 : _GEN_10390; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10392 = 7'h12 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_18 : _GEN_10391; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10393 = 7'h13 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_19 : _GEN_10392; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10394 = 7'h14 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_20 : _GEN_10393; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10395 = 7'h15 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_21 : _GEN_10394; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10396 = 7'h16 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_22 : _GEN_10395; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10397 = 7'h17 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_23 : _GEN_10396; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10398 = 7'h18 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_24 : _GEN_10397; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10399 = 7'h19 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_25 : _GEN_10398; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10400 = 7'h1a == out_payload_1_rob_idx[6:0] ? rob_ingress_id_26 : _GEN_10399; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10401 = 7'h1b == out_payload_1_rob_idx[6:0] ? rob_ingress_id_27 : _GEN_10400; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10402 = 7'h1c == out_payload_1_rob_idx[6:0] ? rob_ingress_id_28 : _GEN_10401; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10403 = 7'h1d == out_payload_1_rob_idx[6:0] ? rob_ingress_id_29 : _GEN_10402; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10404 = 7'h1e == out_payload_1_rob_idx[6:0] ? rob_ingress_id_30 : _GEN_10403; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10405 = 7'h1f == out_payload_1_rob_idx[6:0] ? rob_ingress_id_31 : _GEN_10404; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10406 = 7'h20 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_32 : _GEN_10405; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10407 = 7'h21 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_33 : _GEN_10406; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10408 = 7'h22 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_34 : _GEN_10407; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10409 = 7'h23 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_35 : _GEN_10408; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10410 = 7'h24 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_36 : _GEN_10409; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10411 = 7'h25 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_37 : _GEN_10410; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10412 = 7'h26 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_38 : _GEN_10411; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10413 = 7'h27 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_39 : _GEN_10412; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10414 = 7'h28 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_40 : _GEN_10413; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10415 = 7'h29 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_41 : _GEN_10414; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10416 = 7'h2a == out_payload_1_rob_idx[6:0] ? rob_ingress_id_42 : _GEN_10415; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10417 = 7'h2b == out_payload_1_rob_idx[6:0] ? rob_ingress_id_43 : _GEN_10416; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10418 = 7'h2c == out_payload_1_rob_idx[6:0] ? rob_ingress_id_44 : _GEN_10417; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10419 = 7'h2d == out_payload_1_rob_idx[6:0] ? rob_ingress_id_45 : _GEN_10418; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10420 = 7'h2e == out_payload_1_rob_idx[6:0] ? rob_ingress_id_46 : _GEN_10419; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10421 = 7'h2f == out_payload_1_rob_idx[6:0] ? rob_ingress_id_47 : _GEN_10420; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10422 = 7'h30 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_48 : _GEN_10421; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10423 = 7'h31 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_49 : _GEN_10422; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10424 = 7'h32 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_50 : _GEN_10423; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10425 = 7'h33 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_51 : _GEN_10424; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10426 = 7'h34 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_52 : _GEN_10425; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10427 = 7'h35 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_53 : _GEN_10426; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10428 = 7'h36 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_54 : _GEN_10427; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10429 = 7'h37 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_55 : _GEN_10428; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10430 = 7'h38 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_56 : _GEN_10429; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10431 = 7'h39 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_57 : _GEN_10430; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10432 = 7'h3a == out_payload_1_rob_idx[6:0] ? rob_ingress_id_58 : _GEN_10431; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10433 = 7'h3b == out_payload_1_rob_idx[6:0] ? rob_ingress_id_59 : _GEN_10432; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10434 = 7'h3c == out_payload_1_rob_idx[6:0] ? rob_ingress_id_60 : _GEN_10433; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10435 = 7'h3d == out_payload_1_rob_idx[6:0] ? rob_ingress_id_61 : _GEN_10434; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10436 = 7'h3e == out_payload_1_rob_idx[6:0] ? rob_ingress_id_62 : _GEN_10435; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10437 = 7'h3f == out_payload_1_rob_idx[6:0] ? rob_ingress_id_63 : _GEN_10436; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10438 = 7'h40 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_64 : _GEN_10437; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10439 = 7'h41 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_65 : _GEN_10438; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10440 = 7'h42 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_66 : _GEN_10439; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10441 = 7'h43 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_67 : _GEN_10440; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10442 = 7'h44 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_68 : _GEN_10441; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10443 = 7'h45 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_69 : _GEN_10442; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10444 = 7'h46 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_70 : _GEN_10443; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10445 = 7'h47 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_71 : _GEN_10444; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10446 = 7'h48 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_72 : _GEN_10445; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10447 = 7'h49 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_73 : _GEN_10446; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10448 = 7'h4a == out_payload_1_rob_idx[6:0] ? rob_ingress_id_74 : _GEN_10447; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10449 = 7'h4b == out_payload_1_rob_idx[6:0] ? rob_ingress_id_75 : _GEN_10448; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10450 = 7'h4c == out_payload_1_rob_idx[6:0] ? rob_ingress_id_76 : _GEN_10449; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10451 = 7'h4d == out_payload_1_rob_idx[6:0] ? rob_ingress_id_77 : _GEN_10450; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10452 = 7'h4e == out_payload_1_rob_idx[6:0] ? rob_ingress_id_78 : _GEN_10451; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10453 = 7'h4f == out_payload_1_rob_idx[6:0] ? rob_ingress_id_79 : _GEN_10452; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10454 = 7'h50 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_80 : _GEN_10453; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10455 = 7'h51 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_81 : _GEN_10454; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10456 = 7'h52 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_82 : _GEN_10455; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10457 = 7'h53 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_83 : _GEN_10456; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10458 = 7'h54 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_84 : _GEN_10457; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10459 = 7'h55 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_85 : _GEN_10458; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10460 = 7'h56 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_86 : _GEN_10459; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10461 = 7'h57 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_87 : _GEN_10460; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10462 = 7'h58 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_88 : _GEN_10461; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10463 = 7'h59 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_89 : _GEN_10462; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10464 = 7'h5a == out_payload_1_rob_idx[6:0] ? rob_ingress_id_90 : _GEN_10463; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10465 = 7'h5b == out_payload_1_rob_idx[6:0] ? rob_ingress_id_91 : _GEN_10464; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10466 = 7'h5c == out_payload_1_rob_idx[6:0] ? rob_ingress_id_92 : _GEN_10465; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10467 = 7'h5d == out_payload_1_rob_idx[6:0] ? rob_ingress_id_93 : _GEN_10466; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10468 = 7'h5e == out_payload_1_rob_idx[6:0] ? rob_ingress_id_94 : _GEN_10467; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10469 = 7'h5f == out_payload_1_rob_idx[6:0] ? rob_ingress_id_95 : _GEN_10468; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10470 = 7'h60 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_96 : _GEN_10469; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10471 = 7'h61 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_97 : _GEN_10470; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10472 = 7'h62 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_98 : _GEN_10471; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10473 = 7'h63 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_99 : _GEN_10472; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10474 = 7'h64 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_100 : _GEN_10473; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10475 = 7'h65 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_101 : _GEN_10474; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10476 = 7'h66 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_102 : _GEN_10475; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10477 = 7'h67 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_103 : _GEN_10476; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10478 = 7'h68 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_104 : _GEN_10477; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10479 = 7'h69 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_105 : _GEN_10478; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10480 = 7'h6a == out_payload_1_rob_idx[6:0] ? rob_ingress_id_106 : _GEN_10479; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10481 = 7'h6b == out_payload_1_rob_idx[6:0] ? rob_ingress_id_107 : _GEN_10480; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10482 = 7'h6c == out_payload_1_rob_idx[6:0] ? rob_ingress_id_108 : _GEN_10481; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10483 = 7'h6d == out_payload_1_rob_idx[6:0] ? rob_ingress_id_109 : _GEN_10482; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10484 = 7'h6e == out_payload_1_rob_idx[6:0] ? rob_ingress_id_110 : _GEN_10483; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10485 = 7'h6f == out_payload_1_rob_idx[6:0] ? rob_ingress_id_111 : _GEN_10484; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10486 = 7'h70 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_112 : _GEN_10485; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10487 = 7'h71 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_113 : _GEN_10486; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10488 = 7'h72 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_114 : _GEN_10487; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10489 = 7'h73 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_115 : _GEN_10488; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10490 = 7'h74 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_116 : _GEN_10489; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10491 = 7'h75 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_117 : _GEN_10490; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10492 = 7'h76 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_118 : _GEN_10491; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10493 = 7'h77 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_119 : _GEN_10492; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10494 = 7'h78 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_120 : _GEN_10493; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10495 = 7'h79 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_121 : _GEN_10494; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10496 = 7'h7a == out_payload_1_rob_idx[6:0] ? rob_ingress_id_122 : _GEN_10495; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10497 = 7'h7b == out_payload_1_rob_idx[6:0] ? rob_ingress_id_123 : _GEN_10496; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10498 = 7'h7c == out_payload_1_rob_idx[6:0] ? rob_ingress_id_124 : _GEN_10497; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10499 = 7'h7d == out_payload_1_rob_idx[6:0] ? rob_ingress_id_125 : _GEN_10498; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10500 = 7'h7e == out_payload_1_rob_idx[6:0] ? rob_ingress_id_126 : _GEN_10499; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10501 = 7'h7f == out_payload_1_rob_idx[6:0] ? rob_ingress_id_127 : _GEN_10500; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_10503 = 7'h1 == out_payload_1_rob_idx[6:0] ? rob_egress_id_1 : rob_egress_id_0; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10504 = 7'h2 == out_payload_1_rob_idx[6:0] ? rob_egress_id_2 : _GEN_10503; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10505 = 7'h3 == out_payload_1_rob_idx[6:0] ? rob_egress_id_3 : _GEN_10504; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10506 = 7'h4 == out_payload_1_rob_idx[6:0] ? rob_egress_id_4 : _GEN_10505; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10507 = 7'h5 == out_payload_1_rob_idx[6:0] ? rob_egress_id_5 : _GEN_10506; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10508 = 7'h6 == out_payload_1_rob_idx[6:0] ? rob_egress_id_6 : _GEN_10507; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10509 = 7'h7 == out_payload_1_rob_idx[6:0] ? rob_egress_id_7 : _GEN_10508; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10510 = 7'h8 == out_payload_1_rob_idx[6:0] ? rob_egress_id_8 : _GEN_10509; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10511 = 7'h9 == out_payload_1_rob_idx[6:0] ? rob_egress_id_9 : _GEN_10510; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10512 = 7'ha == out_payload_1_rob_idx[6:0] ? rob_egress_id_10 : _GEN_10511; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10513 = 7'hb == out_payload_1_rob_idx[6:0] ? rob_egress_id_11 : _GEN_10512; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10514 = 7'hc == out_payload_1_rob_idx[6:0] ? rob_egress_id_12 : _GEN_10513; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10515 = 7'hd == out_payload_1_rob_idx[6:0] ? rob_egress_id_13 : _GEN_10514; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10516 = 7'he == out_payload_1_rob_idx[6:0] ? rob_egress_id_14 : _GEN_10515; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10517 = 7'hf == out_payload_1_rob_idx[6:0] ? rob_egress_id_15 : _GEN_10516; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10518 = 7'h10 == out_payload_1_rob_idx[6:0] ? rob_egress_id_16 : _GEN_10517; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10519 = 7'h11 == out_payload_1_rob_idx[6:0] ? rob_egress_id_17 : _GEN_10518; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10520 = 7'h12 == out_payload_1_rob_idx[6:0] ? rob_egress_id_18 : _GEN_10519; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10521 = 7'h13 == out_payload_1_rob_idx[6:0] ? rob_egress_id_19 : _GEN_10520; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10522 = 7'h14 == out_payload_1_rob_idx[6:0] ? rob_egress_id_20 : _GEN_10521; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10523 = 7'h15 == out_payload_1_rob_idx[6:0] ? rob_egress_id_21 : _GEN_10522; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10524 = 7'h16 == out_payload_1_rob_idx[6:0] ? rob_egress_id_22 : _GEN_10523; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10525 = 7'h17 == out_payload_1_rob_idx[6:0] ? rob_egress_id_23 : _GEN_10524; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10526 = 7'h18 == out_payload_1_rob_idx[6:0] ? rob_egress_id_24 : _GEN_10525; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10527 = 7'h19 == out_payload_1_rob_idx[6:0] ? rob_egress_id_25 : _GEN_10526; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10528 = 7'h1a == out_payload_1_rob_idx[6:0] ? rob_egress_id_26 : _GEN_10527; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10529 = 7'h1b == out_payload_1_rob_idx[6:0] ? rob_egress_id_27 : _GEN_10528; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10530 = 7'h1c == out_payload_1_rob_idx[6:0] ? rob_egress_id_28 : _GEN_10529; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10531 = 7'h1d == out_payload_1_rob_idx[6:0] ? rob_egress_id_29 : _GEN_10530; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10532 = 7'h1e == out_payload_1_rob_idx[6:0] ? rob_egress_id_30 : _GEN_10531; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10533 = 7'h1f == out_payload_1_rob_idx[6:0] ? rob_egress_id_31 : _GEN_10532; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10534 = 7'h20 == out_payload_1_rob_idx[6:0] ? rob_egress_id_32 : _GEN_10533; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10535 = 7'h21 == out_payload_1_rob_idx[6:0] ? rob_egress_id_33 : _GEN_10534; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10536 = 7'h22 == out_payload_1_rob_idx[6:0] ? rob_egress_id_34 : _GEN_10535; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10537 = 7'h23 == out_payload_1_rob_idx[6:0] ? rob_egress_id_35 : _GEN_10536; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10538 = 7'h24 == out_payload_1_rob_idx[6:0] ? rob_egress_id_36 : _GEN_10537; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10539 = 7'h25 == out_payload_1_rob_idx[6:0] ? rob_egress_id_37 : _GEN_10538; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10540 = 7'h26 == out_payload_1_rob_idx[6:0] ? rob_egress_id_38 : _GEN_10539; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10541 = 7'h27 == out_payload_1_rob_idx[6:0] ? rob_egress_id_39 : _GEN_10540; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10542 = 7'h28 == out_payload_1_rob_idx[6:0] ? rob_egress_id_40 : _GEN_10541; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10543 = 7'h29 == out_payload_1_rob_idx[6:0] ? rob_egress_id_41 : _GEN_10542; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10544 = 7'h2a == out_payload_1_rob_idx[6:0] ? rob_egress_id_42 : _GEN_10543; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10545 = 7'h2b == out_payload_1_rob_idx[6:0] ? rob_egress_id_43 : _GEN_10544; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10546 = 7'h2c == out_payload_1_rob_idx[6:0] ? rob_egress_id_44 : _GEN_10545; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10547 = 7'h2d == out_payload_1_rob_idx[6:0] ? rob_egress_id_45 : _GEN_10546; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10548 = 7'h2e == out_payload_1_rob_idx[6:0] ? rob_egress_id_46 : _GEN_10547; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10549 = 7'h2f == out_payload_1_rob_idx[6:0] ? rob_egress_id_47 : _GEN_10548; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10550 = 7'h30 == out_payload_1_rob_idx[6:0] ? rob_egress_id_48 : _GEN_10549; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10551 = 7'h31 == out_payload_1_rob_idx[6:0] ? rob_egress_id_49 : _GEN_10550; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10552 = 7'h32 == out_payload_1_rob_idx[6:0] ? rob_egress_id_50 : _GEN_10551; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10553 = 7'h33 == out_payload_1_rob_idx[6:0] ? rob_egress_id_51 : _GEN_10552; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10554 = 7'h34 == out_payload_1_rob_idx[6:0] ? rob_egress_id_52 : _GEN_10553; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10555 = 7'h35 == out_payload_1_rob_idx[6:0] ? rob_egress_id_53 : _GEN_10554; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10556 = 7'h36 == out_payload_1_rob_idx[6:0] ? rob_egress_id_54 : _GEN_10555; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10557 = 7'h37 == out_payload_1_rob_idx[6:0] ? rob_egress_id_55 : _GEN_10556; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10558 = 7'h38 == out_payload_1_rob_idx[6:0] ? rob_egress_id_56 : _GEN_10557; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10559 = 7'h39 == out_payload_1_rob_idx[6:0] ? rob_egress_id_57 : _GEN_10558; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10560 = 7'h3a == out_payload_1_rob_idx[6:0] ? rob_egress_id_58 : _GEN_10559; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10561 = 7'h3b == out_payload_1_rob_idx[6:0] ? rob_egress_id_59 : _GEN_10560; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10562 = 7'h3c == out_payload_1_rob_idx[6:0] ? rob_egress_id_60 : _GEN_10561; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10563 = 7'h3d == out_payload_1_rob_idx[6:0] ? rob_egress_id_61 : _GEN_10562; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10564 = 7'h3e == out_payload_1_rob_idx[6:0] ? rob_egress_id_62 : _GEN_10563; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10565 = 7'h3f == out_payload_1_rob_idx[6:0] ? rob_egress_id_63 : _GEN_10564; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10566 = 7'h40 == out_payload_1_rob_idx[6:0] ? rob_egress_id_64 : _GEN_10565; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10567 = 7'h41 == out_payload_1_rob_idx[6:0] ? rob_egress_id_65 : _GEN_10566; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10568 = 7'h42 == out_payload_1_rob_idx[6:0] ? rob_egress_id_66 : _GEN_10567; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10569 = 7'h43 == out_payload_1_rob_idx[6:0] ? rob_egress_id_67 : _GEN_10568; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10570 = 7'h44 == out_payload_1_rob_idx[6:0] ? rob_egress_id_68 : _GEN_10569; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10571 = 7'h45 == out_payload_1_rob_idx[6:0] ? rob_egress_id_69 : _GEN_10570; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10572 = 7'h46 == out_payload_1_rob_idx[6:0] ? rob_egress_id_70 : _GEN_10571; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10573 = 7'h47 == out_payload_1_rob_idx[6:0] ? rob_egress_id_71 : _GEN_10572; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10574 = 7'h48 == out_payload_1_rob_idx[6:0] ? rob_egress_id_72 : _GEN_10573; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10575 = 7'h49 == out_payload_1_rob_idx[6:0] ? rob_egress_id_73 : _GEN_10574; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10576 = 7'h4a == out_payload_1_rob_idx[6:0] ? rob_egress_id_74 : _GEN_10575; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10577 = 7'h4b == out_payload_1_rob_idx[6:0] ? rob_egress_id_75 : _GEN_10576; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10578 = 7'h4c == out_payload_1_rob_idx[6:0] ? rob_egress_id_76 : _GEN_10577; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10579 = 7'h4d == out_payload_1_rob_idx[6:0] ? rob_egress_id_77 : _GEN_10578; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10580 = 7'h4e == out_payload_1_rob_idx[6:0] ? rob_egress_id_78 : _GEN_10579; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10581 = 7'h4f == out_payload_1_rob_idx[6:0] ? rob_egress_id_79 : _GEN_10580; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10582 = 7'h50 == out_payload_1_rob_idx[6:0] ? rob_egress_id_80 : _GEN_10581; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10583 = 7'h51 == out_payload_1_rob_idx[6:0] ? rob_egress_id_81 : _GEN_10582; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10584 = 7'h52 == out_payload_1_rob_idx[6:0] ? rob_egress_id_82 : _GEN_10583; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10585 = 7'h53 == out_payload_1_rob_idx[6:0] ? rob_egress_id_83 : _GEN_10584; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10586 = 7'h54 == out_payload_1_rob_idx[6:0] ? rob_egress_id_84 : _GEN_10585; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10587 = 7'h55 == out_payload_1_rob_idx[6:0] ? rob_egress_id_85 : _GEN_10586; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10588 = 7'h56 == out_payload_1_rob_idx[6:0] ? rob_egress_id_86 : _GEN_10587; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10589 = 7'h57 == out_payload_1_rob_idx[6:0] ? rob_egress_id_87 : _GEN_10588; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10590 = 7'h58 == out_payload_1_rob_idx[6:0] ? rob_egress_id_88 : _GEN_10589; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10591 = 7'h59 == out_payload_1_rob_idx[6:0] ? rob_egress_id_89 : _GEN_10590; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10592 = 7'h5a == out_payload_1_rob_idx[6:0] ? rob_egress_id_90 : _GEN_10591; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10593 = 7'h5b == out_payload_1_rob_idx[6:0] ? rob_egress_id_91 : _GEN_10592; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10594 = 7'h5c == out_payload_1_rob_idx[6:0] ? rob_egress_id_92 : _GEN_10593; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10595 = 7'h5d == out_payload_1_rob_idx[6:0] ? rob_egress_id_93 : _GEN_10594; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10596 = 7'h5e == out_payload_1_rob_idx[6:0] ? rob_egress_id_94 : _GEN_10595; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10597 = 7'h5f == out_payload_1_rob_idx[6:0] ? rob_egress_id_95 : _GEN_10596; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10598 = 7'h60 == out_payload_1_rob_idx[6:0] ? rob_egress_id_96 : _GEN_10597; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10599 = 7'h61 == out_payload_1_rob_idx[6:0] ? rob_egress_id_97 : _GEN_10598; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10600 = 7'h62 == out_payload_1_rob_idx[6:0] ? rob_egress_id_98 : _GEN_10599; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10601 = 7'h63 == out_payload_1_rob_idx[6:0] ? rob_egress_id_99 : _GEN_10600; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10602 = 7'h64 == out_payload_1_rob_idx[6:0] ? rob_egress_id_100 : _GEN_10601; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10603 = 7'h65 == out_payload_1_rob_idx[6:0] ? rob_egress_id_101 : _GEN_10602; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10604 = 7'h66 == out_payload_1_rob_idx[6:0] ? rob_egress_id_102 : _GEN_10603; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10605 = 7'h67 == out_payload_1_rob_idx[6:0] ? rob_egress_id_103 : _GEN_10604; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10606 = 7'h68 == out_payload_1_rob_idx[6:0] ? rob_egress_id_104 : _GEN_10605; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10607 = 7'h69 == out_payload_1_rob_idx[6:0] ? rob_egress_id_105 : _GEN_10606; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10608 = 7'h6a == out_payload_1_rob_idx[6:0] ? rob_egress_id_106 : _GEN_10607; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10609 = 7'h6b == out_payload_1_rob_idx[6:0] ? rob_egress_id_107 : _GEN_10608; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10610 = 7'h6c == out_payload_1_rob_idx[6:0] ? rob_egress_id_108 : _GEN_10609; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10611 = 7'h6d == out_payload_1_rob_idx[6:0] ? rob_egress_id_109 : _GEN_10610; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10612 = 7'h6e == out_payload_1_rob_idx[6:0] ? rob_egress_id_110 : _GEN_10611; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10613 = 7'h6f == out_payload_1_rob_idx[6:0] ? rob_egress_id_111 : _GEN_10612; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10614 = 7'h70 == out_payload_1_rob_idx[6:0] ? rob_egress_id_112 : _GEN_10613; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10615 = 7'h71 == out_payload_1_rob_idx[6:0] ? rob_egress_id_113 : _GEN_10614; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10616 = 7'h72 == out_payload_1_rob_idx[6:0] ? rob_egress_id_114 : _GEN_10615; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10617 = 7'h73 == out_payload_1_rob_idx[6:0] ? rob_egress_id_115 : _GEN_10616; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10618 = 7'h74 == out_payload_1_rob_idx[6:0] ? rob_egress_id_116 : _GEN_10617; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10619 = 7'h75 == out_payload_1_rob_idx[6:0] ? rob_egress_id_117 : _GEN_10618; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10620 = 7'h76 == out_payload_1_rob_idx[6:0] ? rob_egress_id_118 : _GEN_10619; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10621 = 7'h77 == out_payload_1_rob_idx[6:0] ? rob_egress_id_119 : _GEN_10620; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10622 = 7'h78 == out_payload_1_rob_idx[6:0] ? rob_egress_id_120 : _GEN_10621; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10623 = 7'h79 == out_payload_1_rob_idx[6:0] ? rob_egress_id_121 : _GEN_10622; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10624 = 7'h7a == out_payload_1_rob_idx[6:0] ? rob_egress_id_122 : _GEN_10623; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10625 = 7'h7b == out_payload_1_rob_idx[6:0] ? rob_egress_id_123 : _GEN_10624; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10626 = 7'h7c == out_payload_1_rob_idx[6:0] ? rob_egress_id_124 : _GEN_10625; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10627 = 7'h7d == out_payload_1_rob_idx[6:0] ? rob_egress_id_125 : _GEN_10626; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10628 = 7'h7e == out_payload_1_rob_idx[6:0] ? rob_egress_id_126 : _GEN_10627; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_10629 = 7'h7f == out_payload_1_rob_idx[6:0] ? rob_egress_id_127 : _GEN_10628; // @[TestHarness.scala 204:{18,18}]
  wire [3:0] _GEN_10631 = 7'h1 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_1 : rob_flits_returned_0; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10632 = 7'h2 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_2 : _GEN_10631; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10633 = 7'h3 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_3 : _GEN_10632; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10634 = 7'h4 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_4 : _GEN_10633; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10635 = 7'h5 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_5 : _GEN_10634; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10636 = 7'h6 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_6 : _GEN_10635; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10637 = 7'h7 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_7 : _GEN_10636; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10638 = 7'h8 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_8 : _GEN_10637; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10639 = 7'h9 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_9 : _GEN_10638; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10640 = 7'ha == out_payload_1_rob_idx[6:0] ? rob_flits_returned_10 : _GEN_10639; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10641 = 7'hb == out_payload_1_rob_idx[6:0] ? rob_flits_returned_11 : _GEN_10640; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10642 = 7'hc == out_payload_1_rob_idx[6:0] ? rob_flits_returned_12 : _GEN_10641; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10643 = 7'hd == out_payload_1_rob_idx[6:0] ? rob_flits_returned_13 : _GEN_10642; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10644 = 7'he == out_payload_1_rob_idx[6:0] ? rob_flits_returned_14 : _GEN_10643; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10645 = 7'hf == out_payload_1_rob_idx[6:0] ? rob_flits_returned_15 : _GEN_10644; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10646 = 7'h10 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_16 : _GEN_10645; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10647 = 7'h11 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_17 : _GEN_10646; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10648 = 7'h12 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_18 : _GEN_10647; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10649 = 7'h13 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_19 : _GEN_10648; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10650 = 7'h14 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_20 : _GEN_10649; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10651 = 7'h15 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_21 : _GEN_10650; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10652 = 7'h16 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_22 : _GEN_10651; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10653 = 7'h17 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_23 : _GEN_10652; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10654 = 7'h18 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_24 : _GEN_10653; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10655 = 7'h19 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_25 : _GEN_10654; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10656 = 7'h1a == out_payload_1_rob_idx[6:0] ? rob_flits_returned_26 : _GEN_10655; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10657 = 7'h1b == out_payload_1_rob_idx[6:0] ? rob_flits_returned_27 : _GEN_10656; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10658 = 7'h1c == out_payload_1_rob_idx[6:0] ? rob_flits_returned_28 : _GEN_10657; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10659 = 7'h1d == out_payload_1_rob_idx[6:0] ? rob_flits_returned_29 : _GEN_10658; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10660 = 7'h1e == out_payload_1_rob_idx[6:0] ? rob_flits_returned_30 : _GEN_10659; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10661 = 7'h1f == out_payload_1_rob_idx[6:0] ? rob_flits_returned_31 : _GEN_10660; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10662 = 7'h20 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_32 : _GEN_10661; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10663 = 7'h21 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_33 : _GEN_10662; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10664 = 7'h22 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_34 : _GEN_10663; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10665 = 7'h23 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_35 : _GEN_10664; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10666 = 7'h24 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_36 : _GEN_10665; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10667 = 7'h25 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_37 : _GEN_10666; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10668 = 7'h26 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_38 : _GEN_10667; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10669 = 7'h27 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_39 : _GEN_10668; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10670 = 7'h28 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_40 : _GEN_10669; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10671 = 7'h29 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_41 : _GEN_10670; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10672 = 7'h2a == out_payload_1_rob_idx[6:0] ? rob_flits_returned_42 : _GEN_10671; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10673 = 7'h2b == out_payload_1_rob_idx[6:0] ? rob_flits_returned_43 : _GEN_10672; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10674 = 7'h2c == out_payload_1_rob_idx[6:0] ? rob_flits_returned_44 : _GEN_10673; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10675 = 7'h2d == out_payload_1_rob_idx[6:0] ? rob_flits_returned_45 : _GEN_10674; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10676 = 7'h2e == out_payload_1_rob_idx[6:0] ? rob_flits_returned_46 : _GEN_10675; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10677 = 7'h2f == out_payload_1_rob_idx[6:0] ? rob_flits_returned_47 : _GEN_10676; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10678 = 7'h30 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_48 : _GEN_10677; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10679 = 7'h31 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_49 : _GEN_10678; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10680 = 7'h32 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_50 : _GEN_10679; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10681 = 7'h33 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_51 : _GEN_10680; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10682 = 7'h34 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_52 : _GEN_10681; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10683 = 7'h35 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_53 : _GEN_10682; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10684 = 7'h36 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_54 : _GEN_10683; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10685 = 7'h37 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_55 : _GEN_10684; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10686 = 7'h38 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_56 : _GEN_10685; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10687 = 7'h39 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_57 : _GEN_10686; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10688 = 7'h3a == out_payload_1_rob_idx[6:0] ? rob_flits_returned_58 : _GEN_10687; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10689 = 7'h3b == out_payload_1_rob_idx[6:0] ? rob_flits_returned_59 : _GEN_10688; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10690 = 7'h3c == out_payload_1_rob_idx[6:0] ? rob_flits_returned_60 : _GEN_10689; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10691 = 7'h3d == out_payload_1_rob_idx[6:0] ? rob_flits_returned_61 : _GEN_10690; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10692 = 7'h3e == out_payload_1_rob_idx[6:0] ? rob_flits_returned_62 : _GEN_10691; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10693 = 7'h3f == out_payload_1_rob_idx[6:0] ? rob_flits_returned_63 : _GEN_10692; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10694 = 7'h40 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_64 : _GEN_10693; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10695 = 7'h41 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_65 : _GEN_10694; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10696 = 7'h42 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_66 : _GEN_10695; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10697 = 7'h43 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_67 : _GEN_10696; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10698 = 7'h44 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_68 : _GEN_10697; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10699 = 7'h45 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_69 : _GEN_10698; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10700 = 7'h46 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_70 : _GEN_10699; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10701 = 7'h47 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_71 : _GEN_10700; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10702 = 7'h48 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_72 : _GEN_10701; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10703 = 7'h49 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_73 : _GEN_10702; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10704 = 7'h4a == out_payload_1_rob_idx[6:0] ? rob_flits_returned_74 : _GEN_10703; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10705 = 7'h4b == out_payload_1_rob_idx[6:0] ? rob_flits_returned_75 : _GEN_10704; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10706 = 7'h4c == out_payload_1_rob_idx[6:0] ? rob_flits_returned_76 : _GEN_10705; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10707 = 7'h4d == out_payload_1_rob_idx[6:0] ? rob_flits_returned_77 : _GEN_10706; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10708 = 7'h4e == out_payload_1_rob_idx[6:0] ? rob_flits_returned_78 : _GEN_10707; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10709 = 7'h4f == out_payload_1_rob_idx[6:0] ? rob_flits_returned_79 : _GEN_10708; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10710 = 7'h50 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_80 : _GEN_10709; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10711 = 7'h51 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_81 : _GEN_10710; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10712 = 7'h52 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_82 : _GEN_10711; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10713 = 7'h53 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_83 : _GEN_10712; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10714 = 7'h54 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_84 : _GEN_10713; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10715 = 7'h55 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_85 : _GEN_10714; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10716 = 7'h56 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_86 : _GEN_10715; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10717 = 7'h57 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_87 : _GEN_10716; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10718 = 7'h58 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_88 : _GEN_10717; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10719 = 7'h59 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_89 : _GEN_10718; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10720 = 7'h5a == out_payload_1_rob_idx[6:0] ? rob_flits_returned_90 : _GEN_10719; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10721 = 7'h5b == out_payload_1_rob_idx[6:0] ? rob_flits_returned_91 : _GEN_10720; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10722 = 7'h5c == out_payload_1_rob_idx[6:0] ? rob_flits_returned_92 : _GEN_10721; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10723 = 7'h5d == out_payload_1_rob_idx[6:0] ? rob_flits_returned_93 : _GEN_10722; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10724 = 7'h5e == out_payload_1_rob_idx[6:0] ? rob_flits_returned_94 : _GEN_10723; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10725 = 7'h5f == out_payload_1_rob_idx[6:0] ? rob_flits_returned_95 : _GEN_10724; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10726 = 7'h60 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_96 : _GEN_10725; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10727 = 7'h61 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_97 : _GEN_10726; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10728 = 7'h62 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_98 : _GEN_10727; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10729 = 7'h63 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_99 : _GEN_10728; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10730 = 7'h64 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_100 : _GEN_10729; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10731 = 7'h65 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_101 : _GEN_10730; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10732 = 7'h66 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_102 : _GEN_10731; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10733 = 7'h67 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_103 : _GEN_10732; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10734 = 7'h68 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_104 : _GEN_10733; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10735 = 7'h69 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_105 : _GEN_10734; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10736 = 7'h6a == out_payload_1_rob_idx[6:0] ? rob_flits_returned_106 : _GEN_10735; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10737 = 7'h6b == out_payload_1_rob_idx[6:0] ? rob_flits_returned_107 : _GEN_10736; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10738 = 7'h6c == out_payload_1_rob_idx[6:0] ? rob_flits_returned_108 : _GEN_10737; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10739 = 7'h6d == out_payload_1_rob_idx[6:0] ? rob_flits_returned_109 : _GEN_10738; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10740 = 7'h6e == out_payload_1_rob_idx[6:0] ? rob_flits_returned_110 : _GEN_10739; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10741 = 7'h6f == out_payload_1_rob_idx[6:0] ? rob_flits_returned_111 : _GEN_10740; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10742 = 7'h70 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_112 : _GEN_10741; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10743 = 7'h71 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_113 : _GEN_10742; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10744 = 7'h72 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_114 : _GEN_10743; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10745 = 7'h73 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_115 : _GEN_10744; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10746 = 7'h74 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_116 : _GEN_10745; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10747 = 7'h75 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_117 : _GEN_10746; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10748 = 7'h76 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_118 : _GEN_10747; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10749 = 7'h77 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_119 : _GEN_10748; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10750 = 7'h78 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_120 : _GEN_10749; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10751 = 7'h79 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_121 : _GEN_10750; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10752 = 7'h7a == out_payload_1_rob_idx[6:0] ? rob_flits_returned_122 : _GEN_10751; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10753 = 7'h7b == out_payload_1_rob_idx[6:0] ? rob_flits_returned_123 : _GEN_10752; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10754 = 7'h7c == out_payload_1_rob_idx[6:0] ? rob_flits_returned_124 : _GEN_10753; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10755 = 7'h7d == out_payload_1_rob_idx[6:0] ? rob_flits_returned_125 : _GEN_10754; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10756 = 7'h7e == out_payload_1_rob_idx[6:0] ? rob_flits_returned_126 : _GEN_10755; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10757 = 7'h7f == out_payload_1_rob_idx[6:0] ? rob_flits_returned_127 : _GEN_10756; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10759 = 7'h1 == out_payload_1_rob_idx[6:0] ? rob_n_flits_1 : rob_n_flits_0; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10760 = 7'h2 == out_payload_1_rob_idx[6:0] ? rob_n_flits_2 : _GEN_10759; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10761 = 7'h3 == out_payload_1_rob_idx[6:0] ? rob_n_flits_3 : _GEN_10760; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10762 = 7'h4 == out_payload_1_rob_idx[6:0] ? rob_n_flits_4 : _GEN_10761; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10763 = 7'h5 == out_payload_1_rob_idx[6:0] ? rob_n_flits_5 : _GEN_10762; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10764 = 7'h6 == out_payload_1_rob_idx[6:0] ? rob_n_flits_6 : _GEN_10763; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10765 = 7'h7 == out_payload_1_rob_idx[6:0] ? rob_n_flits_7 : _GEN_10764; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10766 = 7'h8 == out_payload_1_rob_idx[6:0] ? rob_n_flits_8 : _GEN_10765; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10767 = 7'h9 == out_payload_1_rob_idx[6:0] ? rob_n_flits_9 : _GEN_10766; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10768 = 7'ha == out_payload_1_rob_idx[6:0] ? rob_n_flits_10 : _GEN_10767; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10769 = 7'hb == out_payload_1_rob_idx[6:0] ? rob_n_flits_11 : _GEN_10768; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10770 = 7'hc == out_payload_1_rob_idx[6:0] ? rob_n_flits_12 : _GEN_10769; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10771 = 7'hd == out_payload_1_rob_idx[6:0] ? rob_n_flits_13 : _GEN_10770; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10772 = 7'he == out_payload_1_rob_idx[6:0] ? rob_n_flits_14 : _GEN_10771; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10773 = 7'hf == out_payload_1_rob_idx[6:0] ? rob_n_flits_15 : _GEN_10772; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10774 = 7'h10 == out_payload_1_rob_idx[6:0] ? rob_n_flits_16 : _GEN_10773; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10775 = 7'h11 == out_payload_1_rob_idx[6:0] ? rob_n_flits_17 : _GEN_10774; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10776 = 7'h12 == out_payload_1_rob_idx[6:0] ? rob_n_flits_18 : _GEN_10775; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10777 = 7'h13 == out_payload_1_rob_idx[6:0] ? rob_n_flits_19 : _GEN_10776; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10778 = 7'h14 == out_payload_1_rob_idx[6:0] ? rob_n_flits_20 : _GEN_10777; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10779 = 7'h15 == out_payload_1_rob_idx[6:0] ? rob_n_flits_21 : _GEN_10778; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10780 = 7'h16 == out_payload_1_rob_idx[6:0] ? rob_n_flits_22 : _GEN_10779; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10781 = 7'h17 == out_payload_1_rob_idx[6:0] ? rob_n_flits_23 : _GEN_10780; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10782 = 7'h18 == out_payload_1_rob_idx[6:0] ? rob_n_flits_24 : _GEN_10781; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10783 = 7'h19 == out_payload_1_rob_idx[6:0] ? rob_n_flits_25 : _GEN_10782; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10784 = 7'h1a == out_payload_1_rob_idx[6:0] ? rob_n_flits_26 : _GEN_10783; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10785 = 7'h1b == out_payload_1_rob_idx[6:0] ? rob_n_flits_27 : _GEN_10784; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10786 = 7'h1c == out_payload_1_rob_idx[6:0] ? rob_n_flits_28 : _GEN_10785; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10787 = 7'h1d == out_payload_1_rob_idx[6:0] ? rob_n_flits_29 : _GEN_10786; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10788 = 7'h1e == out_payload_1_rob_idx[6:0] ? rob_n_flits_30 : _GEN_10787; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10789 = 7'h1f == out_payload_1_rob_idx[6:0] ? rob_n_flits_31 : _GEN_10788; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10790 = 7'h20 == out_payload_1_rob_idx[6:0] ? rob_n_flits_32 : _GEN_10789; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10791 = 7'h21 == out_payload_1_rob_idx[6:0] ? rob_n_flits_33 : _GEN_10790; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10792 = 7'h22 == out_payload_1_rob_idx[6:0] ? rob_n_flits_34 : _GEN_10791; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10793 = 7'h23 == out_payload_1_rob_idx[6:0] ? rob_n_flits_35 : _GEN_10792; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10794 = 7'h24 == out_payload_1_rob_idx[6:0] ? rob_n_flits_36 : _GEN_10793; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10795 = 7'h25 == out_payload_1_rob_idx[6:0] ? rob_n_flits_37 : _GEN_10794; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10796 = 7'h26 == out_payload_1_rob_idx[6:0] ? rob_n_flits_38 : _GEN_10795; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10797 = 7'h27 == out_payload_1_rob_idx[6:0] ? rob_n_flits_39 : _GEN_10796; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10798 = 7'h28 == out_payload_1_rob_idx[6:0] ? rob_n_flits_40 : _GEN_10797; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10799 = 7'h29 == out_payload_1_rob_idx[6:0] ? rob_n_flits_41 : _GEN_10798; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10800 = 7'h2a == out_payload_1_rob_idx[6:0] ? rob_n_flits_42 : _GEN_10799; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10801 = 7'h2b == out_payload_1_rob_idx[6:0] ? rob_n_flits_43 : _GEN_10800; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10802 = 7'h2c == out_payload_1_rob_idx[6:0] ? rob_n_flits_44 : _GEN_10801; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10803 = 7'h2d == out_payload_1_rob_idx[6:0] ? rob_n_flits_45 : _GEN_10802; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10804 = 7'h2e == out_payload_1_rob_idx[6:0] ? rob_n_flits_46 : _GEN_10803; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10805 = 7'h2f == out_payload_1_rob_idx[6:0] ? rob_n_flits_47 : _GEN_10804; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10806 = 7'h30 == out_payload_1_rob_idx[6:0] ? rob_n_flits_48 : _GEN_10805; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10807 = 7'h31 == out_payload_1_rob_idx[6:0] ? rob_n_flits_49 : _GEN_10806; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10808 = 7'h32 == out_payload_1_rob_idx[6:0] ? rob_n_flits_50 : _GEN_10807; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10809 = 7'h33 == out_payload_1_rob_idx[6:0] ? rob_n_flits_51 : _GEN_10808; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10810 = 7'h34 == out_payload_1_rob_idx[6:0] ? rob_n_flits_52 : _GEN_10809; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10811 = 7'h35 == out_payload_1_rob_idx[6:0] ? rob_n_flits_53 : _GEN_10810; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10812 = 7'h36 == out_payload_1_rob_idx[6:0] ? rob_n_flits_54 : _GEN_10811; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10813 = 7'h37 == out_payload_1_rob_idx[6:0] ? rob_n_flits_55 : _GEN_10812; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10814 = 7'h38 == out_payload_1_rob_idx[6:0] ? rob_n_flits_56 : _GEN_10813; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10815 = 7'h39 == out_payload_1_rob_idx[6:0] ? rob_n_flits_57 : _GEN_10814; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10816 = 7'h3a == out_payload_1_rob_idx[6:0] ? rob_n_flits_58 : _GEN_10815; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10817 = 7'h3b == out_payload_1_rob_idx[6:0] ? rob_n_flits_59 : _GEN_10816; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10818 = 7'h3c == out_payload_1_rob_idx[6:0] ? rob_n_flits_60 : _GEN_10817; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10819 = 7'h3d == out_payload_1_rob_idx[6:0] ? rob_n_flits_61 : _GEN_10818; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10820 = 7'h3e == out_payload_1_rob_idx[6:0] ? rob_n_flits_62 : _GEN_10819; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10821 = 7'h3f == out_payload_1_rob_idx[6:0] ? rob_n_flits_63 : _GEN_10820; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10822 = 7'h40 == out_payload_1_rob_idx[6:0] ? rob_n_flits_64 : _GEN_10821; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10823 = 7'h41 == out_payload_1_rob_idx[6:0] ? rob_n_flits_65 : _GEN_10822; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10824 = 7'h42 == out_payload_1_rob_idx[6:0] ? rob_n_flits_66 : _GEN_10823; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10825 = 7'h43 == out_payload_1_rob_idx[6:0] ? rob_n_flits_67 : _GEN_10824; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10826 = 7'h44 == out_payload_1_rob_idx[6:0] ? rob_n_flits_68 : _GEN_10825; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10827 = 7'h45 == out_payload_1_rob_idx[6:0] ? rob_n_flits_69 : _GEN_10826; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10828 = 7'h46 == out_payload_1_rob_idx[6:0] ? rob_n_flits_70 : _GEN_10827; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10829 = 7'h47 == out_payload_1_rob_idx[6:0] ? rob_n_flits_71 : _GEN_10828; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10830 = 7'h48 == out_payload_1_rob_idx[6:0] ? rob_n_flits_72 : _GEN_10829; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10831 = 7'h49 == out_payload_1_rob_idx[6:0] ? rob_n_flits_73 : _GEN_10830; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10832 = 7'h4a == out_payload_1_rob_idx[6:0] ? rob_n_flits_74 : _GEN_10831; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10833 = 7'h4b == out_payload_1_rob_idx[6:0] ? rob_n_flits_75 : _GEN_10832; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10834 = 7'h4c == out_payload_1_rob_idx[6:0] ? rob_n_flits_76 : _GEN_10833; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10835 = 7'h4d == out_payload_1_rob_idx[6:0] ? rob_n_flits_77 : _GEN_10834; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10836 = 7'h4e == out_payload_1_rob_idx[6:0] ? rob_n_flits_78 : _GEN_10835; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10837 = 7'h4f == out_payload_1_rob_idx[6:0] ? rob_n_flits_79 : _GEN_10836; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10838 = 7'h50 == out_payload_1_rob_idx[6:0] ? rob_n_flits_80 : _GEN_10837; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10839 = 7'h51 == out_payload_1_rob_idx[6:0] ? rob_n_flits_81 : _GEN_10838; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10840 = 7'h52 == out_payload_1_rob_idx[6:0] ? rob_n_flits_82 : _GEN_10839; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10841 = 7'h53 == out_payload_1_rob_idx[6:0] ? rob_n_flits_83 : _GEN_10840; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10842 = 7'h54 == out_payload_1_rob_idx[6:0] ? rob_n_flits_84 : _GEN_10841; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10843 = 7'h55 == out_payload_1_rob_idx[6:0] ? rob_n_flits_85 : _GEN_10842; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10844 = 7'h56 == out_payload_1_rob_idx[6:0] ? rob_n_flits_86 : _GEN_10843; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10845 = 7'h57 == out_payload_1_rob_idx[6:0] ? rob_n_flits_87 : _GEN_10844; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10846 = 7'h58 == out_payload_1_rob_idx[6:0] ? rob_n_flits_88 : _GEN_10845; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10847 = 7'h59 == out_payload_1_rob_idx[6:0] ? rob_n_flits_89 : _GEN_10846; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10848 = 7'h5a == out_payload_1_rob_idx[6:0] ? rob_n_flits_90 : _GEN_10847; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10849 = 7'h5b == out_payload_1_rob_idx[6:0] ? rob_n_flits_91 : _GEN_10848; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10850 = 7'h5c == out_payload_1_rob_idx[6:0] ? rob_n_flits_92 : _GEN_10849; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10851 = 7'h5d == out_payload_1_rob_idx[6:0] ? rob_n_flits_93 : _GEN_10850; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10852 = 7'h5e == out_payload_1_rob_idx[6:0] ? rob_n_flits_94 : _GEN_10851; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10853 = 7'h5f == out_payload_1_rob_idx[6:0] ? rob_n_flits_95 : _GEN_10852; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10854 = 7'h60 == out_payload_1_rob_idx[6:0] ? rob_n_flits_96 : _GEN_10853; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10855 = 7'h61 == out_payload_1_rob_idx[6:0] ? rob_n_flits_97 : _GEN_10854; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10856 = 7'h62 == out_payload_1_rob_idx[6:0] ? rob_n_flits_98 : _GEN_10855; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10857 = 7'h63 == out_payload_1_rob_idx[6:0] ? rob_n_flits_99 : _GEN_10856; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10858 = 7'h64 == out_payload_1_rob_idx[6:0] ? rob_n_flits_100 : _GEN_10857; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10859 = 7'h65 == out_payload_1_rob_idx[6:0] ? rob_n_flits_101 : _GEN_10858; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10860 = 7'h66 == out_payload_1_rob_idx[6:0] ? rob_n_flits_102 : _GEN_10859; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10861 = 7'h67 == out_payload_1_rob_idx[6:0] ? rob_n_flits_103 : _GEN_10860; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10862 = 7'h68 == out_payload_1_rob_idx[6:0] ? rob_n_flits_104 : _GEN_10861; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10863 = 7'h69 == out_payload_1_rob_idx[6:0] ? rob_n_flits_105 : _GEN_10862; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10864 = 7'h6a == out_payload_1_rob_idx[6:0] ? rob_n_flits_106 : _GEN_10863; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10865 = 7'h6b == out_payload_1_rob_idx[6:0] ? rob_n_flits_107 : _GEN_10864; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10866 = 7'h6c == out_payload_1_rob_idx[6:0] ? rob_n_flits_108 : _GEN_10865; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10867 = 7'h6d == out_payload_1_rob_idx[6:0] ? rob_n_flits_109 : _GEN_10866; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10868 = 7'h6e == out_payload_1_rob_idx[6:0] ? rob_n_flits_110 : _GEN_10867; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10869 = 7'h6f == out_payload_1_rob_idx[6:0] ? rob_n_flits_111 : _GEN_10868; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10870 = 7'h70 == out_payload_1_rob_idx[6:0] ? rob_n_flits_112 : _GEN_10869; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10871 = 7'h71 == out_payload_1_rob_idx[6:0] ? rob_n_flits_113 : _GEN_10870; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10872 = 7'h72 == out_payload_1_rob_idx[6:0] ? rob_n_flits_114 : _GEN_10871; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10873 = 7'h73 == out_payload_1_rob_idx[6:0] ? rob_n_flits_115 : _GEN_10872; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10874 = 7'h74 == out_payload_1_rob_idx[6:0] ? rob_n_flits_116 : _GEN_10873; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10875 = 7'h75 == out_payload_1_rob_idx[6:0] ? rob_n_flits_117 : _GEN_10874; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10876 = 7'h76 == out_payload_1_rob_idx[6:0] ? rob_n_flits_118 : _GEN_10875; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10877 = 7'h77 == out_payload_1_rob_idx[6:0] ? rob_n_flits_119 : _GEN_10876; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10878 = 7'h78 == out_payload_1_rob_idx[6:0] ? rob_n_flits_120 : _GEN_10877; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10879 = 7'h79 == out_payload_1_rob_idx[6:0] ? rob_n_flits_121 : _GEN_10878; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10880 = 7'h7a == out_payload_1_rob_idx[6:0] ? rob_n_flits_122 : _GEN_10879; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10881 = 7'h7b == out_payload_1_rob_idx[6:0] ? rob_n_flits_123 : _GEN_10880; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10882 = 7'h7c == out_payload_1_rob_idx[6:0] ? rob_n_flits_124 : _GEN_10881; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10883 = 7'h7d == out_payload_1_rob_idx[6:0] ? rob_n_flits_125 : _GEN_10882; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10884 = 7'h7e == out_payload_1_rob_idx[6:0] ? rob_n_flits_126 : _GEN_10883; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_10885 = 7'h7f == out_payload_1_rob_idx[6:0] ? rob_n_flits_127 : _GEN_10884; // @[TestHarness.scala 205:{42,42}]
  wire [15:0] _GEN_15382 = {{9'd0}, packet_rob_idx_1}; // @[TestHarness.scala 206:61]
  wire  _T_157 = io_from_noc_1_flit_bits_head & enable_print_latency; // @[TestHarness.scala 208:30]
  wire [3:0] _rob_flits_returned_T_5 = _GEN_10757 + 4'h1; // @[TestHarness.scala 213:66]
  wire [3:0] _GEN_11142 = 7'h0 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9732; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11143 = 7'h1 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9733; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11144 = 7'h2 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9734; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11145 = 7'h3 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9735; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11146 = 7'h4 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9736; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11147 = 7'h5 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9737; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11148 = 7'h6 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9738; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11149 = 7'h7 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9739; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11150 = 7'h8 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9740; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11151 = 7'h9 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9741; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11152 = 7'ha == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9742; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11153 = 7'hb == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9743; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11154 = 7'hc == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9744; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11155 = 7'hd == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9745; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11156 = 7'he == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9746; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11157 = 7'hf == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9747; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11158 = 7'h10 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9748; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11159 = 7'h11 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9749; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11160 = 7'h12 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9750; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11161 = 7'h13 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9751; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11162 = 7'h14 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9752; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11163 = 7'h15 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9753; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11164 = 7'h16 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9754; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11165 = 7'h17 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9755; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11166 = 7'h18 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9756; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11167 = 7'h19 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9757; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11168 = 7'h1a == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9758; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11169 = 7'h1b == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9759; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11170 = 7'h1c == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9760; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11171 = 7'h1d == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9761; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11172 = 7'h1e == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9762; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11173 = 7'h1f == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9763; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11174 = 7'h20 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9764; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11175 = 7'h21 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9765; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11176 = 7'h22 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9766; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11177 = 7'h23 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9767; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11178 = 7'h24 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9768; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11179 = 7'h25 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9769; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11180 = 7'h26 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9770; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11181 = 7'h27 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9771; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11182 = 7'h28 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9772; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11183 = 7'h29 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9773; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11184 = 7'h2a == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9774; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11185 = 7'h2b == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9775; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11186 = 7'h2c == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9776; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11187 = 7'h2d == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9777; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11188 = 7'h2e == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9778; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11189 = 7'h2f == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9779; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11190 = 7'h30 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9780; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11191 = 7'h31 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9781; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11192 = 7'h32 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9782; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11193 = 7'h33 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9783; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11194 = 7'h34 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9784; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11195 = 7'h35 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9785; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11196 = 7'h36 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9786; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11197 = 7'h37 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9787; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11198 = 7'h38 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9788; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11199 = 7'h39 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9789; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11200 = 7'h3a == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9790; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11201 = 7'h3b == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9791; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11202 = 7'h3c == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9792; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11203 = 7'h3d == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9793; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11204 = 7'h3e == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9794; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11205 = 7'h3f == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9795; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11206 = 7'h40 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9796; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11207 = 7'h41 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9797; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11208 = 7'h42 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9798; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11209 = 7'h43 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9799; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11210 = 7'h44 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9800; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11211 = 7'h45 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9801; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11212 = 7'h46 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9802; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11213 = 7'h47 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9803; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11214 = 7'h48 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9804; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11215 = 7'h49 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9805; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11216 = 7'h4a == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9806; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11217 = 7'h4b == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9807; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11218 = 7'h4c == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9808; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11219 = 7'h4d == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9809; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11220 = 7'h4e == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9810; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11221 = 7'h4f == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9811; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11222 = 7'h50 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9812; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11223 = 7'h51 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9813; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11224 = 7'h52 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9814; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11225 = 7'h53 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9815; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11226 = 7'h54 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9816; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11227 = 7'h55 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9817; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11228 = 7'h56 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9818; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11229 = 7'h57 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9819; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11230 = 7'h58 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9820; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11231 = 7'h59 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9821; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11232 = 7'h5a == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9822; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11233 = 7'h5b == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9823; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11234 = 7'h5c == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9824; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11235 = 7'h5d == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9825; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11236 = 7'h5e == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9826; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11237 = 7'h5f == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9827; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11238 = 7'h60 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9828; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11239 = 7'h61 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9829; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11240 = 7'h62 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9830; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11241 = 7'h63 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9831; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11242 = 7'h64 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9832; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11243 = 7'h65 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9833; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11244 = 7'h66 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9834; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11245 = 7'h67 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9835; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11246 = 7'h68 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9836; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11247 = 7'h69 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9837; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11248 = 7'h6a == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9838; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11249 = 7'h6b == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9839; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11250 = 7'h6c == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9840; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11251 = 7'h6d == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9841; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11252 = 7'h6e == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9842; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11253 = 7'h6f == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9843; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11254 = 7'h70 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9844; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11255 = 7'h71 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9845; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11256 = 7'h72 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9846; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11257 = 7'h73 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9847; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11258 = 7'h74 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9848; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11259 = 7'h75 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9849; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11260 = 7'h76 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9850; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11261 = 7'h77 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9851; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11262 = 7'h78 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9852; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11263 = 7'h79 == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9853; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11264 = 7'h7a == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9854; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11265 = 7'h7b == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9855; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11266 = 7'h7c == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9856; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11267 = 7'h7d == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9857; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11268 = 7'h7e == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9858; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_11269 = 7'h7f == out_payload_1_rob_idx[6:0] ? _rob_flits_returned_T_5 : _GEN_9859; // @[TestHarness.scala 213:{35,35}]
  wire [15:0] _rob_payload_flits_fired_T_5 = _GEN_10373 + 16'h1; // @[TestHarness.scala 214:76]
  wire [15:0] _GEN_11398 = 7'h0 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9860; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11399 = 7'h1 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9861; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11400 = 7'h2 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9862; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11401 = 7'h3 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9863; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11402 = 7'h4 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9864; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11403 = 7'h5 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9865; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11404 = 7'h6 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9866; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11405 = 7'h7 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9867; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11406 = 7'h8 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9868; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11407 = 7'h9 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9869; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11408 = 7'ha == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9870; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11409 = 7'hb == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9871; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11410 = 7'hc == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9872; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11411 = 7'hd == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9873; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11412 = 7'he == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9874; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11413 = 7'hf == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9875; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11414 = 7'h10 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9876; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11415 = 7'h11 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9877; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11416 = 7'h12 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9878; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11417 = 7'h13 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9879; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11418 = 7'h14 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9880; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11419 = 7'h15 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9881; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11420 = 7'h16 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9882; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11421 = 7'h17 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9883; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11422 = 7'h18 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9884; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11423 = 7'h19 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9885; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11424 = 7'h1a == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9886; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11425 = 7'h1b == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9887; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11426 = 7'h1c == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9888; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11427 = 7'h1d == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9889; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11428 = 7'h1e == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9890; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11429 = 7'h1f == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9891; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11430 = 7'h20 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9892; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11431 = 7'h21 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9893; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11432 = 7'h22 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9894; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11433 = 7'h23 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9895; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11434 = 7'h24 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9896; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11435 = 7'h25 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9897; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11436 = 7'h26 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9898; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11437 = 7'h27 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9899; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11438 = 7'h28 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9900; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11439 = 7'h29 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9901; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11440 = 7'h2a == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9902; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11441 = 7'h2b == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9903; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11442 = 7'h2c == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9904; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11443 = 7'h2d == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9905; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11444 = 7'h2e == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9906; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11445 = 7'h2f == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9907; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11446 = 7'h30 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9908; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11447 = 7'h31 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9909; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11448 = 7'h32 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9910; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11449 = 7'h33 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9911; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11450 = 7'h34 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9912; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11451 = 7'h35 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9913; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11452 = 7'h36 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9914; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11453 = 7'h37 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9915; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11454 = 7'h38 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9916; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11455 = 7'h39 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9917; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11456 = 7'h3a == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9918; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11457 = 7'h3b == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9919; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11458 = 7'h3c == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9920; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11459 = 7'h3d == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9921; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11460 = 7'h3e == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9922; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11461 = 7'h3f == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9923; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11462 = 7'h40 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9924; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11463 = 7'h41 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9925; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11464 = 7'h42 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9926; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11465 = 7'h43 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9927; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11466 = 7'h44 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9928; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11467 = 7'h45 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9929; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11468 = 7'h46 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9930; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11469 = 7'h47 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9931; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11470 = 7'h48 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9932; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11471 = 7'h49 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9933; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11472 = 7'h4a == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9934; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11473 = 7'h4b == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9935; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11474 = 7'h4c == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9936; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11475 = 7'h4d == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9937; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11476 = 7'h4e == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9938; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11477 = 7'h4f == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9939; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11478 = 7'h50 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9940; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11479 = 7'h51 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9941; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11480 = 7'h52 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9942; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11481 = 7'h53 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9943; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11482 = 7'h54 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9944; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11483 = 7'h55 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9945; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11484 = 7'h56 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9946; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11485 = 7'h57 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9947; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11486 = 7'h58 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9948; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11487 = 7'h59 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9949; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11488 = 7'h5a == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9950; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11489 = 7'h5b == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9951; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11490 = 7'h5c == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9952; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11491 = 7'h5d == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9953; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11492 = 7'h5e == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9954; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11493 = 7'h5f == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9955; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11494 = 7'h60 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9956; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11495 = 7'h61 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9957; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11496 = 7'h62 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9958; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11497 = 7'h63 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9959; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11498 = 7'h64 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9960; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11499 = 7'h65 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9961; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11500 = 7'h66 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9962; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11501 = 7'h67 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9963; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11502 = 7'h68 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9964; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11503 = 7'h69 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9965; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11504 = 7'h6a == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9966; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11505 = 7'h6b == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9967; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11506 = 7'h6c == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9968; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11507 = 7'h6d == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9969; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11508 = 7'h6e == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9970; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11509 = 7'h6f == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9971; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11510 = 7'h70 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9972; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11511 = 7'h71 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9973; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11512 = 7'h72 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9974; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11513 = 7'h73 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9975; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11514 = 7'h74 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9976; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11515 = 7'h75 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9977; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11516 = 7'h76 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9978; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11517 = 7'h77 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9979; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11518 = 7'h78 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9980; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11519 = 7'h79 == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9981; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11520 = 7'h7a == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9982; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11521 = 7'h7b == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9983; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11522 = 7'h7c == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9984; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11523 = 7'h7d == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9985; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11524 = 7'h7e == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9986; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_11525 = 7'h7f == out_payload_1_rob_idx[6:0] ? _rob_payload_flits_fired_T_5 : _GEN_9987; // @[TestHarness.scala 214:{40,40}]
  wire  _GEN_11526 = io_from_noc_1_flit_bits_head | packet_valid_1; // @[TestHarness.scala 196:31 215:{31,46}]
  wire [15:0] _GEN_11527 = io_from_noc_1_flit_bits_head ? out_payload_1_rob_idx : {{9'd0}, packet_rob_idx_1}; // @[TestHarness.scala 197:29 215:{31,72}]
  wire [3:0] _GEN_11529 = _T_165 ? _GEN_11142 : _GEN_9732; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11530 = _T_165 ? _GEN_11143 : _GEN_9733; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11531 = _T_165 ? _GEN_11144 : _GEN_9734; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11532 = _T_165 ? _GEN_11145 : _GEN_9735; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11533 = _T_165 ? _GEN_11146 : _GEN_9736; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11534 = _T_165 ? _GEN_11147 : _GEN_9737; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11535 = _T_165 ? _GEN_11148 : _GEN_9738; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11536 = _T_165 ? _GEN_11149 : _GEN_9739; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11537 = _T_165 ? _GEN_11150 : _GEN_9740; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11538 = _T_165 ? _GEN_11151 : _GEN_9741; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11539 = _T_165 ? _GEN_11152 : _GEN_9742; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11540 = _T_165 ? _GEN_11153 : _GEN_9743; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11541 = _T_165 ? _GEN_11154 : _GEN_9744; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11542 = _T_165 ? _GEN_11155 : _GEN_9745; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11543 = _T_165 ? _GEN_11156 : _GEN_9746; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11544 = _T_165 ? _GEN_11157 : _GEN_9747; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11545 = _T_165 ? _GEN_11158 : _GEN_9748; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11546 = _T_165 ? _GEN_11159 : _GEN_9749; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11547 = _T_165 ? _GEN_11160 : _GEN_9750; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11548 = _T_165 ? _GEN_11161 : _GEN_9751; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11549 = _T_165 ? _GEN_11162 : _GEN_9752; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11550 = _T_165 ? _GEN_11163 : _GEN_9753; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11551 = _T_165 ? _GEN_11164 : _GEN_9754; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11552 = _T_165 ? _GEN_11165 : _GEN_9755; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11553 = _T_165 ? _GEN_11166 : _GEN_9756; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11554 = _T_165 ? _GEN_11167 : _GEN_9757; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11555 = _T_165 ? _GEN_11168 : _GEN_9758; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11556 = _T_165 ? _GEN_11169 : _GEN_9759; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11557 = _T_165 ? _GEN_11170 : _GEN_9760; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11558 = _T_165 ? _GEN_11171 : _GEN_9761; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11559 = _T_165 ? _GEN_11172 : _GEN_9762; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11560 = _T_165 ? _GEN_11173 : _GEN_9763; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11561 = _T_165 ? _GEN_11174 : _GEN_9764; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11562 = _T_165 ? _GEN_11175 : _GEN_9765; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11563 = _T_165 ? _GEN_11176 : _GEN_9766; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11564 = _T_165 ? _GEN_11177 : _GEN_9767; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11565 = _T_165 ? _GEN_11178 : _GEN_9768; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11566 = _T_165 ? _GEN_11179 : _GEN_9769; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11567 = _T_165 ? _GEN_11180 : _GEN_9770; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11568 = _T_165 ? _GEN_11181 : _GEN_9771; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11569 = _T_165 ? _GEN_11182 : _GEN_9772; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11570 = _T_165 ? _GEN_11183 : _GEN_9773; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11571 = _T_165 ? _GEN_11184 : _GEN_9774; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11572 = _T_165 ? _GEN_11185 : _GEN_9775; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11573 = _T_165 ? _GEN_11186 : _GEN_9776; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11574 = _T_165 ? _GEN_11187 : _GEN_9777; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11575 = _T_165 ? _GEN_11188 : _GEN_9778; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11576 = _T_165 ? _GEN_11189 : _GEN_9779; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11577 = _T_165 ? _GEN_11190 : _GEN_9780; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11578 = _T_165 ? _GEN_11191 : _GEN_9781; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11579 = _T_165 ? _GEN_11192 : _GEN_9782; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11580 = _T_165 ? _GEN_11193 : _GEN_9783; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11581 = _T_165 ? _GEN_11194 : _GEN_9784; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11582 = _T_165 ? _GEN_11195 : _GEN_9785; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11583 = _T_165 ? _GEN_11196 : _GEN_9786; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11584 = _T_165 ? _GEN_11197 : _GEN_9787; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11585 = _T_165 ? _GEN_11198 : _GEN_9788; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11586 = _T_165 ? _GEN_11199 : _GEN_9789; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11587 = _T_165 ? _GEN_11200 : _GEN_9790; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11588 = _T_165 ? _GEN_11201 : _GEN_9791; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11589 = _T_165 ? _GEN_11202 : _GEN_9792; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11590 = _T_165 ? _GEN_11203 : _GEN_9793; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11591 = _T_165 ? _GEN_11204 : _GEN_9794; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11592 = _T_165 ? _GEN_11205 : _GEN_9795; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11593 = _T_165 ? _GEN_11206 : _GEN_9796; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11594 = _T_165 ? _GEN_11207 : _GEN_9797; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11595 = _T_165 ? _GEN_11208 : _GEN_9798; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11596 = _T_165 ? _GEN_11209 : _GEN_9799; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11597 = _T_165 ? _GEN_11210 : _GEN_9800; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11598 = _T_165 ? _GEN_11211 : _GEN_9801; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11599 = _T_165 ? _GEN_11212 : _GEN_9802; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11600 = _T_165 ? _GEN_11213 : _GEN_9803; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11601 = _T_165 ? _GEN_11214 : _GEN_9804; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11602 = _T_165 ? _GEN_11215 : _GEN_9805; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11603 = _T_165 ? _GEN_11216 : _GEN_9806; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11604 = _T_165 ? _GEN_11217 : _GEN_9807; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11605 = _T_165 ? _GEN_11218 : _GEN_9808; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11606 = _T_165 ? _GEN_11219 : _GEN_9809; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11607 = _T_165 ? _GEN_11220 : _GEN_9810; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11608 = _T_165 ? _GEN_11221 : _GEN_9811; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11609 = _T_165 ? _GEN_11222 : _GEN_9812; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11610 = _T_165 ? _GEN_11223 : _GEN_9813; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11611 = _T_165 ? _GEN_11224 : _GEN_9814; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11612 = _T_165 ? _GEN_11225 : _GEN_9815; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11613 = _T_165 ? _GEN_11226 : _GEN_9816; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11614 = _T_165 ? _GEN_11227 : _GEN_9817; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11615 = _T_165 ? _GEN_11228 : _GEN_9818; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11616 = _T_165 ? _GEN_11229 : _GEN_9819; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11617 = _T_165 ? _GEN_11230 : _GEN_9820; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11618 = _T_165 ? _GEN_11231 : _GEN_9821; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11619 = _T_165 ? _GEN_11232 : _GEN_9822; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11620 = _T_165 ? _GEN_11233 : _GEN_9823; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11621 = _T_165 ? _GEN_11234 : _GEN_9824; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11622 = _T_165 ? _GEN_11235 : _GEN_9825; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11623 = _T_165 ? _GEN_11236 : _GEN_9826; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11624 = _T_165 ? _GEN_11237 : _GEN_9827; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11625 = _T_165 ? _GEN_11238 : _GEN_9828; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11626 = _T_165 ? _GEN_11239 : _GEN_9829; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11627 = _T_165 ? _GEN_11240 : _GEN_9830; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11628 = _T_165 ? _GEN_11241 : _GEN_9831; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11629 = _T_165 ? _GEN_11242 : _GEN_9832; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11630 = _T_165 ? _GEN_11243 : _GEN_9833; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11631 = _T_165 ? _GEN_11244 : _GEN_9834; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11632 = _T_165 ? _GEN_11245 : _GEN_9835; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11633 = _T_165 ? _GEN_11246 : _GEN_9836; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11634 = _T_165 ? _GEN_11247 : _GEN_9837; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11635 = _T_165 ? _GEN_11248 : _GEN_9838; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11636 = _T_165 ? _GEN_11249 : _GEN_9839; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11637 = _T_165 ? _GEN_11250 : _GEN_9840; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11638 = _T_165 ? _GEN_11251 : _GEN_9841; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11639 = _T_165 ? _GEN_11252 : _GEN_9842; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11640 = _T_165 ? _GEN_11253 : _GEN_9843; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11641 = _T_165 ? _GEN_11254 : _GEN_9844; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11642 = _T_165 ? _GEN_11255 : _GEN_9845; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11643 = _T_165 ? _GEN_11256 : _GEN_9846; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11644 = _T_165 ? _GEN_11257 : _GEN_9847; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11645 = _T_165 ? _GEN_11258 : _GEN_9848; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11646 = _T_165 ? _GEN_11259 : _GEN_9849; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11647 = _T_165 ? _GEN_11260 : _GEN_9850; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11648 = _T_165 ? _GEN_11261 : _GEN_9851; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11649 = _T_165 ? _GEN_11262 : _GEN_9852; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11650 = _T_165 ? _GEN_11263 : _GEN_9853; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11651 = _T_165 ? _GEN_11264 : _GEN_9854; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11652 = _T_165 ? _GEN_11265 : _GEN_9855; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11653 = _T_165 ? _GEN_11266 : _GEN_9856; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11654 = _T_165 ? _GEN_11267 : _GEN_9857; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11655 = _T_165 ? _GEN_11268 : _GEN_9858; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_11656 = _T_165 ? _GEN_11269 : _GEN_9859; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11657 = _T_165 ? _GEN_11398 : _GEN_9860; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11658 = _T_165 ? _GEN_11399 : _GEN_9861; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11659 = _T_165 ? _GEN_11400 : _GEN_9862; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11660 = _T_165 ? _GEN_11401 : _GEN_9863; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11661 = _T_165 ? _GEN_11402 : _GEN_9864; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11662 = _T_165 ? _GEN_11403 : _GEN_9865; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11663 = _T_165 ? _GEN_11404 : _GEN_9866; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11664 = _T_165 ? _GEN_11405 : _GEN_9867; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11665 = _T_165 ? _GEN_11406 : _GEN_9868; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11666 = _T_165 ? _GEN_11407 : _GEN_9869; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11667 = _T_165 ? _GEN_11408 : _GEN_9870; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11668 = _T_165 ? _GEN_11409 : _GEN_9871; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11669 = _T_165 ? _GEN_11410 : _GEN_9872; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11670 = _T_165 ? _GEN_11411 : _GEN_9873; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11671 = _T_165 ? _GEN_11412 : _GEN_9874; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11672 = _T_165 ? _GEN_11413 : _GEN_9875; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11673 = _T_165 ? _GEN_11414 : _GEN_9876; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11674 = _T_165 ? _GEN_11415 : _GEN_9877; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11675 = _T_165 ? _GEN_11416 : _GEN_9878; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11676 = _T_165 ? _GEN_11417 : _GEN_9879; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11677 = _T_165 ? _GEN_11418 : _GEN_9880; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11678 = _T_165 ? _GEN_11419 : _GEN_9881; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11679 = _T_165 ? _GEN_11420 : _GEN_9882; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11680 = _T_165 ? _GEN_11421 : _GEN_9883; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11681 = _T_165 ? _GEN_11422 : _GEN_9884; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11682 = _T_165 ? _GEN_11423 : _GEN_9885; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11683 = _T_165 ? _GEN_11424 : _GEN_9886; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11684 = _T_165 ? _GEN_11425 : _GEN_9887; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11685 = _T_165 ? _GEN_11426 : _GEN_9888; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11686 = _T_165 ? _GEN_11427 : _GEN_9889; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11687 = _T_165 ? _GEN_11428 : _GEN_9890; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11688 = _T_165 ? _GEN_11429 : _GEN_9891; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11689 = _T_165 ? _GEN_11430 : _GEN_9892; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11690 = _T_165 ? _GEN_11431 : _GEN_9893; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11691 = _T_165 ? _GEN_11432 : _GEN_9894; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11692 = _T_165 ? _GEN_11433 : _GEN_9895; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11693 = _T_165 ? _GEN_11434 : _GEN_9896; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11694 = _T_165 ? _GEN_11435 : _GEN_9897; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11695 = _T_165 ? _GEN_11436 : _GEN_9898; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11696 = _T_165 ? _GEN_11437 : _GEN_9899; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11697 = _T_165 ? _GEN_11438 : _GEN_9900; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11698 = _T_165 ? _GEN_11439 : _GEN_9901; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11699 = _T_165 ? _GEN_11440 : _GEN_9902; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11700 = _T_165 ? _GEN_11441 : _GEN_9903; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11701 = _T_165 ? _GEN_11442 : _GEN_9904; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11702 = _T_165 ? _GEN_11443 : _GEN_9905; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11703 = _T_165 ? _GEN_11444 : _GEN_9906; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11704 = _T_165 ? _GEN_11445 : _GEN_9907; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11705 = _T_165 ? _GEN_11446 : _GEN_9908; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11706 = _T_165 ? _GEN_11447 : _GEN_9909; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11707 = _T_165 ? _GEN_11448 : _GEN_9910; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11708 = _T_165 ? _GEN_11449 : _GEN_9911; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11709 = _T_165 ? _GEN_11450 : _GEN_9912; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11710 = _T_165 ? _GEN_11451 : _GEN_9913; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11711 = _T_165 ? _GEN_11452 : _GEN_9914; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11712 = _T_165 ? _GEN_11453 : _GEN_9915; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11713 = _T_165 ? _GEN_11454 : _GEN_9916; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11714 = _T_165 ? _GEN_11455 : _GEN_9917; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11715 = _T_165 ? _GEN_11456 : _GEN_9918; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11716 = _T_165 ? _GEN_11457 : _GEN_9919; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11717 = _T_165 ? _GEN_11458 : _GEN_9920; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11718 = _T_165 ? _GEN_11459 : _GEN_9921; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11719 = _T_165 ? _GEN_11460 : _GEN_9922; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11720 = _T_165 ? _GEN_11461 : _GEN_9923; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11721 = _T_165 ? _GEN_11462 : _GEN_9924; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11722 = _T_165 ? _GEN_11463 : _GEN_9925; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11723 = _T_165 ? _GEN_11464 : _GEN_9926; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11724 = _T_165 ? _GEN_11465 : _GEN_9927; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11725 = _T_165 ? _GEN_11466 : _GEN_9928; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11726 = _T_165 ? _GEN_11467 : _GEN_9929; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11727 = _T_165 ? _GEN_11468 : _GEN_9930; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11728 = _T_165 ? _GEN_11469 : _GEN_9931; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11729 = _T_165 ? _GEN_11470 : _GEN_9932; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11730 = _T_165 ? _GEN_11471 : _GEN_9933; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11731 = _T_165 ? _GEN_11472 : _GEN_9934; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11732 = _T_165 ? _GEN_11473 : _GEN_9935; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11733 = _T_165 ? _GEN_11474 : _GEN_9936; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11734 = _T_165 ? _GEN_11475 : _GEN_9937; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11735 = _T_165 ? _GEN_11476 : _GEN_9938; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11736 = _T_165 ? _GEN_11477 : _GEN_9939; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11737 = _T_165 ? _GEN_11478 : _GEN_9940; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11738 = _T_165 ? _GEN_11479 : _GEN_9941; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11739 = _T_165 ? _GEN_11480 : _GEN_9942; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11740 = _T_165 ? _GEN_11481 : _GEN_9943; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11741 = _T_165 ? _GEN_11482 : _GEN_9944; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11742 = _T_165 ? _GEN_11483 : _GEN_9945; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11743 = _T_165 ? _GEN_11484 : _GEN_9946; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11744 = _T_165 ? _GEN_11485 : _GEN_9947; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11745 = _T_165 ? _GEN_11486 : _GEN_9948; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11746 = _T_165 ? _GEN_11487 : _GEN_9949; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11747 = _T_165 ? _GEN_11488 : _GEN_9950; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11748 = _T_165 ? _GEN_11489 : _GEN_9951; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11749 = _T_165 ? _GEN_11490 : _GEN_9952; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11750 = _T_165 ? _GEN_11491 : _GEN_9953; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11751 = _T_165 ? _GEN_11492 : _GEN_9954; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11752 = _T_165 ? _GEN_11493 : _GEN_9955; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11753 = _T_165 ? _GEN_11494 : _GEN_9956; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11754 = _T_165 ? _GEN_11495 : _GEN_9957; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11755 = _T_165 ? _GEN_11496 : _GEN_9958; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11756 = _T_165 ? _GEN_11497 : _GEN_9959; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11757 = _T_165 ? _GEN_11498 : _GEN_9960; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11758 = _T_165 ? _GEN_11499 : _GEN_9961; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11759 = _T_165 ? _GEN_11500 : _GEN_9962; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11760 = _T_165 ? _GEN_11501 : _GEN_9963; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11761 = _T_165 ? _GEN_11502 : _GEN_9964; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11762 = _T_165 ? _GEN_11503 : _GEN_9965; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11763 = _T_165 ? _GEN_11504 : _GEN_9966; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11764 = _T_165 ? _GEN_11505 : _GEN_9967; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11765 = _T_165 ? _GEN_11506 : _GEN_9968; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11766 = _T_165 ? _GEN_11507 : _GEN_9969; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11767 = _T_165 ? _GEN_11508 : _GEN_9970; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11768 = _T_165 ? _GEN_11509 : _GEN_9971; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11769 = _T_165 ? _GEN_11510 : _GEN_9972; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11770 = _T_165 ? _GEN_11511 : _GEN_9973; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11771 = _T_165 ? _GEN_11512 : _GEN_9974; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11772 = _T_165 ? _GEN_11513 : _GEN_9975; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11773 = _T_165 ? _GEN_11514 : _GEN_9976; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11774 = _T_165 ? _GEN_11515 : _GEN_9977; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11775 = _T_165 ? _GEN_11516 : _GEN_9978; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11776 = _T_165 ? _GEN_11517 : _GEN_9979; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11777 = _T_165 ? _GEN_11518 : _GEN_9980; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11778 = _T_165 ? _GEN_11519 : _GEN_9981; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11779 = _T_165 ? _GEN_11520 : _GEN_9982; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11780 = _T_165 ? _GEN_11521 : _GEN_9983; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11781 = _T_165 ? _GEN_11522 : _GEN_9984; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11782 = _T_165 ? _GEN_11523 : _GEN_9985; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11783 = _T_165 ? _GEN_11524 : _GEN_9986; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11784 = _T_165 ? _GEN_11525 : _GEN_9987; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_11786 = _T_165 ? _GEN_11527 : {{9'd0}, packet_rob_idx_1}; // @[TestHarness.scala 199:26 197:29]
  wire [31:0] out_payload_2_tsc = io_from_noc_2_flit_bits_payload[63:32]; // @[TestHarness.scala 194:51]
  reg  packet_valid_2; // @[TestHarness.scala 196:31]
  reg [6:0] packet_rob_idx_2; // @[TestHarness.scala 197:29]
  wire [127:0] _T_170 = rob_valids >> out_payload_2_rob_idx; // @[TestHarness.scala 201:24]
  wire [31:0] _GEN_11788 = 7'h1 == out_payload_2_rob_idx[6:0] ? rob_payload_1_tsc : rob_payload_0_tsc; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11789 = 7'h2 == out_payload_2_rob_idx[6:0] ? rob_payload_2_tsc : _GEN_11788; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11790 = 7'h3 == out_payload_2_rob_idx[6:0] ? rob_payload_3_tsc : _GEN_11789; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11791 = 7'h4 == out_payload_2_rob_idx[6:0] ? rob_payload_4_tsc : _GEN_11790; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11792 = 7'h5 == out_payload_2_rob_idx[6:0] ? rob_payload_5_tsc : _GEN_11791; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11793 = 7'h6 == out_payload_2_rob_idx[6:0] ? rob_payload_6_tsc : _GEN_11792; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11794 = 7'h7 == out_payload_2_rob_idx[6:0] ? rob_payload_7_tsc : _GEN_11793; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11795 = 7'h8 == out_payload_2_rob_idx[6:0] ? rob_payload_8_tsc : _GEN_11794; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11796 = 7'h9 == out_payload_2_rob_idx[6:0] ? rob_payload_9_tsc : _GEN_11795; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11797 = 7'ha == out_payload_2_rob_idx[6:0] ? rob_payload_10_tsc : _GEN_11796; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11798 = 7'hb == out_payload_2_rob_idx[6:0] ? rob_payload_11_tsc : _GEN_11797; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11799 = 7'hc == out_payload_2_rob_idx[6:0] ? rob_payload_12_tsc : _GEN_11798; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11800 = 7'hd == out_payload_2_rob_idx[6:0] ? rob_payload_13_tsc : _GEN_11799; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11801 = 7'he == out_payload_2_rob_idx[6:0] ? rob_payload_14_tsc : _GEN_11800; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11802 = 7'hf == out_payload_2_rob_idx[6:0] ? rob_payload_15_tsc : _GEN_11801; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11803 = 7'h10 == out_payload_2_rob_idx[6:0] ? rob_payload_16_tsc : _GEN_11802; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11804 = 7'h11 == out_payload_2_rob_idx[6:0] ? rob_payload_17_tsc : _GEN_11803; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11805 = 7'h12 == out_payload_2_rob_idx[6:0] ? rob_payload_18_tsc : _GEN_11804; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11806 = 7'h13 == out_payload_2_rob_idx[6:0] ? rob_payload_19_tsc : _GEN_11805; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11807 = 7'h14 == out_payload_2_rob_idx[6:0] ? rob_payload_20_tsc : _GEN_11806; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11808 = 7'h15 == out_payload_2_rob_idx[6:0] ? rob_payload_21_tsc : _GEN_11807; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11809 = 7'h16 == out_payload_2_rob_idx[6:0] ? rob_payload_22_tsc : _GEN_11808; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11810 = 7'h17 == out_payload_2_rob_idx[6:0] ? rob_payload_23_tsc : _GEN_11809; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11811 = 7'h18 == out_payload_2_rob_idx[6:0] ? rob_payload_24_tsc : _GEN_11810; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11812 = 7'h19 == out_payload_2_rob_idx[6:0] ? rob_payload_25_tsc : _GEN_11811; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11813 = 7'h1a == out_payload_2_rob_idx[6:0] ? rob_payload_26_tsc : _GEN_11812; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11814 = 7'h1b == out_payload_2_rob_idx[6:0] ? rob_payload_27_tsc : _GEN_11813; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11815 = 7'h1c == out_payload_2_rob_idx[6:0] ? rob_payload_28_tsc : _GEN_11814; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11816 = 7'h1d == out_payload_2_rob_idx[6:0] ? rob_payload_29_tsc : _GEN_11815; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11817 = 7'h1e == out_payload_2_rob_idx[6:0] ? rob_payload_30_tsc : _GEN_11816; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11818 = 7'h1f == out_payload_2_rob_idx[6:0] ? rob_payload_31_tsc : _GEN_11817; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11819 = 7'h20 == out_payload_2_rob_idx[6:0] ? rob_payload_32_tsc : _GEN_11818; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11820 = 7'h21 == out_payload_2_rob_idx[6:0] ? rob_payload_33_tsc : _GEN_11819; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11821 = 7'h22 == out_payload_2_rob_idx[6:0] ? rob_payload_34_tsc : _GEN_11820; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11822 = 7'h23 == out_payload_2_rob_idx[6:0] ? rob_payload_35_tsc : _GEN_11821; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11823 = 7'h24 == out_payload_2_rob_idx[6:0] ? rob_payload_36_tsc : _GEN_11822; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11824 = 7'h25 == out_payload_2_rob_idx[6:0] ? rob_payload_37_tsc : _GEN_11823; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11825 = 7'h26 == out_payload_2_rob_idx[6:0] ? rob_payload_38_tsc : _GEN_11824; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11826 = 7'h27 == out_payload_2_rob_idx[6:0] ? rob_payload_39_tsc : _GEN_11825; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11827 = 7'h28 == out_payload_2_rob_idx[6:0] ? rob_payload_40_tsc : _GEN_11826; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11828 = 7'h29 == out_payload_2_rob_idx[6:0] ? rob_payload_41_tsc : _GEN_11827; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11829 = 7'h2a == out_payload_2_rob_idx[6:0] ? rob_payload_42_tsc : _GEN_11828; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11830 = 7'h2b == out_payload_2_rob_idx[6:0] ? rob_payload_43_tsc : _GEN_11829; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11831 = 7'h2c == out_payload_2_rob_idx[6:0] ? rob_payload_44_tsc : _GEN_11830; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11832 = 7'h2d == out_payload_2_rob_idx[6:0] ? rob_payload_45_tsc : _GEN_11831; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11833 = 7'h2e == out_payload_2_rob_idx[6:0] ? rob_payload_46_tsc : _GEN_11832; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11834 = 7'h2f == out_payload_2_rob_idx[6:0] ? rob_payload_47_tsc : _GEN_11833; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11835 = 7'h30 == out_payload_2_rob_idx[6:0] ? rob_payload_48_tsc : _GEN_11834; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11836 = 7'h31 == out_payload_2_rob_idx[6:0] ? rob_payload_49_tsc : _GEN_11835; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11837 = 7'h32 == out_payload_2_rob_idx[6:0] ? rob_payload_50_tsc : _GEN_11836; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11838 = 7'h33 == out_payload_2_rob_idx[6:0] ? rob_payload_51_tsc : _GEN_11837; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11839 = 7'h34 == out_payload_2_rob_idx[6:0] ? rob_payload_52_tsc : _GEN_11838; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11840 = 7'h35 == out_payload_2_rob_idx[6:0] ? rob_payload_53_tsc : _GEN_11839; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11841 = 7'h36 == out_payload_2_rob_idx[6:0] ? rob_payload_54_tsc : _GEN_11840; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11842 = 7'h37 == out_payload_2_rob_idx[6:0] ? rob_payload_55_tsc : _GEN_11841; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11843 = 7'h38 == out_payload_2_rob_idx[6:0] ? rob_payload_56_tsc : _GEN_11842; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11844 = 7'h39 == out_payload_2_rob_idx[6:0] ? rob_payload_57_tsc : _GEN_11843; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11845 = 7'h3a == out_payload_2_rob_idx[6:0] ? rob_payload_58_tsc : _GEN_11844; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11846 = 7'h3b == out_payload_2_rob_idx[6:0] ? rob_payload_59_tsc : _GEN_11845; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11847 = 7'h3c == out_payload_2_rob_idx[6:0] ? rob_payload_60_tsc : _GEN_11846; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11848 = 7'h3d == out_payload_2_rob_idx[6:0] ? rob_payload_61_tsc : _GEN_11847; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11849 = 7'h3e == out_payload_2_rob_idx[6:0] ? rob_payload_62_tsc : _GEN_11848; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11850 = 7'h3f == out_payload_2_rob_idx[6:0] ? rob_payload_63_tsc : _GEN_11849; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11851 = 7'h40 == out_payload_2_rob_idx[6:0] ? rob_payload_64_tsc : _GEN_11850; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11852 = 7'h41 == out_payload_2_rob_idx[6:0] ? rob_payload_65_tsc : _GEN_11851; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11853 = 7'h42 == out_payload_2_rob_idx[6:0] ? rob_payload_66_tsc : _GEN_11852; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11854 = 7'h43 == out_payload_2_rob_idx[6:0] ? rob_payload_67_tsc : _GEN_11853; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11855 = 7'h44 == out_payload_2_rob_idx[6:0] ? rob_payload_68_tsc : _GEN_11854; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11856 = 7'h45 == out_payload_2_rob_idx[6:0] ? rob_payload_69_tsc : _GEN_11855; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11857 = 7'h46 == out_payload_2_rob_idx[6:0] ? rob_payload_70_tsc : _GEN_11856; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11858 = 7'h47 == out_payload_2_rob_idx[6:0] ? rob_payload_71_tsc : _GEN_11857; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11859 = 7'h48 == out_payload_2_rob_idx[6:0] ? rob_payload_72_tsc : _GEN_11858; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11860 = 7'h49 == out_payload_2_rob_idx[6:0] ? rob_payload_73_tsc : _GEN_11859; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11861 = 7'h4a == out_payload_2_rob_idx[6:0] ? rob_payload_74_tsc : _GEN_11860; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11862 = 7'h4b == out_payload_2_rob_idx[6:0] ? rob_payload_75_tsc : _GEN_11861; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11863 = 7'h4c == out_payload_2_rob_idx[6:0] ? rob_payload_76_tsc : _GEN_11862; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11864 = 7'h4d == out_payload_2_rob_idx[6:0] ? rob_payload_77_tsc : _GEN_11863; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11865 = 7'h4e == out_payload_2_rob_idx[6:0] ? rob_payload_78_tsc : _GEN_11864; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11866 = 7'h4f == out_payload_2_rob_idx[6:0] ? rob_payload_79_tsc : _GEN_11865; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11867 = 7'h50 == out_payload_2_rob_idx[6:0] ? rob_payload_80_tsc : _GEN_11866; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11868 = 7'h51 == out_payload_2_rob_idx[6:0] ? rob_payload_81_tsc : _GEN_11867; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11869 = 7'h52 == out_payload_2_rob_idx[6:0] ? rob_payload_82_tsc : _GEN_11868; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11870 = 7'h53 == out_payload_2_rob_idx[6:0] ? rob_payload_83_tsc : _GEN_11869; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11871 = 7'h54 == out_payload_2_rob_idx[6:0] ? rob_payload_84_tsc : _GEN_11870; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11872 = 7'h55 == out_payload_2_rob_idx[6:0] ? rob_payload_85_tsc : _GEN_11871; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11873 = 7'h56 == out_payload_2_rob_idx[6:0] ? rob_payload_86_tsc : _GEN_11872; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11874 = 7'h57 == out_payload_2_rob_idx[6:0] ? rob_payload_87_tsc : _GEN_11873; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11875 = 7'h58 == out_payload_2_rob_idx[6:0] ? rob_payload_88_tsc : _GEN_11874; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11876 = 7'h59 == out_payload_2_rob_idx[6:0] ? rob_payload_89_tsc : _GEN_11875; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11877 = 7'h5a == out_payload_2_rob_idx[6:0] ? rob_payload_90_tsc : _GEN_11876; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11878 = 7'h5b == out_payload_2_rob_idx[6:0] ? rob_payload_91_tsc : _GEN_11877; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11879 = 7'h5c == out_payload_2_rob_idx[6:0] ? rob_payload_92_tsc : _GEN_11878; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11880 = 7'h5d == out_payload_2_rob_idx[6:0] ? rob_payload_93_tsc : _GEN_11879; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11881 = 7'h5e == out_payload_2_rob_idx[6:0] ? rob_payload_94_tsc : _GEN_11880; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11882 = 7'h5f == out_payload_2_rob_idx[6:0] ? rob_payload_95_tsc : _GEN_11881; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11883 = 7'h60 == out_payload_2_rob_idx[6:0] ? rob_payload_96_tsc : _GEN_11882; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11884 = 7'h61 == out_payload_2_rob_idx[6:0] ? rob_payload_97_tsc : _GEN_11883; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11885 = 7'h62 == out_payload_2_rob_idx[6:0] ? rob_payload_98_tsc : _GEN_11884; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11886 = 7'h63 == out_payload_2_rob_idx[6:0] ? rob_payload_99_tsc : _GEN_11885; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11887 = 7'h64 == out_payload_2_rob_idx[6:0] ? rob_payload_100_tsc : _GEN_11886; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11888 = 7'h65 == out_payload_2_rob_idx[6:0] ? rob_payload_101_tsc : _GEN_11887; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11889 = 7'h66 == out_payload_2_rob_idx[6:0] ? rob_payload_102_tsc : _GEN_11888; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11890 = 7'h67 == out_payload_2_rob_idx[6:0] ? rob_payload_103_tsc : _GEN_11889; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11891 = 7'h68 == out_payload_2_rob_idx[6:0] ? rob_payload_104_tsc : _GEN_11890; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11892 = 7'h69 == out_payload_2_rob_idx[6:0] ? rob_payload_105_tsc : _GEN_11891; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11893 = 7'h6a == out_payload_2_rob_idx[6:0] ? rob_payload_106_tsc : _GEN_11892; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11894 = 7'h6b == out_payload_2_rob_idx[6:0] ? rob_payload_107_tsc : _GEN_11893; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11895 = 7'h6c == out_payload_2_rob_idx[6:0] ? rob_payload_108_tsc : _GEN_11894; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11896 = 7'h6d == out_payload_2_rob_idx[6:0] ? rob_payload_109_tsc : _GEN_11895; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11897 = 7'h6e == out_payload_2_rob_idx[6:0] ? rob_payload_110_tsc : _GEN_11896; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11898 = 7'h6f == out_payload_2_rob_idx[6:0] ? rob_payload_111_tsc : _GEN_11897; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11899 = 7'h70 == out_payload_2_rob_idx[6:0] ? rob_payload_112_tsc : _GEN_11898; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11900 = 7'h71 == out_payload_2_rob_idx[6:0] ? rob_payload_113_tsc : _GEN_11899; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11901 = 7'h72 == out_payload_2_rob_idx[6:0] ? rob_payload_114_tsc : _GEN_11900; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11902 = 7'h73 == out_payload_2_rob_idx[6:0] ? rob_payload_115_tsc : _GEN_11901; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11903 = 7'h74 == out_payload_2_rob_idx[6:0] ? rob_payload_116_tsc : _GEN_11902; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11904 = 7'h75 == out_payload_2_rob_idx[6:0] ? rob_payload_117_tsc : _GEN_11903; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11905 = 7'h76 == out_payload_2_rob_idx[6:0] ? rob_payload_118_tsc : _GEN_11904; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11906 = 7'h77 == out_payload_2_rob_idx[6:0] ? rob_payload_119_tsc : _GEN_11905; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11907 = 7'h78 == out_payload_2_rob_idx[6:0] ? rob_payload_120_tsc : _GEN_11906; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11908 = 7'h79 == out_payload_2_rob_idx[6:0] ? rob_payload_121_tsc : _GEN_11907; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11909 = 7'h7a == out_payload_2_rob_idx[6:0] ? rob_payload_122_tsc : _GEN_11908; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11910 = 7'h7b == out_payload_2_rob_idx[6:0] ? rob_payload_123_tsc : _GEN_11909; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11911 = 7'h7c == out_payload_2_rob_idx[6:0] ? rob_payload_124_tsc : _GEN_11910; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11912 = 7'h7d == out_payload_2_rob_idx[6:0] ? rob_payload_125_tsc : _GEN_11911; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11913 = 7'h7e == out_payload_2_rob_idx[6:0] ? rob_payload_126_tsc : _GEN_11912; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_11914 = 7'h7f == out_payload_2_rob_idx[6:0] ? rob_payload_127_tsc : _GEN_11913; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11916 = 7'h1 == out_payload_2_rob_idx[6:0] ? rob_payload_1_rob_idx : rob_payload_0_rob_idx; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11917 = 7'h2 == out_payload_2_rob_idx[6:0] ? rob_payload_2_rob_idx : _GEN_11916; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11918 = 7'h3 == out_payload_2_rob_idx[6:0] ? rob_payload_3_rob_idx : _GEN_11917; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11919 = 7'h4 == out_payload_2_rob_idx[6:0] ? rob_payload_4_rob_idx : _GEN_11918; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11920 = 7'h5 == out_payload_2_rob_idx[6:0] ? rob_payload_5_rob_idx : _GEN_11919; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11921 = 7'h6 == out_payload_2_rob_idx[6:0] ? rob_payload_6_rob_idx : _GEN_11920; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11922 = 7'h7 == out_payload_2_rob_idx[6:0] ? rob_payload_7_rob_idx : _GEN_11921; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11923 = 7'h8 == out_payload_2_rob_idx[6:0] ? rob_payload_8_rob_idx : _GEN_11922; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11924 = 7'h9 == out_payload_2_rob_idx[6:0] ? rob_payload_9_rob_idx : _GEN_11923; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11925 = 7'ha == out_payload_2_rob_idx[6:0] ? rob_payload_10_rob_idx : _GEN_11924; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11926 = 7'hb == out_payload_2_rob_idx[6:0] ? rob_payload_11_rob_idx : _GEN_11925; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11927 = 7'hc == out_payload_2_rob_idx[6:0] ? rob_payload_12_rob_idx : _GEN_11926; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11928 = 7'hd == out_payload_2_rob_idx[6:0] ? rob_payload_13_rob_idx : _GEN_11927; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11929 = 7'he == out_payload_2_rob_idx[6:0] ? rob_payload_14_rob_idx : _GEN_11928; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11930 = 7'hf == out_payload_2_rob_idx[6:0] ? rob_payload_15_rob_idx : _GEN_11929; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11931 = 7'h10 == out_payload_2_rob_idx[6:0] ? rob_payload_16_rob_idx : _GEN_11930; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11932 = 7'h11 == out_payload_2_rob_idx[6:0] ? rob_payload_17_rob_idx : _GEN_11931; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11933 = 7'h12 == out_payload_2_rob_idx[6:0] ? rob_payload_18_rob_idx : _GEN_11932; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11934 = 7'h13 == out_payload_2_rob_idx[6:0] ? rob_payload_19_rob_idx : _GEN_11933; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11935 = 7'h14 == out_payload_2_rob_idx[6:0] ? rob_payload_20_rob_idx : _GEN_11934; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11936 = 7'h15 == out_payload_2_rob_idx[6:0] ? rob_payload_21_rob_idx : _GEN_11935; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11937 = 7'h16 == out_payload_2_rob_idx[6:0] ? rob_payload_22_rob_idx : _GEN_11936; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11938 = 7'h17 == out_payload_2_rob_idx[6:0] ? rob_payload_23_rob_idx : _GEN_11937; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11939 = 7'h18 == out_payload_2_rob_idx[6:0] ? rob_payload_24_rob_idx : _GEN_11938; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11940 = 7'h19 == out_payload_2_rob_idx[6:0] ? rob_payload_25_rob_idx : _GEN_11939; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11941 = 7'h1a == out_payload_2_rob_idx[6:0] ? rob_payload_26_rob_idx : _GEN_11940; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11942 = 7'h1b == out_payload_2_rob_idx[6:0] ? rob_payload_27_rob_idx : _GEN_11941; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11943 = 7'h1c == out_payload_2_rob_idx[6:0] ? rob_payload_28_rob_idx : _GEN_11942; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11944 = 7'h1d == out_payload_2_rob_idx[6:0] ? rob_payload_29_rob_idx : _GEN_11943; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11945 = 7'h1e == out_payload_2_rob_idx[6:0] ? rob_payload_30_rob_idx : _GEN_11944; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11946 = 7'h1f == out_payload_2_rob_idx[6:0] ? rob_payload_31_rob_idx : _GEN_11945; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11947 = 7'h20 == out_payload_2_rob_idx[6:0] ? rob_payload_32_rob_idx : _GEN_11946; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11948 = 7'h21 == out_payload_2_rob_idx[6:0] ? rob_payload_33_rob_idx : _GEN_11947; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11949 = 7'h22 == out_payload_2_rob_idx[6:0] ? rob_payload_34_rob_idx : _GEN_11948; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11950 = 7'h23 == out_payload_2_rob_idx[6:0] ? rob_payload_35_rob_idx : _GEN_11949; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11951 = 7'h24 == out_payload_2_rob_idx[6:0] ? rob_payload_36_rob_idx : _GEN_11950; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11952 = 7'h25 == out_payload_2_rob_idx[6:0] ? rob_payload_37_rob_idx : _GEN_11951; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11953 = 7'h26 == out_payload_2_rob_idx[6:0] ? rob_payload_38_rob_idx : _GEN_11952; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11954 = 7'h27 == out_payload_2_rob_idx[6:0] ? rob_payload_39_rob_idx : _GEN_11953; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11955 = 7'h28 == out_payload_2_rob_idx[6:0] ? rob_payload_40_rob_idx : _GEN_11954; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11956 = 7'h29 == out_payload_2_rob_idx[6:0] ? rob_payload_41_rob_idx : _GEN_11955; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11957 = 7'h2a == out_payload_2_rob_idx[6:0] ? rob_payload_42_rob_idx : _GEN_11956; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11958 = 7'h2b == out_payload_2_rob_idx[6:0] ? rob_payload_43_rob_idx : _GEN_11957; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11959 = 7'h2c == out_payload_2_rob_idx[6:0] ? rob_payload_44_rob_idx : _GEN_11958; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11960 = 7'h2d == out_payload_2_rob_idx[6:0] ? rob_payload_45_rob_idx : _GEN_11959; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11961 = 7'h2e == out_payload_2_rob_idx[6:0] ? rob_payload_46_rob_idx : _GEN_11960; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11962 = 7'h2f == out_payload_2_rob_idx[6:0] ? rob_payload_47_rob_idx : _GEN_11961; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11963 = 7'h30 == out_payload_2_rob_idx[6:0] ? rob_payload_48_rob_idx : _GEN_11962; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11964 = 7'h31 == out_payload_2_rob_idx[6:0] ? rob_payload_49_rob_idx : _GEN_11963; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11965 = 7'h32 == out_payload_2_rob_idx[6:0] ? rob_payload_50_rob_idx : _GEN_11964; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11966 = 7'h33 == out_payload_2_rob_idx[6:0] ? rob_payload_51_rob_idx : _GEN_11965; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11967 = 7'h34 == out_payload_2_rob_idx[6:0] ? rob_payload_52_rob_idx : _GEN_11966; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11968 = 7'h35 == out_payload_2_rob_idx[6:0] ? rob_payload_53_rob_idx : _GEN_11967; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11969 = 7'h36 == out_payload_2_rob_idx[6:0] ? rob_payload_54_rob_idx : _GEN_11968; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11970 = 7'h37 == out_payload_2_rob_idx[6:0] ? rob_payload_55_rob_idx : _GEN_11969; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11971 = 7'h38 == out_payload_2_rob_idx[6:0] ? rob_payload_56_rob_idx : _GEN_11970; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11972 = 7'h39 == out_payload_2_rob_idx[6:0] ? rob_payload_57_rob_idx : _GEN_11971; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11973 = 7'h3a == out_payload_2_rob_idx[6:0] ? rob_payload_58_rob_idx : _GEN_11972; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11974 = 7'h3b == out_payload_2_rob_idx[6:0] ? rob_payload_59_rob_idx : _GEN_11973; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11975 = 7'h3c == out_payload_2_rob_idx[6:0] ? rob_payload_60_rob_idx : _GEN_11974; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11976 = 7'h3d == out_payload_2_rob_idx[6:0] ? rob_payload_61_rob_idx : _GEN_11975; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11977 = 7'h3e == out_payload_2_rob_idx[6:0] ? rob_payload_62_rob_idx : _GEN_11976; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11978 = 7'h3f == out_payload_2_rob_idx[6:0] ? rob_payload_63_rob_idx : _GEN_11977; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11979 = 7'h40 == out_payload_2_rob_idx[6:0] ? rob_payload_64_rob_idx : _GEN_11978; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11980 = 7'h41 == out_payload_2_rob_idx[6:0] ? rob_payload_65_rob_idx : _GEN_11979; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11981 = 7'h42 == out_payload_2_rob_idx[6:0] ? rob_payload_66_rob_idx : _GEN_11980; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11982 = 7'h43 == out_payload_2_rob_idx[6:0] ? rob_payload_67_rob_idx : _GEN_11981; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11983 = 7'h44 == out_payload_2_rob_idx[6:0] ? rob_payload_68_rob_idx : _GEN_11982; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11984 = 7'h45 == out_payload_2_rob_idx[6:0] ? rob_payload_69_rob_idx : _GEN_11983; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11985 = 7'h46 == out_payload_2_rob_idx[6:0] ? rob_payload_70_rob_idx : _GEN_11984; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11986 = 7'h47 == out_payload_2_rob_idx[6:0] ? rob_payload_71_rob_idx : _GEN_11985; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11987 = 7'h48 == out_payload_2_rob_idx[6:0] ? rob_payload_72_rob_idx : _GEN_11986; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11988 = 7'h49 == out_payload_2_rob_idx[6:0] ? rob_payload_73_rob_idx : _GEN_11987; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11989 = 7'h4a == out_payload_2_rob_idx[6:0] ? rob_payload_74_rob_idx : _GEN_11988; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11990 = 7'h4b == out_payload_2_rob_idx[6:0] ? rob_payload_75_rob_idx : _GEN_11989; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11991 = 7'h4c == out_payload_2_rob_idx[6:0] ? rob_payload_76_rob_idx : _GEN_11990; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11992 = 7'h4d == out_payload_2_rob_idx[6:0] ? rob_payload_77_rob_idx : _GEN_11991; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11993 = 7'h4e == out_payload_2_rob_idx[6:0] ? rob_payload_78_rob_idx : _GEN_11992; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11994 = 7'h4f == out_payload_2_rob_idx[6:0] ? rob_payload_79_rob_idx : _GEN_11993; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11995 = 7'h50 == out_payload_2_rob_idx[6:0] ? rob_payload_80_rob_idx : _GEN_11994; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11996 = 7'h51 == out_payload_2_rob_idx[6:0] ? rob_payload_81_rob_idx : _GEN_11995; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11997 = 7'h52 == out_payload_2_rob_idx[6:0] ? rob_payload_82_rob_idx : _GEN_11996; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11998 = 7'h53 == out_payload_2_rob_idx[6:0] ? rob_payload_83_rob_idx : _GEN_11997; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_11999 = 7'h54 == out_payload_2_rob_idx[6:0] ? rob_payload_84_rob_idx : _GEN_11998; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12000 = 7'h55 == out_payload_2_rob_idx[6:0] ? rob_payload_85_rob_idx : _GEN_11999; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12001 = 7'h56 == out_payload_2_rob_idx[6:0] ? rob_payload_86_rob_idx : _GEN_12000; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12002 = 7'h57 == out_payload_2_rob_idx[6:0] ? rob_payload_87_rob_idx : _GEN_12001; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12003 = 7'h58 == out_payload_2_rob_idx[6:0] ? rob_payload_88_rob_idx : _GEN_12002; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12004 = 7'h59 == out_payload_2_rob_idx[6:0] ? rob_payload_89_rob_idx : _GEN_12003; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12005 = 7'h5a == out_payload_2_rob_idx[6:0] ? rob_payload_90_rob_idx : _GEN_12004; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12006 = 7'h5b == out_payload_2_rob_idx[6:0] ? rob_payload_91_rob_idx : _GEN_12005; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12007 = 7'h5c == out_payload_2_rob_idx[6:0] ? rob_payload_92_rob_idx : _GEN_12006; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12008 = 7'h5d == out_payload_2_rob_idx[6:0] ? rob_payload_93_rob_idx : _GEN_12007; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12009 = 7'h5e == out_payload_2_rob_idx[6:0] ? rob_payload_94_rob_idx : _GEN_12008; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12010 = 7'h5f == out_payload_2_rob_idx[6:0] ? rob_payload_95_rob_idx : _GEN_12009; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12011 = 7'h60 == out_payload_2_rob_idx[6:0] ? rob_payload_96_rob_idx : _GEN_12010; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12012 = 7'h61 == out_payload_2_rob_idx[6:0] ? rob_payload_97_rob_idx : _GEN_12011; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12013 = 7'h62 == out_payload_2_rob_idx[6:0] ? rob_payload_98_rob_idx : _GEN_12012; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12014 = 7'h63 == out_payload_2_rob_idx[6:0] ? rob_payload_99_rob_idx : _GEN_12013; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12015 = 7'h64 == out_payload_2_rob_idx[6:0] ? rob_payload_100_rob_idx : _GEN_12014; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12016 = 7'h65 == out_payload_2_rob_idx[6:0] ? rob_payload_101_rob_idx : _GEN_12015; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12017 = 7'h66 == out_payload_2_rob_idx[6:0] ? rob_payload_102_rob_idx : _GEN_12016; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12018 = 7'h67 == out_payload_2_rob_idx[6:0] ? rob_payload_103_rob_idx : _GEN_12017; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12019 = 7'h68 == out_payload_2_rob_idx[6:0] ? rob_payload_104_rob_idx : _GEN_12018; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12020 = 7'h69 == out_payload_2_rob_idx[6:0] ? rob_payload_105_rob_idx : _GEN_12019; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12021 = 7'h6a == out_payload_2_rob_idx[6:0] ? rob_payload_106_rob_idx : _GEN_12020; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12022 = 7'h6b == out_payload_2_rob_idx[6:0] ? rob_payload_107_rob_idx : _GEN_12021; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12023 = 7'h6c == out_payload_2_rob_idx[6:0] ? rob_payload_108_rob_idx : _GEN_12022; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12024 = 7'h6d == out_payload_2_rob_idx[6:0] ? rob_payload_109_rob_idx : _GEN_12023; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12025 = 7'h6e == out_payload_2_rob_idx[6:0] ? rob_payload_110_rob_idx : _GEN_12024; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12026 = 7'h6f == out_payload_2_rob_idx[6:0] ? rob_payload_111_rob_idx : _GEN_12025; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12027 = 7'h70 == out_payload_2_rob_idx[6:0] ? rob_payload_112_rob_idx : _GEN_12026; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12028 = 7'h71 == out_payload_2_rob_idx[6:0] ? rob_payload_113_rob_idx : _GEN_12027; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12029 = 7'h72 == out_payload_2_rob_idx[6:0] ? rob_payload_114_rob_idx : _GEN_12028; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12030 = 7'h73 == out_payload_2_rob_idx[6:0] ? rob_payload_115_rob_idx : _GEN_12029; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12031 = 7'h74 == out_payload_2_rob_idx[6:0] ? rob_payload_116_rob_idx : _GEN_12030; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12032 = 7'h75 == out_payload_2_rob_idx[6:0] ? rob_payload_117_rob_idx : _GEN_12031; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12033 = 7'h76 == out_payload_2_rob_idx[6:0] ? rob_payload_118_rob_idx : _GEN_12032; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12034 = 7'h77 == out_payload_2_rob_idx[6:0] ? rob_payload_119_rob_idx : _GEN_12033; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12035 = 7'h78 == out_payload_2_rob_idx[6:0] ? rob_payload_120_rob_idx : _GEN_12034; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12036 = 7'h79 == out_payload_2_rob_idx[6:0] ? rob_payload_121_rob_idx : _GEN_12035; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12037 = 7'h7a == out_payload_2_rob_idx[6:0] ? rob_payload_122_rob_idx : _GEN_12036; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12038 = 7'h7b == out_payload_2_rob_idx[6:0] ? rob_payload_123_rob_idx : _GEN_12037; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12039 = 7'h7c == out_payload_2_rob_idx[6:0] ? rob_payload_124_rob_idx : _GEN_12038; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12040 = 7'h7d == out_payload_2_rob_idx[6:0] ? rob_payload_125_rob_idx : _GEN_12039; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12041 = 7'h7e == out_payload_2_rob_idx[6:0] ? rob_payload_126_rob_idx : _GEN_12040; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12042 = 7'h7f == out_payload_2_rob_idx[6:0] ? rob_payload_127_rob_idx : _GEN_12041; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12044 = 7'h1 == out_payload_2_rob_idx[6:0] ? rob_payload_1_flits_fired : rob_payload_0_flits_fired; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12045 = 7'h2 == out_payload_2_rob_idx[6:0] ? rob_payload_2_flits_fired : _GEN_12044; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12046 = 7'h3 == out_payload_2_rob_idx[6:0] ? rob_payload_3_flits_fired : _GEN_12045; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12047 = 7'h4 == out_payload_2_rob_idx[6:0] ? rob_payload_4_flits_fired : _GEN_12046; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12048 = 7'h5 == out_payload_2_rob_idx[6:0] ? rob_payload_5_flits_fired : _GEN_12047; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12049 = 7'h6 == out_payload_2_rob_idx[6:0] ? rob_payload_6_flits_fired : _GEN_12048; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12050 = 7'h7 == out_payload_2_rob_idx[6:0] ? rob_payload_7_flits_fired : _GEN_12049; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12051 = 7'h8 == out_payload_2_rob_idx[6:0] ? rob_payload_8_flits_fired : _GEN_12050; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12052 = 7'h9 == out_payload_2_rob_idx[6:0] ? rob_payload_9_flits_fired : _GEN_12051; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12053 = 7'ha == out_payload_2_rob_idx[6:0] ? rob_payload_10_flits_fired : _GEN_12052; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12054 = 7'hb == out_payload_2_rob_idx[6:0] ? rob_payload_11_flits_fired : _GEN_12053; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12055 = 7'hc == out_payload_2_rob_idx[6:0] ? rob_payload_12_flits_fired : _GEN_12054; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12056 = 7'hd == out_payload_2_rob_idx[6:0] ? rob_payload_13_flits_fired : _GEN_12055; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12057 = 7'he == out_payload_2_rob_idx[6:0] ? rob_payload_14_flits_fired : _GEN_12056; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12058 = 7'hf == out_payload_2_rob_idx[6:0] ? rob_payload_15_flits_fired : _GEN_12057; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12059 = 7'h10 == out_payload_2_rob_idx[6:0] ? rob_payload_16_flits_fired : _GEN_12058; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12060 = 7'h11 == out_payload_2_rob_idx[6:0] ? rob_payload_17_flits_fired : _GEN_12059; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12061 = 7'h12 == out_payload_2_rob_idx[6:0] ? rob_payload_18_flits_fired : _GEN_12060; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12062 = 7'h13 == out_payload_2_rob_idx[6:0] ? rob_payload_19_flits_fired : _GEN_12061; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12063 = 7'h14 == out_payload_2_rob_idx[6:0] ? rob_payload_20_flits_fired : _GEN_12062; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12064 = 7'h15 == out_payload_2_rob_idx[6:0] ? rob_payload_21_flits_fired : _GEN_12063; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12065 = 7'h16 == out_payload_2_rob_idx[6:0] ? rob_payload_22_flits_fired : _GEN_12064; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12066 = 7'h17 == out_payload_2_rob_idx[6:0] ? rob_payload_23_flits_fired : _GEN_12065; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12067 = 7'h18 == out_payload_2_rob_idx[6:0] ? rob_payload_24_flits_fired : _GEN_12066; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12068 = 7'h19 == out_payload_2_rob_idx[6:0] ? rob_payload_25_flits_fired : _GEN_12067; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12069 = 7'h1a == out_payload_2_rob_idx[6:0] ? rob_payload_26_flits_fired : _GEN_12068; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12070 = 7'h1b == out_payload_2_rob_idx[6:0] ? rob_payload_27_flits_fired : _GEN_12069; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12071 = 7'h1c == out_payload_2_rob_idx[6:0] ? rob_payload_28_flits_fired : _GEN_12070; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12072 = 7'h1d == out_payload_2_rob_idx[6:0] ? rob_payload_29_flits_fired : _GEN_12071; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12073 = 7'h1e == out_payload_2_rob_idx[6:0] ? rob_payload_30_flits_fired : _GEN_12072; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12074 = 7'h1f == out_payload_2_rob_idx[6:0] ? rob_payload_31_flits_fired : _GEN_12073; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12075 = 7'h20 == out_payload_2_rob_idx[6:0] ? rob_payload_32_flits_fired : _GEN_12074; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12076 = 7'h21 == out_payload_2_rob_idx[6:0] ? rob_payload_33_flits_fired : _GEN_12075; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12077 = 7'h22 == out_payload_2_rob_idx[6:0] ? rob_payload_34_flits_fired : _GEN_12076; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12078 = 7'h23 == out_payload_2_rob_idx[6:0] ? rob_payload_35_flits_fired : _GEN_12077; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12079 = 7'h24 == out_payload_2_rob_idx[6:0] ? rob_payload_36_flits_fired : _GEN_12078; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12080 = 7'h25 == out_payload_2_rob_idx[6:0] ? rob_payload_37_flits_fired : _GEN_12079; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12081 = 7'h26 == out_payload_2_rob_idx[6:0] ? rob_payload_38_flits_fired : _GEN_12080; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12082 = 7'h27 == out_payload_2_rob_idx[6:0] ? rob_payload_39_flits_fired : _GEN_12081; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12083 = 7'h28 == out_payload_2_rob_idx[6:0] ? rob_payload_40_flits_fired : _GEN_12082; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12084 = 7'h29 == out_payload_2_rob_idx[6:0] ? rob_payload_41_flits_fired : _GEN_12083; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12085 = 7'h2a == out_payload_2_rob_idx[6:0] ? rob_payload_42_flits_fired : _GEN_12084; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12086 = 7'h2b == out_payload_2_rob_idx[6:0] ? rob_payload_43_flits_fired : _GEN_12085; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12087 = 7'h2c == out_payload_2_rob_idx[6:0] ? rob_payload_44_flits_fired : _GEN_12086; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12088 = 7'h2d == out_payload_2_rob_idx[6:0] ? rob_payload_45_flits_fired : _GEN_12087; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12089 = 7'h2e == out_payload_2_rob_idx[6:0] ? rob_payload_46_flits_fired : _GEN_12088; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12090 = 7'h2f == out_payload_2_rob_idx[6:0] ? rob_payload_47_flits_fired : _GEN_12089; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12091 = 7'h30 == out_payload_2_rob_idx[6:0] ? rob_payload_48_flits_fired : _GEN_12090; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12092 = 7'h31 == out_payload_2_rob_idx[6:0] ? rob_payload_49_flits_fired : _GEN_12091; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12093 = 7'h32 == out_payload_2_rob_idx[6:0] ? rob_payload_50_flits_fired : _GEN_12092; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12094 = 7'h33 == out_payload_2_rob_idx[6:0] ? rob_payload_51_flits_fired : _GEN_12093; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12095 = 7'h34 == out_payload_2_rob_idx[6:0] ? rob_payload_52_flits_fired : _GEN_12094; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12096 = 7'h35 == out_payload_2_rob_idx[6:0] ? rob_payload_53_flits_fired : _GEN_12095; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12097 = 7'h36 == out_payload_2_rob_idx[6:0] ? rob_payload_54_flits_fired : _GEN_12096; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12098 = 7'h37 == out_payload_2_rob_idx[6:0] ? rob_payload_55_flits_fired : _GEN_12097; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12099 = 7'h38 == out_payload_2_rob_idx[6:0] ? rob_payload_56_flits_fired : _GEN_12098; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12100 = 7'h39 == out_payload_2_rob_idx[6:0] ? rob_payload_57_flits_fired : _GEN_12099; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12101 = 7'h3a == out_payload_2_rob_idx[6:0] ? rob_payload_58_flits_fired : _GEN_12100; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12102 = 7'h3b == out_payload_2_rob_idx[6:0] ? rob_payload_59_flits_fired : _GEN_12101; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12103 = 7'h3c == out_payload_2_rob_idx[6:0] ? rob_payload_60_flits_fired : _GEN_12102; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12104 = 7'h3d == out_payload_2_rob_idx[6:0] ? rob_payload_61_flits_fired : _GEN_12103; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12105 = 7'h3e == out_payload_2_rob_idx[6:0] ? rob_payload_62_flits_fired : _GEN_12104; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12106 = 7'h3f == out_payload_2_rob_idx[6:0] ? rob_payload_63_flits_fired : _GEN_12105; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12107 = 7'h40 == out_payload_2_rob_idx[6:0] ? rob_payload_64_flits_fired : _GEN_12106; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12108 = 7'h41 == out_payload_2_rob_idx[6:0] ? rob_payload_65_flits_fired : _GEN_12107; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12109 = 7'h42 == out_payload_2_rob_idx[6:0] ? rob_payload_66_flits_fired : _GEN_12108; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12110 = 7'h43 == out_payload_2_rob_idx[6:0] ? rob_payload_67_flits_fired : _GEN_12109; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12111 = 7'h44 == out_payload_2_rob_idx[6:0] ? rob_payload_68_flits_fired : _GEN_12110; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12112 = 7'h45 == out_payload_2_rob_idx[6:0] ? rob_payload_69_flits_fired : _GEN_12111; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12113 = 7'h46 == out_payload_2_rob_idx[6:0] ? rob_payload_70_flits_fired : _GEN_12112; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12114 = 7'h47 == out_payload_2_rob_idx[6:0] ? rob_payload_71_flits_fired : _GEN_12113; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12115 = 7'h48 == out_payload_2_rob_idx[6:0] ? rob_payload_72_flits_fired : _GEN_12114; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12116 = 7'h49 == out_payload_2_rob_idx[6:0] ? rob_payload_73_flits_fired : _GEN_12115; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12117 = 7'h4a == out_payload_2_rob_idx[6:0] ? rob_payload_74_flits_fired : _GEN_12116; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12118 = 7'h4b == out_payload_2_rob_idx[6:0] ? rob_payload_75_flits_fired : _GEN_12117; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12119 = 7'h4c == out_payload_2_rob_idx[6:0] ? rob_payload_76_flits_fired : _GEN_12118; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12120 = 7'h4d == out_payload_2_rob_idx[6:0] ? rob_payload_77_flits_fired : _GEN_12119; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12121 = 7'h4e == out_payload_2_rob_idx[6:0] ? rob_payload_78_flits_fired : _GEN_12120; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12122 = 7'h4f == out_payload_2_rob_idx[6:0] ? rob_payload_79_flits_fired : _GEN_12121; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12123 = 7'h50 == out_payload_2_rob_idx[6:0] ? rob_payload_80_flits_fired : _GEN_12122; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12124 = 7'h51 == out_payload_2_rob_idx[6:0] ? rob_payload_81_flits_fired : _GEN_12123; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12125 = 7'h52 == out_payload_2_rob_idx[6:0] ? rob_payload_82_flits_fired : _GEN_12124; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12126 = 7'h53 == out_payload_2_rob_idx[6:0] ? rob_payload_83_flits_fired : _GEN_12125; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12127 = 7'h54 == out_payload_2_rob_idx[6:0] ? rob_payload_84_flits_fired : _GEN_12126; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12128 = 7'h55 == out_payload_2_rob_idx[6:0] ? rob_payload_85_flits_fired : _GEN_12127; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12129 = 7'h56 == out_payload_2_rob_idx[6:0] ? rob_payload_86_flits_fired : _GEN_12128; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12130 = 7'h57 == out_payload_2_rob_idx[6:0] ? rob_payload_87_flits_fired : _GEN_12129; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12131 = 7'h58 == out_payload_2_rob_idx[6:0] ? rob_payload_88_flits_fired : _GEN_12130; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12132 = 7'h59 == out_payload_2_rob_idx[6:0] ? rob_payload_89_flits_fired : _GEN_12131; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12133 = 7'h5a == out_payload_2_rob_idx[6:0] ? rob_payload_90_flits_fired : _GEN_12132; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12134 = 7'h5b == out_payload_2_rob_idx[6:0] ? rob_payload_91_flits_fired : _GEN_12133; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12135 = 7'h5c == out_payload_2_rob_idx[6:0] ? rob_payload_92_flits_fired : _GEN_12134; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12136 = 7'h5d == out_payload_2_rob_idx[6:0] ? rob_payload_93_flits_fired : _GEN_12135; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12137 = 7'h5e == out_payload_2_rob_idx[6:0] ? rob_payload_94_flits_fired : _GEN_12136; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12138 = 7'h5f == out_payload_2_rob_idx[6:0] ? rob_payload_95_flits_fired : _GEN_12137; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12139 = 7'h60 == out_payload_2_rob_idx[6:0] ? rob_payload_96_flits_fired : _GEN_12138; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12140 = 7'h61 == out_payload_2_rob_idx[6:0] ? rob_payload_97_flits_fired : _GEN_12139; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12141 = 7'h62 == out_payload_2_rob_idx[6:0] ? rob_payload_98_flits_fired : _GEN_12140; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12142 = 7'h63 == out_payload_2_rob_idx[6:0] ? rob_payload_99_flits_fired : _GEN_12141; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12143 = 7'h64 == out_payload_2_rob_idx[6:0] ? rob_payload_100_flits_fired : _GEN_12142; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12144 = 7'h65 == out_payload_2_rob_idx[6:0] ? rob_payload_101_flits_fired : _GEN_12143; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12145 = 7'h66 == out_payload_2_rob_idx[6:0] ? rob_payload_102_flits_fired : _GEN_12144; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12146 = 7'h67 == out_payload_2_rob_idx[6:0] ? rob_payload_103_flits_fired : _GEN_12145; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12147 = 7'h68 == out_payload_2_rob_idx[6:0] ? rob_payload_104_flits_fired : _GEN_12146; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12148 = 7'h69 == out_payload_2_rob_idx[6:0] ? rob_payload_105_flits_fired : _GEN_12147; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12149 = 7'h6a == out_payload_2_rob_idx[6:0] ? rob_payload_106_flits_fired : _GEN_12148; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12150 = 7'h6b == out_payload_2_rob_idx[6:0] ? rob_payload_107_flits_fired : _GEN_12149; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12151 = 7'h6c == out_payload_2_rob_idx[6:0] ? rob_payload_108_flits_fired : _GEN_12150; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12152 = 7'h6d == out_payload_2_rob_idx[6:0] ? rob_payload_109_flits_fired : _GEN_12151; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12153 = 7'h6e == out_payload_2_rob_idx[6:0] ? rob_payload_110_flits_fired : _GEN_12152; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12154 = 7'h6f == out_payload_2_rob_idx[6:0] ? rob_payload_111_flits_fired : _GEN_12153; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12155 = 7'h70 == out_payload_2_rob_idx[6:0] ? rob_payload_112_flits_fired : _GEN_12154; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12156 = 7'h71 == out_payload_2_rob_idx[6:0] ? rob_payload_113_flits_fired : _GEN_12155; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12157 = 7'h72 == out_payload_2_rob_idx[6:0] ? rob_payload_114_flits_fired : _GEN_12156; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12158 = 7'h73 == out_payload_2_rob_idx[6:0] ? rob_payload_115_flits_fired : _GEN_12157; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12159 = 7'h74 == out_payload_2_rob_idx[6:0] ? rob_payload_116_flits_fired : _GEN_12158; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12160 = 7'h75 == out_payload_2_rob_idx[6:0] ? rob_payload_117_flits_fired : _GEN_12159; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12161 = 7'h76 == out_payload_2_rob_idx[6:0] ? rob_payload_118_flits_fired : _GEN_12160; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12162 = 7'h77 == out_payload_2_rob_idx[6:0] ? rob_payload_119_flits_fired : _GEN_12161; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12163 = 7'h78 == out_payload_2_rob_idx[6:0] ? rob_payload_120_flits_fired : _GEN_12162; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12164 = 7'h79 == out_payload_2_rob_idx[6:0] ? rob_payload_121_flits_fired : _GEN_12163; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12165 = 7'h7a == out_payload_2_rob_idx[6:0] ? rob_payload_122_flits_fired : _GEN_12164; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12166 = 7'h7b == out_payload_2_rob_idx[6:0] ? rob_payload_123_flits_fired : _GEN_12165; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12167 = 7'h7c == out_payload_2_rob_idx[6:0] ? rob_payload_124_flits_fired : _GEN_12166; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12168 = 7'h7d == out_payload_2_rob_idx[6:0] ? rob_payload_125_flits_fired : _GEN_12167; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12169 = 7'h7e == out_payload_2_rob_idx[6:0] ? rob_payload_126_flits_fired : _GEN_12168; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_12170 = 7'h7f == out_payload_2_rob_idx[6:0] ? rob_payload_127_flits_fired : _GEN_12169; // @[TestHarness.scala 202:{35,35}]
  wire [63:0] _T_176 = {_GEN_11914,_GEN_12042,_GEN_12170}; // @[TestHarness.scala 202:35]
  wire [1:0] _GEN_12172 = 7'h1 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_1 : rob_ingress_id_0; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12173 = 7'h2 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_2 : _GEN_12172; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12174 = 7'h3 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_3 : _GEN_12173; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12175 = 7'h4 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_4 : _GEN_12174; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12176 = 7'h5 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_5 : _GEN_12175; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12177 = 7'h6 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_6 : _GEN_12176; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12178 = 7'h7 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_7 : _GEN_12177; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12179 = 7'h8 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_8 : _GEN_12178; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12180 = 7'h9 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_9 : _GEN_12179; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12181 = 7'ha == out_payload_2_rob_idx[6:0] ? rob_ingress_id_10 : _GEN_12180; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12182 = 7'hb == out_payload_2_rob_idx[6:0] ? rob_ingress_id_11 : _GEN_12181; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12183 = 7'hc == out_payload_2_rob_idx[6:0] ? rob_ingress_id_12 : _GEN_12182; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12184 = 7'hd == out_payload_2_rob_idx[6:0] ? rob_ingress_id_13 : _GEN_12183; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12185 = 7'he == out_payload_2_rob_idx[6:0] ? rob_ingress_id_14 : _GEN_12184; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12186 = 7'hf == out_payload_2_rob_idx[6:0] ? rob_ingress_id_15 : _GEN_12185; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12187 = 7'h10 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_16 : _GEN_12186; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12188 = 7'h11 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_17 : _GEN_12187; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12189 = 7'h12 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_18 : _GEN_12188; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12190 = 7'h13 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_19 : _GEN_12189; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12191 = 7'h14 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_20 : _GEN_12190; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12192 = 7'h15 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_21 : _GEN_12191; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12193 = 7'h16 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_22 : _GEN_12192; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12194 = 7'h17 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_23 : _GEN_12193; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12195 = 7'h18 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_24 : _GEN_12194; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12196 = 7'h19 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_25 : _GEN_12195; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12197 = 7'h1a == out_payload_2_rob_idx[6:0] ? rob_ingress_id_26 : _GEN_12196; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12198 = 7'h1b == out_payload_2_rob_idx[6:0] ? rob_ingress_id_27 : _GEN_12197; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12199 = 7'h1c == out_payload_2_rob_idx[6:0] ? rob_ingress_id_28 : _GEN_12198; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12200 = 7'h1d == out_payload_2_rob_idx[6:0] ? rob_ingress_id_29 : _GEN_12199; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12201 = 7'h1e == out_payload_2_rob_idx[6:0] ? rob_ingress_id_30 : _GEN_12200; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12202 = 7'h1f == out_payload_2_rob_idx[6:0] ? rob_ingress_id_31 : _GEN_12201; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12203 = 7'h20 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_32 : _GEN_12202; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12204 = 7'h21 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_33 : _GEN_12203; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12205 = 7'h22 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_34 : _GEN_12204; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12206 = 7'h23 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_35 : _GEN_12205; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12207 = 7'h24 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_36 : _GEN_12206; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12208 = 7'h25 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_37 : _GEN_12207; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12209 = 7'h26 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_38 : _GEN_12208; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12210 = 7'h27 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_39 : _GEN_12209; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12211 = 7'h28 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_40 : _GEN_12210; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12212 = 7'h29 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_41 : _GEN_12211; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12213 = 7'h2a == out_payload_2_rob_idx[6:0] ? rob_ingress_id_42 : _GEN_12212; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12214 = 7'h2b == out_payload_2_rob_idx[6:0] ? rob_ingress_id_43 : _GEN_12213; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12215 = 7'h2c == out_payload_2_rob_idx[6:0] ? rob_ingress_id_44 : _GEN_12214; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12216 = 7'h2d == out_payload_2_rob_idx[6:0] ? rob_ingress_id_45 : _GEN_12215; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12217 = 7'h2e == out_payload_2_rob_idx[6:0] ? rob_ingress_id_46 : _GEN_12216; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12218 = 7'h2f == out_payload_2_rob_idx[6:0] ? rob_ingress_id_47 : _GEN_12217; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12219 = 7'h30 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_48 : _GEN_12218; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12220 = 7'h31 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_49 : _GEN_12219; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12221 = 7'h32 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_50 : _GEN_12220; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12222 = 7'h33 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_51 : _GEN_12221; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12223 = 7'h34 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_52 : _GEN_12222; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12224 = 7'h35 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_53 : _GEN_12223; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12225 = 7'h36 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_54 : _GEN_12224; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12226 = 7'h37 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_55 : _GEN_12225; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12227 = 7'h38 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_56 : _GEN_12226; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12228 = 7'h39 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_57 : _GEN_12227; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12229 = 7'h3a == out_payload_2_rob_idx[6:0] ? rob_ingress_id_58 : _GEN_12228; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12230 = 7'h3b == out_payload_2_rob_idx[6:0] ? rob_ingress_id_59 : _GEN_12229; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12231 = 7'h3c == out_payload_2_rob_idx[6:0] ? rob_ingress_id_60 : _GEN_12230; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12232 = 7'h3d == out_payload_2_rob_idx[6:0] ? rob_ingress_id_61 : _GEN_12231; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12233 = 7'h3e == out_payload_2_rob_idx[6:0] ? rob_ingress_id_62 : _GEN_12232; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12234 = 7'h3f == out_payload_2_rob_idx[6:0] ? rob_ingress_id_63 : _GEN_12233; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12235 = 7'h40 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_64 : _GEN_12234; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12236 = 7'h41 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_65 : _GEN_12235; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12237 = 7'h42 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_66 : _GEN_12236; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12238 = 7'h43 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_67 : _GEN_12237; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12239 = 7'h44 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_68 : _GEN_12238; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12240 = 7'h45 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_69 : _GEN_12239; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12241 = 7'h46 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_70 : _GEN_12240; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12242 = 7'h47 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_71 : _GEN_12241; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12243 = 7'h48 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_72 : _GEN_12242; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12244 = 7'h49 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_73 : _GEN_12243; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12245 = 7'h4a == out_payload_2_rob_idx[6:0] ? rob_ingress_id_74 : _GEN_12244; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12246 = 7'h4b == out_payload_2_rob_idx[6:0] ? rob_ingress_id_75 : _GEN_12245; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12247 = 7'h4c == out_payload_2_rob_idx[6:0] ? rob_ingress_id_76 : _GEN_12246; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12248 = 7'h4d == out_payload_2_rob_idx[6:0] ? rob_ingress_id_77 : _GEN_12247; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12249 = 7'h4e == out_payload_2_rob_idx[6:0] ? rob_ingress_id_78 : _GEN_12248; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12250 = 7'h4f == out_payload_2_rob_idx[6:0] ? rob_ingress_id_79 : _GEN_12249; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12251 = 7'h50 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_80 : _GEN_12250; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12252 = 7'h51 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_81 : _GEN_12251; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12253 = 7'h52 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_82 : _GEN_12252; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12254 = 7'h53 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_83 : _GEN_12253; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12255 = 7'h54 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_84 : _GEN_12254; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12256 = 7'h55 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_85 : _GEN_12255; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12257 = 7'h56 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_86 : _GEN_12256; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12258 = 7'h57 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_87 : _GEN_12257; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12259 = 7'h58 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_88 : _GEN_12258; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12260 = 7'h59 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_89 : _GEN_12259; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12261 = 7'h5a == out_payload_2_rob_idx[6:0] ? rob_ingress_id_90 : _GEN_12260; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12262 = 7'h5b == out_payload_2_rob_idx[6:0] ? rob_ingress_id_91 : _GEN_12261; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12263 = 7'h5c == out_payload_2_rob_idx[6:0] ? rob_ingress_id_92 : _GEN_12262; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12264 = 7'h5d == out_payload_2_rob_idx[6:0] ? rob_ingress_id_93 : _GEN_12263; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12265 = 7'h5e == out_payload_2_rob_idx[6:0] ? rob_ingress_id_94 : _GEN_12264; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12266 = 7'h5f == out_payload_2_rob_idx[6:0] ? rob_ingress_id_95 : _GEN_12265; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12267 = 7'h60 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_96 : _GEN_12266; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12268 = 7'h61 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_97 : _GEN_12267; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12269 = 7'h62 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_98 : _GEN_12268; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12270 = 7'h63 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_99 : _GEN_12269; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12271 = 7'h64 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_100 : _GEN_12270; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12272 = 7'h65 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_101 : _GEN_12271; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12273 = 7'h66 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_102 : _GEN_12272; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12274 = 7'h67 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_103 : _GEN_12273; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12275 = 7'h68 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_104 : _GEN_12274; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12276 = 7'h69 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_105 : _GEN_12275; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12277 = 7'h6a == out_payload_2_rob_idx[6:0] ? rob_ingress_id_106 : _GEN_12276; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12278 = 7'h6b == out_payload_2_rob_idx[6:0] ? rob_ingress_id_107 : _GEN_12277; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12279 = 7'h6c == out_payload_2_rob_idx[6:0] ? rob_ingress_id_108 : _GEN_12278; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12280 = 7'h6d == out_payload_2_rob_idx[6:0] ? rob_ingress_id_109 : _GEN_12279; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12281 = 7'h6e == out_payload_2_rob_idx[6:0] ? rob_ingress_id_110 : _GEN_12280; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12282 = 7'h6f == out_payload_2_rob_idx[6:0] ? rob_ingress_id_111 : _GEN_12281; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12283 = 7'h70 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_112 : _GEN_12282; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12284 = 7'h71 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_113 : _GEN_12283; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12285 = 7'h72 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_114 : _GEN_12284; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12286 = 7'h73 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_115 : _GEN_12285; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12287 = 7'h74 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_116 : _GEN_12286; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12288 = 7'h75 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_117 : _GEN_12287; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12289 = 7'h76 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_118 : _GEN_12288; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12290 = 7'h77 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_119 : _GEN_12289; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12291 = 7'h78 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_120 : _GEN_12290; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12292 = 7'h79 == out_payload_2_rob_idx[6:0] ? rob_ingress_id_121 : _GEN_12291; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12293 = 7'h7a == out_payload_2_rob_idx[6:0] ? rob_ingress_id_122 : _GEN_12292; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12294 = 7'h7b == out_payload_2_rob_idx[6:0] ? rob_ingress_id_123 : _GEN_12293; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12295 = 7'h7c == out_payload_2_rob_idx[6:0] ? rob_ingress_id_124 : _GEN_12294; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12296 = 7'h7d == out_payload_2_rob_idx[6:0] ? rob_ingress_id_125 : _GEN_12295; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12297 = 7'h7e == out_payload_2_rob_idx[6:0] ? rob_ingress_id_126 : _GEN_12296; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12298 = 7'h7f == out_payload_2_rob_idx[6:0] ? rob_ingress_id_127 : _GEN_12297; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_12300 = 7'h1 == out_payload_2_rob_idx[6:0] ? rob_egress_id_1 : rob_egress_id_0; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12301 = 7'h2 == out_payload_2_rob_idx[6:0] ? rob_egress_id_2 : _GEN_12300; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12302 = 7'h3 == out_payload_2_rob_idx[6:0] ? rob_egress_id_3 : _GEN_12301; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12303 = 7'h4 == out_payload_2_rob_idx[6:0] ? rob_egress_id_4 : _GEN_12302; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12304 = 7'h5 == out_payload_2_rob_idx[6:0] ? rob_egress_id_5 : _GEN_12303; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12305 = 7'h6 == out_payload_2_rob_idx[6:0] ? rob_egress_id_6 : _GEN_12304; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12306 = 7'h7 == out_payload_2_rob_idx[6:0] ? rob_egress_id_7 : _GEN_12305; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12307 = 7'h8 == out_payload_2_rob_idx[6:0] ? rob_egress_id_8 : _GEN_12306; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12308 = 7'h9 == out_payload_2_rob_idx[6:0] ? rob_egress_id_9 : _GEN_12307; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12309 = 7'ha == out_payload_2_rob_idx[6:0] ? rob_egress_id_10 : _GEN_12308; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12310 = 7'hb == out_payload_2_rob_idx[6:0] ? rob_egress_id_11 : _GEN_12309; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12311 = 7'hc == out_payload_2_rob_idx[6:0] ? rob_egress_id_12 : _GEN_12310; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12312 = 7'hd == out_payload_2_rob_idx[6:0] ? rob_egress_id_13 : _GEN_12311; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12313 = 7'he == out_payload_2_rob_idx[6:0] ? rob_egress_id_14 : _GEN_12312; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12314 = 7'hf == out_payload_2_rob_idx[6:0] ? rob_egress_id_15 : _GEN_12313; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12315 = 7'h10 == out_payload_2_rob_idx[6:0] ? rob_egress_id_16 : _GEN_12314; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12316 = 7'h11 == out_payload_2_rob_idx[6:0] ? rob_egress_id_17 : _GEN_12315; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12317 = 7'h12 == out_payload_2_rob_idx[6:0] ? rob_egress_id_18 : _GEN_12316; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12318 = 7'h13 == out_payload_2_rob_idx[6:0] ? rob_egress_id_19 : _GEN_12317; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12319 = 7'h14 == out_payload_2_rob_idx[6:0] ? rob_egress_id_20 : _GEN_12318; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12320 = 7'h15 == out_payload_2_rob_idx[6:0] ? rob_egress_id_21 : _GEN_12319; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12321 = 7'h16 == out_payload_2_rob_idx[6:0] ? rob_egress_id_22 : _GEN_12320; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12322 = 7'h17 == out_payload_2_rob_idx[6:0] ? rob_egress_id_23 : _GEN_12321; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12323 = 7'h18 == out_payload_2_rob_idx[6:0] ? rob_egress_id_24 : _GEN_12322; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12324 = 7'h19 == out_payload_2_rob_idx[6:0] ? rob_egress_id_25 : _GEN_12323; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12325 = 7'h1a == out_payload_2_rob_idx[6:0] ? rob_egress_id_26 : _GEN_12324; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12326 = 7'h1b == out_payload_2_rob_idx[6:0] ? rob_egress_id_27 : _GEN_12325; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12327 = 7'h1c == out_payload_2_rob_idx[6:0] ? rob_egress_id_28 : _GEN_12326; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12328 = 7'h1d == out_payload_2_rob_idx[6:0] ? rob_egress_id_29 : _GEN_12327; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12329 = 7'h1e == out_payload_2_rob_idx[6:0] ? rob_egress_id_30 : _GEN_12328; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12330 = 7'h1f == out_payload_2_rob_idx[6:0] ? rob_egress_id_31 : _GEN_12329; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12331 = 7'h20 == out_payload_2_rob_idx[6:0] ? rob_egress_id_32 : _GEN_12330; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12332 = 7'h21 == out_payload_2_rob_idx[6:0] ? rob_egress_id_33 : _GEN_12331; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12333 = 7'h22 == out_payload_2_rob_idx[6:0] ? rob_egress_id_34 : _GEN_12332; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12334 = 7'h23 == out_payload_2_rob_idx[6:0] ? rob_egress_id_35 : _GEN_12333; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12335 = 7'h24 == out_payload_2_rob_idx[6:0] ? rob_egress_id_36 : _GEN_12334; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12336 = 7'h25 == out_payload_2_rob_idx[6:0] ? rob_egress_id_37 : _GEN_12335; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12337 = 7'h26 == out_payload_2_rob_idx[6:0] ? rob_egress_id_38 : _GEN_12336; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12338 = 7'h27 == out_payload_2_rob_idx[6:0] ? rob_egress_id_39 : _GEN_12337; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12339 = 7'h28 == out_payload_2_rob_idx[6:0] ? rob_egress_id_40 : _GEN_12338; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12340 = 7'h29 == out_payload_2_rob_idx[6:0] ? rob_egress_id_41 : _GEN_12339; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12341 = 7'h2a == out_payload_2_rob_idx[6:0] ? rob_egress_id_42 : _GEN_12340; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12342 = 7'h2b == out_payload_2_rob_idx[6:0] ? rob_egress_id_43 : _GEN_12341; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12343 = 7'h2c == out_payload_2_rob_idx[6:0] ? rob_egress_id_44 : _GEN_12342; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12344 = 7'h2d == out_payload_2_rob_idx[6:0] ? rob_egress_id_45 : _GEN_12343; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12345 = 7'h2e == out_payload_2_rob_idx[6:0] ? rob_egress_id_46 : _GEN_12344; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12346 = 7'h2f == out_payload_2_rob_idx[6:0] ? rob_egress_id_47 : _GEN_12345; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12347 = 7'h30 == out_payload_2_rob_idx[6:0] ? rob_egress_id_48 : _GEN_12346; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12348 = 7'h31 == out_payload_2_rob_idx[6:0] ? rob_egress_id_49 : _GEN_12347; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12349 = 7'h32 == out_payload_2_rob_idx[6:0] ? rob_egress_id_50 : _GEN_12348; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12350 = 7'h33 == out_payload_2_rob_idx[6:0] ? rob_egress_id_51 : _GEN_12349; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12351 = 7'h34 == out_payload_2_rob_idx[6:0] ? rob_egress_id_52 : _GEN_12350; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12352 = 7'h35 == out_payload_2_rob_idx[6:0] ? rob_egress_id_53 : _GEN_12351; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12353 = 7'h36 == out_payload_2_rob_idx[6:0] ? rob_egress_id_54 : _GEN_12352; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12354 = 7'h37 == out_payload_2_rob_idx[6:0] ? rob_egress_id_55 : _GEN_12353; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12355 = 7'h38 == out_payload_2_rob_idx[6:0] ? rob_egress_id_56 : _GEN_12354; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12356 = 7'h39 == out_payload_2_rob_idx[6:0] ? rob_egress_id_57 : _GEN_12355; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12357 = 7'h3a == out_payload_2_rob_idx[6:0] ? rob_egress_id_58 : _GEN_12356; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12358 = 7'h3b == out_payload_2_rob_idx[6:0] ? rob_egress_id_59 : _GEN_12357; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12359 = 7'h3c == out_payload_2_rob_idx[6:0] ? rob_egress_id_60 : _GEN_12358; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12360 = 7'h3d == out_payload_2_rob_idx[6:0] ? rob_egress_id_61 : _GEN_12359; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12361 = 7'h3e == out_payload_2_rob_idx[6:0] ? rob_egress_id_62 : _GEN_12360; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12362 = 7'h3f == out_payload_2_rob_idx[6:0] ? rob_egress_id_63 : _GEN_12361; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12363 = 7'h40 == out_payload_2_rob_idx[6:0] ? rob_egress_id_64 : _GEN_12362; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12364 = 7'h41 == out_payload_2_rob_idx[6:0] ? rob_egress_id_65 : _GEN_12363; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12365 = 7'h42 == out_payload_2_rob_idx[6:0] ? rob_egress_id_66 : _GEN_12364; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12366 = 7'h43 == out_payload_2_rob_idx[6:0] ? rob_egress_id_67 : _GEN_12365; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12367 = 7'h44 == out_payload_2_rob_idx[6:0] ? rob_egress_id_68 : _GEN_12366; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12368 = 7'h45 == out_payload_2_rob_idx[6:0] ? rob_egress_id_69 : _GEN_12367; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12369 = 7'h46 == out_payload_2_rob_idx[6:0] ? rob_egress_id_70 : _GEN_12368; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12370 = 7'h47 == out_payload_2_rob_idx[6:0] ? rob_egress_id_71 : _GEN_12369; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12371 = 7'h48 == out_payload_2_rob_idx[6:0] ? rob_egress_id_72 : _GEN_12370; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12372 = 7'h49 == out_payload_2_rob_idx[6:0] ? rob_egress_id_73 : _GEN_12371; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12373 = 7'h4a == out_payload_2_rob_idx[6:0] ? rob_egress_id_74 : _GEN_12372; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12374 = 7'h4b == out_payload_2_rob_idx[6:0] ? rob_egress_id_75 : _GEN_12373; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12375 = 7'h4c == out_payload_2_rob_idx[6:0] ? rob_egress_id_76 : _GEN_12374; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12376 = 7'h4d == out_payload_2_rob_idx[6:0] ? rob_egress_id_77 : _GEN_12375; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12377 = 7'h4e == out_payload_2_rob_idx[6:0] ? rob_egress_id_78 : _GEN_12376; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12378 = 7'h4f == out_payload_2_rob_idx[6:0] ? rob_egress_id_79 : _GEN_12377; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12379 = 7'h50 == out_payload_2_rob_idx[6:0] ? rob_egress_id_80 : _GEN_12378; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12380 = 7'h51 == out_payload_2_rob_idx[6:0] ? rob_egress_id_81 : _GEN_12379; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12381 = 7'h52 == out_payload_2_rob_idx[6:0] ? rob_egress_id_82 : _GEN_12380; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12382 = 7'h53 == out_payload_2_rob_idx[6:0] ? rob_egress_id_83 : _GEN_12381; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12383 = 7'h54 == out_payload_2_rob_idx[6:0] ? rob_egress_id_84 : _GEN_12382; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12384 = 7'h55 == out_payload_2_rob_idx[6:0] ? rob_egress_id_85 : _GEN_12383; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12385 = 7'h56 == out_payload_2_rob_idx[6:0] ? rob_egress_id_86 : _GEN_12384; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12386 = 7'h57 == out_payload_2_rob_idx[6:0] ? rob_egress_id_87 : _GEN_12385; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12387 = 7'h58 == out_payload_2_rob_idx[6:0] ? rob_egress_id_88 : _GEN_12386; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12388 = 7'h59 == out_payload_2_rob_idx[6:0] ? rob_egress_id_89 : _GEN_12387; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12389 = 7'h5a == out_payload_2_rob_idx[6:0] ? rob_egress_id_90 : _GEN_12388; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12390 = 7'h5b == out_payload_2_rob_idx[6:0] ? rob_egress_id_91 : _GEN_12389; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12391 = 7'h5c == out_payload_2_rob_idx[6:0] ? rob_egress_id_92 : _GEN_12390; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12392 = 7'h5d == out_payload_2_rob_idx[6:0] ? rob_egress_id_93 : _GEN_12391; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12393 = 7'h5e == out_payload_2_rob_idx[6:0] ? rob_egress_id_94 : _GEN_12392; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12394 = 7'h5f == out_payload_2_rob_idx[6:0] ? rob_egress_id_95 : _GEN_12393; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12395 = 7'h60 == out_payload_2_rob_idx[6:0] ? rob_egress_id_96 : _GEN_12394; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12396 = 7'h61 == out_payload_2_rob_idx[6:0] ? rob_egress_id_97 : _GEN_12395; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12397 = 7'h62 == out_payload_2_rob_idx[6:0] ? rob_egress_id_98 : _GEN_12396; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12398 = 7'h63 == out_payload_2_rob_idx[6:0] ? rob_egress_id_99 : _GEN_12397; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12399 = 7'h64 == out_payload_2_rob_idx[6:0] ? rob_egress_id_100 : _GEN_12398; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12400 = 7'h65 == out_payload_2_rob_idx[6:0] ? rob_egress_id_101 : _GEN_12399; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12401 = 7'h66 == out_payload_2_rob_idx[6:0] ? rob_egress_id_102 : _GEN_12400; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12402 = 7'h67 == out_payload_2_rob_idx[6:0] ? rob_egress_id_103 : _GEN_12401; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12403 = 7'h68 == out_payload_2_rob_idx[6:0] ? rob_egress_id_104 : _GEN_12402; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12404 = 7'h69 == out_payload_2_rob_idx[6:0] ? rob_egress_id_105 : _GEN_12403; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12405 = 7'h6a == out_payload_2_rob_idx[6:0] ? rob_egress_id_106 : _GEN_12404; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12406 = 7'h6b == out_payload_2_rob_idx[6:0] ? rob_egress_id_107 : _GEN_12405; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12407 = 7'h6c == out_payload_2_rob_idx[6:0] ? rob_egress_id_108 : _GEN_12406; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12408 = 7'h6d == out_payload_2_rob_idx[6:0] ? rob_egress_id_109 : _GEN_12407; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12409 = 7'h6e == out_payload_2_rob_idx[6:0] ? rob_egress_id_110 : _GEN_12408; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12410 = 7'h6f == out_payload_2_rob_idx[6:0] ? rob_egress_id_111 : _GEN_12409; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12411 = 7'h70 == out_payload_2_rob_idx[6:0] ? rob_egress_id_112 : _GEN_12410; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12412 = 7'h71 == out_payload_2_rob_idx[6:0] ? rob_egress_id_113 : _GEN_12411; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12413 = 7'h72 == out_payload_2_rob_idx[6:0] ? rob_egress_id_114 : _GEN_12412; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12414 = 7'h73 == out_payload_2_rob_idx[6:0] ? rob_egress_id_115 : _GEN_12413; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12415 = 7'h74 == out_payload_2_rob_idx[6:0] ? rob_egress_id_116 : _GEN_12414; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12416 = 7'h75 == out_payload_2_rob_idx[6:0] ? rob_egress_id_117 : _GEN_12415; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12417 = 7'h76 == out_payload_2_rob_idx[6:0] ? rob_egress_id_118 : _GEN_12416; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12418 = 7'h77 == out_payload_2_rob_idx[6:0] ? rob_egress_id_119 : _GEN_12417; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12419 = 7'h78 == out_payload_2_rob_idx[6:0] ? rob_egress_id_120 : _GEN_12418; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12420 = 7'h79 == out_payload_2_rob_idx[6:0] ? rob_egress_id_121 : _GEN_12419; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12421 = 7'h7a == out_payload_2_rob_idx[6:0] ? rob_egress_id_122 : _GEN_12420; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12422 = 7'h7b == out_payload_2_rob_idx[6:0] ? rob_egress_id_123 : _GEN_12421; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12423 = 7'h7c == out_payload_2_rob_idx[6:0] ? rob_egress_id_124 : _GEN_12422; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12424 = 7'h7d == out_payload_2_rob_idx[6:0] ? rob_egress_id_125 : _GEN_12423; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12425 = 7'h7e == out_payload_2_rob_idx[6:0] ? rob_egress_id_126 : _GEN_12424; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_12426 = 7'h7f == out_payload_2_rob_idx[6:0] ? rob_egress_id_127 : _GEN_12425; // @[TestHarness.scala 204:{18,18}]
  wire [3:0] _GEN_12428 = 7'h1 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_1 : rob_flits_returned_0; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12429 = 7'h2 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_2 : _GEN_12428; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12430 = 7'h3 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_3 : _GEN_12429; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12431 = 7'h4 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_4 : _GEN_12430; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12432 = 7'h5 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_5 : _GEN_12431; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12433 = 7'h6 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_6 : _GEN_12432; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12434 = 7'h7 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_7 : _GEN_12433; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12435 = 7'h8 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_8 : _GEN_12434; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12436 = 7'h9 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_9 : _GEN_12435; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12437 = 7'ha == out_payload_2_rob_idx[6:0] ? rob_flits_returned_10 : _GEN_12436; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12438 = 7'hb == out_payload_2_rob_idx[6:0] ? rob_flits_returned_11 : _GEN_12437; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12439 = 7'hc == out_payload_2_rob_idx[6:0] ? rob_flits_returned_12 : _GEN_12438; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12440 = 7'hd == out_payload_2_rob_idx[6:0] ? rob_flits_returned_13 : _GEN_12439; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12441 = 7'he == out_payload_2_rob_idx[6:0] ? rob_flits_returned_14 : _GEN_12440; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12442 = 7'hf == out_payload_2_rob_idx[6:0] ? rob_flits_returned_15 : _GEN_12441; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12443 = 7'h10 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_16 : _GEN_12442; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12444 = 7'h11 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_17 : _GEN_12443; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12445 = 7'h12 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_18 : _GEN_12444; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12446 = 7'h13 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_19 : _GEN_12445; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12447 = 7'h14 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_20 : _GEN_12446; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12448 = 7'h15 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_21 : _GEN_12447; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12449 = 7'h16 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_22 : _GEN_12448; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12450 = 7'h17 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_23 : _GEN_12449; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12451 = 7'h18 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_24 : _GEN_12450; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12452 = 7'h19 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_25 : _GEN_12451; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12453 = 7'h1a == out_payload_2_rob_idx[6:0] ? rob_flits_returned_26 : _GEN_12452; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12454 = 7'h1b == out_payload_2_rob_idx[6:0] ? rob_flits_returned_27 : _GEN_12453; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12455 = 7'h1c == out_payload_2_rob_idx[6:0] ? rob_flits_returned_28 : _GEN_12454; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12456 = 7'h1d == out_payload_2_rob_idx[6:0] ? rob_flits_returned_29 : _GEN_12455; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12457 = 7'h1e == out_payload_2_rob_idx[6:0] ? rob_flits_returned_30 : _GEN_12456; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12458 = 7'h1f == out_payload_2_rob_idx[6:0] ? rob_flits_returned_31 : _GEN_12457; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12459 = 7'h20 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_32 : _GEN_12458; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12460 = 7'h21 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_33 : _GEN_12459; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12461 = 7'h22 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_34 : _GEN_12460; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12462 = 7'h23 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_35 : _GEN_12461; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12463 = 7'h24 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_36 : _GEN_12462; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12464 = 7'h25 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_37 : _GEN_12463; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12465 = 7'h26 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_38 : _GEN_12464; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12466 = 7'h27 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_39 : _GEN_12465; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12467 = 7'h28 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_40 : _GEN_12466; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12468 = 7'h29 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_41 : _GEN_12467; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12469 = 7'h2a == out_payload_2_rob_idx[6:0] ? rob_flits_returned_42 : _GEN_12468; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12470 = 7'h2b == out_payload_2_rob_idx[6:0] ? rob_flits_returned_43 : _GEN_12469; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12471 = 7'h2c == out_payload_2_rob_idx[6:0] ? rob_flits_returned_44 : _GEN_12470; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12472 = 7'h2d == out_payload_2_rob_idx[6:0] ? rob_flits_returned_45 : _GEN_12471; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12473 = 7'h2e == out_payload_2_rob_idx[6:0] ? rob_flits_returned_46 : _GEN_12472; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12474 = 7'h2f == out_payload_2_rob_idx[6:0] ? rob_flits_returned_47 : _GEN_12473; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12475 = 7'h30 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_48 : _GEN_12474; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12476 = 7'h31 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_49 : _GEN_12475; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12477 = 7'h32 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_50 : _GEN_12476; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12478 = 7'h33 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_51 : _GEN_12477; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12479 = 7'h34 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_52 : _GEN_12478; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12480 = 7'h35 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_53 : _GEN_12479; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12481 = 7'h36 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_54 : _GEN_12480; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12482 = 7'h37 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_55 : _GEN_12481; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12483 = 7'h38 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_56 : _GEN_12482; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12484 = 7'h39 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_57 : _GEN_12483; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12485 = 7'h3a == out_payload_2_rob_idx[6:0] ? rob_flits_returned_58 : _GEN_12484; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12486 = 7'h3b == out_payload_2_rob_idx[6:0] ? rob_flits_returned_59 : _GEN_12485; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12487 = 7'h3c == out_payload_2_rob_idx[6:0] ? rob_flits_returned_60 : _GEN_12486; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12488 = 7'h3d == out_payload_2_rob_idx[6:0] ? rob_flits_returned_61 : _GEN_12487; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12489 = 7'h3e == out_payload_2_rob_idx[6:0] ? rob_flits_returned_62 : _GEN_12488; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12490 = 7'h3f == out_payload_2_rob_idx[6:0] ? rob_flits_returned_63 : _GEN_12489; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12491 = 7'h40 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_64 : _GEN_12490; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12492 = 7'h41 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_65 : _GEN_12491; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12493 = 7'h42 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_66 : _GEN_12492; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12494 = 7'h43 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_67 : _GEN_12493; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12495 = 7'h44 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_68 : _GEN_12494; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12496 = 7'h45 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_69 : _GEN_12495; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12497 = 7'h46 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_70 : _GEN_12496; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12498 = 7'h47 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_71 : _GEN_12497; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12499 = 7'h48 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_72 : _GEN_12498; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12500 = 7'h49 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_73 : _GEN_12499; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12501 = 7'h4a == out_payload_2_rob_idx[6:0] ? rob_flits_returned_74 : _GEN_12500; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12502 = 7'h4b == out_payload_2_rob_idx[6:0] ? rob_flits_returned_75 : _GEN_12501; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12503 = 7'h4c == out_payload_2_rob_idx[6:0] ? rob_flits_returned_76 : _GEN_12502; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12504 = 7'h4d == out_payload_2_rob_idx[6:0] ? rob_flits_returned_77 : _GEN_12503; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12505 = 7'h4e == out_payload_2_rob_idx[6:0] ? rob_flits_returned_78 : _GEN_12504; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12506 = 7'h4f == out_payload_2_rob_idx[6:0] ? rob_flits_returned_79 : _GEN_12505; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12507 = 7'h50 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_80 : _GEN_12506; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12508 = 7'h51 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_81 : _GEN_12507; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12509 = 7'h52 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_82 : _GEN_12508; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12510 = 7'h53 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_83 : _GEN_12509; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12511 = 7'h54 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_84 : _GEN_12510; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12512 = 7'h55 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_85 : _GEN_12511; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12513 = 7'h56 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_86 : _GEN_12512; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12514 = 7'h57 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_87 : _GEN_12513; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12515 = 7'h58 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_88 : _GEN_12514; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12516 = 7'h59 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_89 : _GEN_12515; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12517 = 7'h5a == out_payload_2_rob_idx[6:0] ? rob_flits_returned_90 : _GEN_12516; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12518 = 7'h5b == out_payload_2_rob_idx[6:0] ? rob_flits_returned_91 : _GEN_12517; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12519 = 7'h5c == out_payload_2_rob_idx[6:0] ? rob_flits_returned_92 : _GEN_12518; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12520 = 7'h5d == out_payload_2_rob_idx[6:0] ? rob_flits_returned_93 : _GEN_12519; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12521 = 7'h5e == out_payload_2_rob_idx[6:0] ? rob_flits_returned_94 : _GEN_12520; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12522 = 7'h5f == out_payload_2_rob_idx[6:0] ? rob_flits_returned_95 : _GEN_12521; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12523 = 7'h60 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_96 : _GEN_12522; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12524 = 7'h61 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_97 : _GEN_12523; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12525 = 7'h62 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_98 : _GEN_12524; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12526 = 7'h63 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_99 : _GEN_12525; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12527 = 7'h64 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_100 : _GEN_12526; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12528 = 7'h65 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_101 : _GEN_12527; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12529 = 7'h66 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_102 : _GEN_12528; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12530 = 7'h67 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_103 : _GEN_12529; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12531 = 7'h68 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_104 : _GEN_12530; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12532 = 7'h69 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_105 : _GEN_12531; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12533 = 7'h6a == out_payload_2_rob_idx[6:0] ? rob_flits_returned_106 : _GEN_12532; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12534 = 7'h6b == out_payload_2_rob_idx[6:0] ? rob_flits_returned_107 : _GEN_12533; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12535 = 7'h6c == out_payload_2_rob_idx[6:0] ? rob_flits_returned_108 : _GEN_12534; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12536 = 7'h6d == out_payload_2_rob_idx[6:0] ? rob_flits_returned_109 : _GEN_12535; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12537 = 7'h6e == out_payload_2_rob_idx[6:0] ? rob_flits_returned_110 : _GEN_12536; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12538 = 7'h6f == out_payload_2_rob_idx[6:0] ? rob_flits_returned_111 : _GEN_12537; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12539 = 7'h70 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_112 : _GEN_12538; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12540 = 7'h71 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_113 : _GEN_12539; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12541 = 7'h72 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_114 : _GEN_12540; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12542 = 7'h73 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_115 : _GEN_12541; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12543 = 7'h74 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_116 : _GEN_12542; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12544 = 7'h75 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_117 : _GEN_12543; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12545 = 7'h76 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_118 : _GEN_12544; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12546 = 7'h77 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_119 : _GEN_12545; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12547 = 7'h78 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_120 : _GEN_12546; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12548 = 7'h79 == out_payload_2_rob_idx[6:0] ? rob_flits_returned_121 : _GEN_12547; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12549 = 7'h7a == out_payload_2_rob_idx[6:0] ? rob_flits_returned_122 : _GEN_12548; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12550 = 7'h7b == out_payload_2_rob_idx[6:0] ? rob_flits_returned_123 : _GEN_12549; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12551 = 7'h7c == out_payload_2_rob_idx[6:0] ? rob_flits_returned_124 : _GEN_12550; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12552 = 7'h7d == out_payload_2_rob_idx[6:0] ? rob_flits_returned_125 : _GEN_12551; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12553 = 7'h7e == out_payload_2_rob_idx[6:0] ? rob_flits_returned_126 : _GEN_12552; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12554 = 7'h7f == out_payload_2_rob_idx[6:0] ? rob_flits_returned_127 : _GEN_12553; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12556 = 7'h1 == out_payload_2_rob_idx[6:0] ? rob_n_flits_1 : rob_n_flits_0; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12557 = 7'h2 == out_payload_2_rob_idx[6:0] ? rob_n_flits_2 : _GEN_12556; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12558 = 7'h3 == out_payload_2_rob_idx[6:0] ? rob_n_flits_3 : _GEN_12557; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12559 = 7'h4 == out_payload_2_rob_idx[6:0] ? rob_n_flits_4 : _GEN_12558; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12560 = 7'h5 == out_payload_2_rob_idx[6:0] ? rob_n_flits_5 : _GEN_12559; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12561 = 7'h6 == out_payload_2_rob_idx[6:0] ? rob_n_flits_6 : _GEN_12560; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12562 = 7'h7 == out_payload_2_rob_idx[6:0] ? rob_n_flits_7 : _GEN_12561; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12563 = 7'h8 == out_payload_2_rob_idx[6:0] ? rob_n_flits_8 : _GEN_12562; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12564 = 7'h9 == out_payload_2_rob_idx[6:0] ? rob_n_flits_9 : _GEN_12563; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12565 = 7'ha == out_payload_2_rob_idx[6:0] ? rob_n_flits_10 : _GEN_12564; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12566 = 7'hb == out_payload_2_rob_idx[6:0] ? rob_n_flits_11 : _GEN_12565; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12567 = 7'hc == out_payload_2_rob_idx[6:0] ? rob_n_flits_12 : _GEN_12566; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12568 = 7'hd == out_payload_2_rob_idx[6:0] ? rob_n_flits_13 : _GEN_12567; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12569 = 7'he == out_payload_2_rob_idx[6:0] ? rob_n_flits_14 : _GEN_12568; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12570 = 7'hf == out_payload_2_rob_idx[6:0] ? rob_n_flits_15 : _GEN_12569; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12571 = 7'h10 == out_payload_2_rob_idx[6:0] ? rob_n_flits_16 : _GEN_12570; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12572 = 7'h11 == out_payload_2_rob_idx[6:0] ? rob_n_flits_17 : _GEN_12571; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12573 = 7'h12 == out_payload_2_rob_idx[6:0] ? rob_n_flits_18 : _GEN_12572; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12574 = 7'h13 == out_payload_2_rob_idx[6:0] ? rob_n_flits_19 : _GEN_12573; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12575 = 7'h14 == out_payload_2_rob_idx[6:0] ? rob_n_flits_20 : _GEN_12574; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12576 = 7'h15 == out_payload_2_rob_idx[6:0] ? rob_n_flits_21 : _GEN_12575; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12577 = 7'h16 == out_payload_2_rob_idx[6:0] ? rob_n_flits_22 : _GEN_12576; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12578 = 7'h17 == out_payload_2_rob_idx[6:0] ? rob_n_flits_23 : _GEN_12577; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12579 = 7'h18 == out_payload_2_rob_idx[6:0] ? rob_n_flits_24 : _GEN_12578; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12580 = 7'h19 == out_payload_2_rob_idx[6:0] ? rob_n_flits_25 : _GEN_12579; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12581 = 7'h1a == out_payload_2_rob_idx[6:0] ? rob_n_flits_26 : _GEN_12580; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12582 = 7'h1b == out_payload_2_rob_idx[6:0] ? rob_n_flits_27 : _GEN_12581; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12583 = 7'h1c == out_payload_2_rob_idx[6:0] ? rob_n_flits_28 : _GEN_12582; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12584 = 7'h1d == out_payload_2_rob_idx[6:0] ? rob_n_flits_29 : _GEN_12583; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12585 = 7'h1e == out_payload_2_rob_idx[6:0] ? rob_n_flits_30 : _GEN_12584; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12586 = 7'h1f == out_payload_2_rob_idx[6:0] ? rob_n_flits_31 : _GEN_12585; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12587 = 7'h20 == out_payload_2_rob_idx[6:0] ? rob_n_flits_32 : _GEN_12586; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12588 = 7'h21 == out_payload_2_rob_idx[6:0] ? rob_n_flits_33 : _GEN_12587; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12589 = 7'h22 == out_payload_2_rob_idx[6:0] ? rob_n_flits_34 : _GEN_12588; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12590 = 7'h23 == out_payload_2_rob_idx[6:0] ? rob_n_flits_35 : _GEN_12589; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12591 = 7'h24 == out_payload_2_rob_idx[6:0] ? rob_n_flits_36 : _GEN_12590; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12592 = 7'h25 == out_payload_2_rob_idx[6:0] ? rob_n_flits_37 : _GEN_12591; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12593 = 7'h26 == out_payload_2_rob_idx[6:0] ? rob_n_flits_38 : _GEN_12592; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12594 = 7'h27 == out_payload_2_rob_idx[6:0] ? rob_n_flits_39 : _GEN_12593; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12595 = 7'h28 == out_payload_2_rob_idx[6:0] ? rob_n_flits_40 : _GEN_12594; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12596 = 7'h29 == out_payload_2_rob_idx[6:0] ? rob_n_flits_41 : _GEN_12595; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12597 = 7'h2a == out_payload_2_rob_idx[6:0] ? rob_n_flits_42 : _GEN_12596; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12598 = 7'h2b == out_payload_2_rob_idx[6:0] ? rob_n_flits_43 : _GEN_12597; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12599 = 7'h2c == out_payload_2_rob_idx[6:0] ? rob_n_flits_44 : _GEN_12598; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12600 = 7'h2d == out_payload_2_rob_idx[6:0] ? rob_n_flits_45 : _GEN_12599; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12601 = 7'h2e == out_payload_2_rob_idx[6:0] ? rob_n_flits_46 : _GEN_12600; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12602 = 7'h2f == out_payload_2_rob_idx[6:0] ? rob_n_flits_47 : _GEN_12601; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12603 = 7'h30 == out_payload_2_rob_idx[6:0] ? rob_n_flits_48 : _GEN_12602; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12604 = 7'h31 == out_payload_2_rob_idx[6:0] ? rob_n_flits_49 : _GEN_12603; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12605 = 7'h32 == out_payload_2_rob_idx[6:0] ? rob_n_flits_50 : _GEN_12604; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12606 = 7'h33 == out_payload_2_rob_idx[6:0] ? rob_n_flits_51 : _GEN_12605; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12607 = 7'h34 == out_payload_2_rob_idx[6:0] ? rob_n_flits_52 : _GEN_12606; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12608 = 7'h35 == out_payload_2_rob_idx[6:0] ? rob_n_flits_53 : _GEN_12607; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12609 = 7'h36 == out_payload_2_rob_idx[6:0] ? rob_n_flits_54 : _GEN_12608; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12610 = 7'h37 == out_payload_2_rob_idx[6:0] ? rob_n_flits_55 : _GEN_12609; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12611 = 7'h38 == out_payload_2_rob_idx[6:0] ? rob_n_flits_56 : _GEN_12610; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12612 = 7'h39 == out_payload_2_rob_idx[6:0] ? rob_n_flits_57 : _GEN_12611; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12613 = 7'h3a == out_payload_2_rob_idx[6:0] ? rob_n_flits_58 : _GEN_12612; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12614 = 7'h3b == out_payload_2_rob_idx[6:0] ? rob_n_flits_59 : _GEN_12613; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12615 = 7'h3c == out_payload_2_rob_idx[6:0] ? rob_n_flits_60 : _GEN_12614; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12616 = 7'h3d == out_payload_2_rob_idx[6:0] ? rob_n_flits_61 : _GEN_12615; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12617 = 7'h3e == out_payload_2_rob_idx[6:0] ? rob_n_flits_62 : _GEN_12616; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12618 = 7'h3f == out_payload_2_rob_idx[6:0] ? rob_n_flits_63 : _GEN_12617; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12619 = 7'h40 == out_payload_2_rob_idx[6:0] ? rob_n_flits_64 : _GEN_12618; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12620 = 7'h41 == out_payload_2_rob_idx[6:0] ? rob_n_flits_65 : _GEN_12619; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12621 = 7'h42 == out_payload_2_rob_idx[6:0] ? rob_n_flits_66 : _GEN_12620; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12622 = 7'h43 == out_payload_2_rob_idx[6:0] ? rob_n_flits_67 : _GEN_12621; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12623 = 7'h44 == out_payload_2_rob_idx[6:0] ? rob_n_flits_68 : _GEN_12622; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12624 = 7'h45 == out_payload_2_rob_idx[6:0] ? rob_n_flits_69 : _GEN_12623; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12625 = 7'h46 == out_payload_2_rob_idx[6:0] ? rob_n_flits_70 : _GEN_12624; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12626 = 7'h47 == out_payload_2_rob_idx[6:0] ? rob_n_flits_71 : _GEN_12625; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12627 = 7'h48 == out_payload_2_rob_idx[6:0] ? rob_n_flits_72 : _GEN_12626; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12628 = 7'h49 == out_payload_2_rob_idx[6:0] ? rob_n_flits_73 : _GEN_12627; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12629 = 7'h4a == out_payload_2_rob_idx[6:0] ? rob_n_flits_74 : _GEN_12628; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12630 = 7'h4b == out_payload_2_rob_idx[6:0] ? rob_n_flits_75 : _GEN_12629; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12631 = 7'h4c == out_payload_2_rob_idx[6:0] ? rob_n_flits_76 : _GEN_12630; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12632 = 7'h4d == out_payload_2_rob_idx[6:0] ? rob_n_flits_77 : _GEN_12631; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12633 = 7'h4e == out_payload_2_rob_idx[6:0] ? rob_n_flits_78 : _GEN_12632; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12634 = 7'h4f == out_payload_2_rob_idx[6:0] ? rob_n_flits_79 : _GEN_12633; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12635 = 7'h50 == out_payload_2_rob_idx[6:0] ? rob_n_flits_80 : _GEN_12634; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12636 = 7'h51 == out_payload_2_rob_idx[6:0] ? rob_n_flits_81 : _GEN_12635; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12637 = 7'h52 == out_payload_2_rob_idx[6:0] ? rob_n_flits_82 : _GEN_12636; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12638 = 7'h53 == out_payload_2_rob_idx[6:0] ? rob_n_flits_83 : _GEN_12637; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12639 = 7'h54 == out_payload_2_rob_idx[6:0] ? rob_n_flits_84 : _GEN_12638; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12640 = 7'h55 == out_payload_2_rob_idx[6:0] ? rob_n_flits_85 : _GEN_12639; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12641 = 7'h56 == out_payload_2_rob_idx[6:0] ? rob_n_flits_86 : _GEN_12640; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12642 = 7'h57 == out_payload_2_rob_idx[6:0] ? rob_n_flits_87 : _GEN_12641; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12643 = 7'h58 == out_payload_2_rob_idx[6:0] ? rob_n_flits_88 : _GEN_12642; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12644 = 7'h59 == out_payload_2_rob_idx[6:0] ? rob_n_flits_89 : _GEN_12643; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12645 = 7'h5a == out_payload_2_rob_idx[6:0] ? rob_n_flits_90 : _GEN_12644; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12646 = 7'h5b == out_payload_2_rob_idx[6:0] ? rob_n_flits_91 : _GEN_12645; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12647 = 7'h5c == out_payload_2_rob_idx[6:0] ? rob_n_flits_92 : _GEN_12646; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12648 = 7'h5d == out_payload_2_rob_idx[6:0] ? rob_n_flits_93 : _GEN_12647; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12649 = 7'h5e == out_payload_2_rob_idx[6:0] ? rob_n_flits_94 : _GEN_12648; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12650 = 7'h5f == out_payload_2_rob_idx[6:0] ? rob_n_flits_95 : _GEN_12649; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12651 = 7'h60 == out_payload_2_rob_idx[6:0] ? rob_n_flits_96 : _GEN_12650; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12652 = 7'h61 == out_payload_2_rob_idx[6:0] ? rob_n_flits_97 : _GEN_12651; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12653 = 7'h62 == out_payload_2_rob_idx[6:0] ? rob_n_flits_98 : _GEN_12652; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12654 = 7'h63 == out_payload_2_rob_idx[6:0] ? rob_n_flits_99 : _GEN_12653; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12655 = 7'h64 == out_payload_2_rob_idx[6:0] ? rob_n_flits_100 : _GEN_12654; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12656 = 7'h65 == out_payload_2_rob_idx[6:0] ? rob_n_flits_101 : _GEN_12655; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12657 = 7'h66 == out_payload_2_rob_idx[6:0] ? rob_n_flits_102 : _GEN_12656; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12658 = 7'h67 == out_payload_2_rob_idx[6:0] ? rob_n_flits_103 : _GEN_12657; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12659 = 7'h68 == out_payload_2_rob_idx[6:0] ? rob_n_flits_104 : _GEN_12658; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12660 = 7'h69 == out_payload_2_rob_idx[6:0] ? rob_n_flits_105 : _GEN_12659; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12661 = 7'h6a == out_payload_2_rob_idx[6:0] ? rob_n_flits_106 : _GEN_12660; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12662 = 7'h6b == out_payload_2_rob_idx[6:0] ? rob_n_flits_107 : _GEN_12661; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12663 = 7'h6c == out_payload_2_rob_idx[6:0] ? rob_n_flits_108 : _GEN_12662; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12664 = 7'h6d == out_payload_2_rob_idx[6:0] ? rob_n_flits_109 : _GEN_12663; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12665 = 7'h6e == out_payload_2_rob_idx[6:0] ? rob_n_flits_110 : _GEN_12664; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12666 = 7'h6f == out_payload_2_rob_idx[6:0] ? rob_n_flits_111 : _GEN_12665; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12667 = 7'h70 == out_payload_2_rob_idx[6:0] ? rob_n_flits_112 : _GEN_12666; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12668 = 7'h71 == out_payload_2_rob_idx[6:0] ? rob_n_flits_113 : _GEN_12667; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12669 = 7'h72 == out_payload_2_rob_idx[6:0] ? rob_n_flits_114 : _GEN_12668; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12670 = 7'h73 == out_payload_2_rob_idx[6:0] ? rob_n_flits_115 : _GEN_12669; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12671 = 7'h74 == out_payload_2_rob_idx[6:0] ? rob_n_flits_116 : _GEN_12670; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12672 = 7'h75 == out_payload_2_rob_idx[6:0] ? rob_n_flits_117 : _GEN_12671; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12673 = 7'h76 == out_payload_2_rob_idx[6:0] ? rob_n_flits_118 : _GEN_12672; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12674 = 7'h77 == out_payload_2_rob_idx[6:0] ? rob_n_flits_119 : _GEN_12673; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12675 = 7'h78 == out_payload_2_rob_idx[6:0] ? rob_n_flits_120 : _GEN_12674; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12676 = 7'h79 == out_payload_2_rob_idx[6:0] ? rob_n_flits_121 : _GEN_12675; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12677 = 7'h7a == out_payload_2_rob_idx[6:0] ? rob_n_flits_122 : _GEN_12676; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12678 = 7'h7b == out_payload_2_rob_idx[6:0] ? rob_n_flits_123 : _GEN_12677; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12679 = 7'h7c == out_payload_2_rob_idx[6:0] ? rob_n_flits_124 : _GEN_12678; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12680 = 7'h7d == out_payload_2_rob_idx[6:0] ? rob_n_flits_125 : _GEN_12679; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12681 = 7'h7e == out_payload_2_rob_idx[6:0] ? rob_n_flits_126 : _GEN_12680; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_12682 = 7'h7f == out_payload_2_rob_idx[6:0] ? rob_n_flits_127 : _GEN_12681; // @[TestHarness.scala 205:{42,42}]
  wire [15:0] _GEN_15383 = {{9'd0}, packet_rob_idx_2}; // @[TestHarness.scala 206:61]
  wire  _T_204 = io_from_noc_2_flit_bits_head & enable_print_latency; // @[TestHarness.scala 208:30]
  wire [3:0] _rob_flits_returned_T_8 = _GEN_12554 + 4'h1; // @[TestHarness.scala 213:66]
  wire [3:0] _GEN_12939 = 7'h0 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11529; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12940 = 7'h1 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11530; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12941 = 7'h2 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11531; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12942 = 7'h3 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11532; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12943 = 7'h4 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11533; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12944 = 7'h5 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11534; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12945 = 7'h6 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11535; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12946 = 7'h7 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11536; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12947 = 7'h8 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11537; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12948 = 7'h9 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11538; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12949 = 7'ha == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11539; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12950 = 7'hb == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11540; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12951 = 7'hc == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11541; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12952 = 7'hd == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11542; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12953 = 7'he == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11543; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12954 = 7'hf == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11544; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12955 = 7'h10 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11545; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12956 = 7'h11 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11546; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12957 = 7'h12 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11547; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12958 = 7'h13 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11548; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12959 = 7'h14 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11549; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12960 = 7'h15 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11550; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12961 = 7'h16 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11551; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12962 = 7'h17 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11552; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12963 = 7'h18 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11553; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12964 = 7'h19 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11554; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12965 = 7'h1a == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11555; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12966 = 7'h1b == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11556; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12967 = 7'h1c == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11557; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12968 = 7'h1d == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11558; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12969 = 7'h1e == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11559; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12970 = 7'h1f == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11560; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12971 = 7'h20 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11561; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12972 = 7'h21 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11562; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12973 = 7'h22 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11563; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12974 = 7'h23 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11564; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12975 = 7'h24 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11565; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12976 = 7'h25 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11566; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12977 = 7'h26 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11567; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12978 = 7'h27 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11568; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12979 = 7'h28 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11569; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12980 = 7'h29 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11570; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12981 = 7'h2a == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11571; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12982 = 7'h2b == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11572; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12983 = 7'h2c == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11573; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12984 = 7'h2d == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11574; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12985 = 7'h2e == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11575; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12986 = 7'h2f == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11576; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12987 = 7'h30 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11577; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12988 = 7'h31 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11578; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12989 = 7'h32 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11579; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12990 = 7'h33 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11580; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12991 = 7'h34 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11581; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12992 = 7'h35 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11582; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12993 = 7'h36 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11583; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12994 = 7'h37 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11584; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12995 = 7'h38 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11585; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12996 = 7'h39 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11586; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12997 = 7'h3a == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11587; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12998 = 7'h3b == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11588; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_12999 = 7'h3c == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11589; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13000 = 7'h3d == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11590; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13001 = 7'h3e == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11591; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13002 = 7'h3f == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11592; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13003 = 7'h40 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11593; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13004 = 7'h41 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11594; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13005 = 7'h42 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11595; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13006 = 7'h43 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11596; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13007 = 7'h44 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11597; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13008 = 7'h45 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11598; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13009 = 7'h46 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11599; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13010 = 7'h47 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11600; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13011 = 7'h48 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11601; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13012 = 7'h49 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11602; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13013 = 7'h4a == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11603; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13014 = 7'h4b == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11604; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13015 = 7'h4c == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11605; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13016 = 7'h4d == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11606; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13017 = 7'h4e == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11607; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13018 = 7'h4f == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11608; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13019 = 7'h50 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11609; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13020 = 7'h51 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11610; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13021 = 7'h52 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11611; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13022 = 7'h53 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11612; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13023 = 7'h54 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11613; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13024 = 7'h55 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11614; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13025 = 7'h56 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11615; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13026 = 7'h57 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11616; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13027 = 7'h58 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11617; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13028 = 7'h59 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11618; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13029 = 7'h5a == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11619; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13030 = 7'h5b == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11620; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13031 = 7'h5c == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11621; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13032 = 7'h5d == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11622; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13033 = 7'h5e == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11623; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13034 = 7'h5f == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11624; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13035 = 7'h60 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11625; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13036 = 7'h61 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11626; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13037 = 7'h62 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11627; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13038 = 7'h63 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11628; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13039 = 7'h64 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11629; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13040 = 7'h65 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11630; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13041 = 7'h66 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11631; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13042 = 7'h67 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11632; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13043 = 7'h68 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11633; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13044 = 7'h69 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11634; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13045 = 7'h6a == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11635; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13046 = 7'h6b == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11636; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13047 = 7'h6c == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11637; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13048 = 7'h6d == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11638; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13049 = 7'h6e == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11639; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13050 = 7'h6f == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11640; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13051 = 7'h70 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11641; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13052 = 7'h71 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11642; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13053 = 7'h72 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11643; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13054 = 7'h73 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11644; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13055 = 7'h74 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11645; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13056 = 7'h75 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11646; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13057 = 7'h76 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11647; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13058 = 7'h77 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11648; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13059 = 7'h78 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11649; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13060 = 7'h79 == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11650; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13061 = 7'h7a == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11651; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13062 = 7'h7b == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11652; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13063 = 7'h7c == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11653; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13064 = 7'h7d == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11654; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13065 = 7'h7e == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11655; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_13066 = 7'h7f == out_payload_2_rob_idx[6:0] ? _rob_flits_returned_T_8 : _GEN_11656; // @[TestHarness.scala 213:{35,35}]
  wire [15:0] _rob_payload_flits_fired_T_8 = _GEN_12170 + 16'h1; // @[TestHarness.scala 214:76]
  wire [15:0] _GEN_13195 = 7'h0 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11657; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13196 = 7'h1 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11658; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13197 = 7'h2 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11659; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13198 = 7'h3 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11660; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13199 = 7'h4 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11661; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13200 = 7'h5 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11662; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13201 = 7'h6 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11663; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13202 = 7'h7 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11664; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13203 = 7'h8 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11665; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13204 = 7'h9 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11666; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13205 = 7'ha == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11667; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13206 = 7'hb == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11668; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13207 = 7'hc == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11669; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13208 = 7'hd == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11670; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13209 = 7'he == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11671; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13210 = 7'hf == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11672; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13211 = 7'h10 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11673; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13212 = 7'h11 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11674; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13213 = 7'h12 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11675; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13214 = 7'h13 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11676; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13215 = 7'h14 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11677; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13216 = 7'h15 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11678; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13217 = 7'h16 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11679; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13218 = 7'h17 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11680; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13219 = 7'h18 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11681; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13220 = 7'h19 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11682; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13221 = 7'h1a == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11683; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13222 = 7'h1b == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11684; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13223 = 7'h1c == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11685; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13224 = 7'h1d == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11686; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13225 = 7'h1e == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11687; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13226 = 7'h1f == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11688; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13227 = 7'h20 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11689; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13228 = 7'h21 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11690; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13229 = 7'h22 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11691; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13230 = 7'h23 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11692; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13231 = 7'h24 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11693; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13232 = 7'h25 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11694; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13233 = 7'h26 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11695; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13234 = 7'h27 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11696; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13235 = 7'h28 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11697; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13236 = 7'h29 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11698; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13237 = 7'h2a == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11699; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13238 = 7'h2b == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11700; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13239 = 7'h2c == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11701; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13240 = 7'h2d == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11702; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13241 = 7'h2e == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11703; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13242 = 7'h2f == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11704; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13243 = 7'h30 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11705; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13244 = 7'h31 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11706; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13245 = 7'h32 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11707; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13246 = 7'h33 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11708; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13247 = 7'h34 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11709; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13248 = 7'h35 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11710; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13249 = 7'h36 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11711; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13250 = 7'h37 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11712; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13251 = 7'h38 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11713; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13252 = 7'h39 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11714; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13253 = 7'h3a == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11715; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13254 = 7'h3b == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11716; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13255 = 7'h3c == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11717; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13256 = 7'h3d == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11718; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13257 = 7'h3e == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11719; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13258 = 7'h3f == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11720; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13259 = 7'h40 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11721; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13260 = 7'h41 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11722; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13261 = 7'h42 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11723; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13262 = 7'h43 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11724; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13263 = 7'h44 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11725; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13264 = 7'h45 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11726; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13265 = 7'h46 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11727; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13266 = 7'h47 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11728; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13267 = 7'h48 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11729; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13268 = 7'h49 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11730; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13269 = 7'h4a == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11731; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13270 = 7'h4b == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11732; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13271 = 7'h4c == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11733; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13272 = 7'h4d == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11734; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13273 = 7'h4e == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11735; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13274 = 7'h4f == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11736; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13275 = 7'h50 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11737; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13276 = 7'h51 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11738; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13277 = 7'h52 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11739; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13278 = 7'h53 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11740; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13279 = 7'h54 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11741; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13280 = 7'h55 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11742; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13281 = 7'h56 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11743; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13282 = 7'h57 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11744; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13283 = 7'h58 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11745; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13284 = 7'h59 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11746; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13285 = 7'h5a == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11747; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13286 = 7'h5b == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11748; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13287 = 7'h5c == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11749; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13288 = 7'h5d == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11750; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13289 = 7'h5e == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11751; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13290 = 7'h5f == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11752; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13291 = 7'h60 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11753; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13292 = 7'h61 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11754; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13293 = 7'h62 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11755; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13294 = 7'h63 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11756; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13295 = 7'h64 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11757; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13296 = 7'h65 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11758; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13297 = 7'h66 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11759; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13298 = 7'h67 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11760; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13299 = 7'h68 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11761; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13300 = 7'h69 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11762; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13301 = 7'h6a == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11763; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13302 = 7'h6b == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11764; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13303 = 7'h6c == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11765; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13304 = 7'h6d == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11766; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13305 = 7'h6e == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11767; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13306 = 7'h6f == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11768; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13307 = 7'h70 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11769; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13308 = 7'h71 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11770; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13309 = 7'h72 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11771; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13310 = 7'h73 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11772; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13311 = 7'h74 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11773; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13312 = 7'h75 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11774; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13313 = 7'h76 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11775; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13314 = 7'h77 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11776; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13315 = 7'h78 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11777; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13316 = 7'h79 == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11778; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13317 = 7'h7a == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11779; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13318 = 7'h7b == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11780; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13319 = 7'h7c == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11781; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13320 = 7'h7d == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11782; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13321 = 7'h7e == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11783; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_13322 = 7'h7f == out_payload_2_rob_idx[6:0] ? _rob_payload_flits_fired_T_8 : _GEN_11784; // @[TestHarness.scala 214:{40,40}]
  wire  _GEN_13323 = io_from_noc_2_flit_bits_head | packet_valid_2; // @[TestHarness.scala 196:31 215:{31,46}]
  wire [15:0] _GEN_13324 = io_from_noc_2_flit_bits_head ? out_payload_2_rob_idx : {{9'd0}, packet_rob_idx_2}; // @[TestHarness.scala 197:29 215:{31,72}]
  wire [3:0] _GEN_13326 = _T_212 ? _GEN_12939 : _GEN_11529; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13327 = _T_212 ? _GEN_12940 : _GEN_11530; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13328 = _T_212 ? _GEN_12941 : _GEN_11531; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13329 = _T_212 ? _GEN_12942 : _GEN_11532; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13330 = _T_212 ? _GEN_12943 : _GEN_11533; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13331 = _T_212 ? _GEN_12944 : _GEN_11534; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13332 = _T_212 ? _GEN_12945 : _GEN_11535; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13333 = _T_212 ? _GEN_12946 : _GEN_11536; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13334 = _T_212 ? _GEN_12947 : _GEN_11537; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13335 = _T_212 ? _GEN_12948 : _GEN_11538; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13336 = _T_212 ? _GEN_12949 : _GEN_11539; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13337 = _T_212 ? _GEN_12950 : _GEN_11540; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13338 = _T_212 ? _GEN_12951 : _GEN_11541; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13339 = _T_212 ? _GEN_12952 : _GEN_11542; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13340 = _T_212 ? _GEN_12953 : _GEN_11543; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13341 = _T_212 ? _GEN_12954 : _GEN_11544; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13342 = _T_212 ? _GEN_12955 : _GEN_11545; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13343 = _T_212 ? _GEN_12956 : _GEN_11546; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13344 = _T_212 ? _GEN_12957 : _GEN_11547; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13345 = _T_212 ? _GEN_12958 : _GEN_11548; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13346 = _T_212 ? _GEN_12959 : _GEN_11549; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13347 = _T_212 ? _GEN_12960 : _GEN_11550; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13348 = _T_212 ? _GEN_12961 : _GEN_11551; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13349 = _T_212 ? _GEN_12962 : _GEN_11552; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13350 = _T_212 ? _GEN_12963 : _GEN_11553; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13351 = _T_212 ? _GEN_12964 : _GEN_11554; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13352 = _T_212 ? _GEN_12965 : _GEN_11555; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13353 = _T_212 ? _GEN_12966 : _GEN_11556; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13354 = _T_212 ? _GEN_12967 : _GEN_11557; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13355 = _T_212 ? _GEN_12968 : _GEN_11558; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13356 = _T_212 ? _GEN_12969 : _GEN_11559; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13357 = _T_212 ? _GEN_12970 : _GEN_11560; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13358 = _T_212 ? _GEN_12971 : _GEN_11561; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13359 = _T_212 ? _GEN_12972 : _GEN_11562; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13360 = _T_212 ? _GEN_12973 : _GEN_11563; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13361 = _T_212 ? _GEN_12974 : _GEN_11564; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13362 = _T_212 ? _GEN_12975 : _GEN_11565; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13363 = _T_212 ? _GEN_12976 : _GEN_11566; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13364 = _T_212 ? _GEN_12977 : _GEN_11567; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13365 = _T_212 ? _GEN_12978 : _GEN_11568; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13366 = _T_212 ? _GEN_12979 : _GEN_11569; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13367 = _T_212 ? _GEN_12980 : _GEN_11570; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13368 = _T_212 ? _GEN_12981 : _GEN_11571; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13369 = _T_212 ? _GEN_12982 : _GEN_11572; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13370 = _T_212 ? _GEN_12983 : _GEN_11573; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13371 = _T_212 ? _GEN_12984 : _GEN_11574; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13372 = _T_212 ? _GEN_12985 : _GEN_11575; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13373 = _T_212 ? _GEN_12986 : _GEN_11576; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13374 = _T_212 ? _GEN_12987 : _GEN_11577; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13375 = _T_212 ? _GEN_12988 : _GEN_11578; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13376 = _T_212 ? _GEN_12989 : _GEN_11579; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13377 = _T_212 ? _GEN_12990 : _GEN_11580; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13378 = _T_212 ? _GEN_12991 : _GEN_11581; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13379 = _T_212 ? _GEN_12992 : _GEN_11582; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13380 = _T_212 ? _GEN_12993 : _GEN_11583; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13381 = _T_212 ? _GEN_12994 : _GEN_11584; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13382 = _T_212 ? _GEN_12995 : _GEN_11585; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13383 = _T_212 ? _GEN_12996 : _GEN_11586; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13384 = _T_212 ? _GEN_12997 : _GEN_11587; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13385 = _T_212 ? _GEN_12998 : _GEN_11588; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13386 = _T_212 ? _GEN_12999 : _GEN_11589; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13387 = _T_212 ? _GEN_13000 : _GEN_11590; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13388 = _T_212 ? _GEN_13001 : _GEN_11591; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13389 = _T_212 ? _GEN_13002 : _GEN_11592; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13390 = _T_212 ? _GEN_13003 : _GEN_11593; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13391 = _T_212 ? _GEN_13004 : _GEN_11594; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13392 = _T_212 ? _GEN_13005 : _GEN_11595; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13393 = _T_212 ? _GEN_13006 : _GEN_11596; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13394 = _T_212 ? _GEN_13007 : _GEN_11597; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13395 = _T_212 ? _GEN_13008 : _GEN_11598; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13396 = _T_212 ? _GEN_13009 : _GEN_11599; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13397 = _T_212 ? _GEN_13010 : _GEN_11600; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13398 = _T_212 ? _GEN_13011 : _GEN_11601; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13399 = _T_212 ? _GEN_13012 : _GEN_11602; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13400 = _T_212 ? _GEN_13013 : _GEN_11603; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13401 = _T_212 ? _GEN_13014 : _GEN_11604; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13402 = _T_212 ? _GEN_13015 : _GEN_11605; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13403 = _T_212 ? _GEN_13016 : _GEN_11606; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13404 = _T_212 ? _GEN_13017 : _GEN_11607; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13405 = _T_212 ? _GEN_13018 : _GEN_11608; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13406 = _T_212 ? _GEN_13019 : _GEN_11609; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13407 = _T_212 ? _GEN_13020 : _GEN_11610; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13408 = _T_212 ? _GEN_13021 : _GEN_11611; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13409 = _T_212 ? _GEN_13022 : _GEN_11612; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13410 = _T_212 ? _GEN_13023 : _GEN_11613; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13411 = _T_212 ? _GEN_13024 : _GEN_11614; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13412 = _T_212 ? _GEN_13025 : _GEN_11615; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13413 = _T_212 ? _GEN_13026 : _GEN_11616; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13414 = _T_212 ? _GEN_13027 : _GEN_11617; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13415 = _T_212 ? _GEN_13028 : _GEN_11618; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13416 = _T_212 ? _GEN_13029 : _GEN_11619; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13417 = _T_212 ? _GEN_13030 : _GEN_11620; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13418 = _T_212 ? _GEN_13031 : _GEN_11621; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13419 = _T_212 ? _GEN_13032 : _GEN_11622; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13420 = _T_212 ? _GEN_13033 : _GEN_11623; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13421 = _T_212 ? _GEN_13034 : _GEN_11624; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13422 = _T_212 ? _GEN_13035 : _GEN_11625; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13423 = _T_212 ? _GEN_13036 : _GEN_11626; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13424 = _T_212 ? _GEN_13037 : _GEN_11627; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13425 = _T_212 ? _GEN_13038 : _GEN_11628; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13426 = _T_212 ? _GEN_13039 : _GEN_11629; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13427 = _T_212 ? _GEN_13040 : _GEN_11630; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13428 = _T_212 ? _GEN_13041 : _GEN_11631; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13429 = _T_212 ? _GEN_13042 : _GEN_11632; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13430 = _T_212 ? _GEN_13043 : _GEN_11633; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13431 = _T_212 ? _GEN_13044 : _GEN_11634; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13432 = _T_212 ? _GEN_13045 : _GEN_11635; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13433 = _T_212 ? _GEN_13046 : _GEN_11636; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13434 = _T_212 ? _GEN_13047 : _GEN_11637; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13435 = _T_212 ? _GEN_13048 : _GEN_11638; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13436 = _T_212 ? _GEN_13049 : _GEN_11639; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13437 = _T_212 ? _GEN_13050 : _GEN_11640; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13438 = _T_212 ? _GEN_13051 : _GEN_11641; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13439 = _T_212 ? _GEN_13052 : _GEN_11642; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13440 = _T_212 ? _GEN_13053 : _GEN_11643; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13441 = _T_212 ? _GEN_13054 : _GEN_11644; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13442 = _T_212 ? _GEN_13055 : _GEN_11645; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13443 = _T_212 ? _GEN_13056 : _GEN_11646; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13444 = _T_212 ? _GEN_13057 : _GEN_11647; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13445 = _T_212 ? _GEN_13058 : _GEN_11648; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13446 = _T_212 ? _GEN_13059 : _GEN_11649; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13447 = _T_212 ? _GEN_13060 : _GEN_11650; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13448 = _T_212 ? _GEN_13061 : _GEN_11651; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13449 = _T_212 ? _GEN_13062 : _GEN_11652; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13450 = _T_212 ? _GEN_13063 : _GEN_11653; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13451 = _T_212 ? _GEN_13064 : _GEN_11654; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13452 = _T_212 ? _GEN_13065 : _GEN_11655; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_13453 = _T_212 ? _GEN_13066 : _GEN_11656; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13454 = _T_212 ? _GEN_13195 : _GEN_11657; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13455 = _T_212 ? _GEN_13196 : _GEN_11658; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13456 = _T_212 ? _GEN_13197 : _GEN_11659; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13457 = _T_212 ? _GEN_13198 : _GEN_11660; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13458 = _T_212 ? _GEN_13199 : _GEN_11661; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13459 = _T_212 ? _GEN_13200 : _GEN_11662; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13460 = _T_212 ? _GEN_13201 : _GEN_11663; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13461 = _T_212 ? _GEN_13202 : _GEN_11664; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13462 = _T_212 ? _GEN_13203 : _GEN_11665; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13463 = _T_212 ? _GEN_13204 : _GEN_11666; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13464 = _T_212 ? _GEN_13205 : _GEN_11667; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13465 = _T_212 ? _GEN_13206 : _GEN_11668; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13466 = _T_212 ? _GEN_13207 : _GEN_11669; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13467 = _T_212 ? _GEN_13208 : _GEN_11670; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13468 = _T_212 ? _GEN_13209 : _GEN_11671; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13469 = _T_212 ? _GEN_13210 : _GEN_11672; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13470 = _T_212 ? _GEN_13211 : _GEN_11673; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13471 = _T_212 ? _GEN_13212 : _GEN_11674; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13472 = _T_212 ? _GEN_13213 : _GEN_11675; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13473 = _T_212 ? _GEN_13214 : _GEN_11676; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13474 = _T_212 ? _GEN_13215 : _GEN_11677; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13475 = _T_212 ? _GEN_13216 : _GEN_11678; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13476 = _T_212 ? _GEN_13217 : _GEN_11679; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13477 = _T_212 ? _GEN_13218 : _GEN_11680; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13478 = _T_212 ? _GEN_13219 : _GEN_11681; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13479 = _T_212 ? _GEN_13220 : _GEN_11682; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13480 = _T_212 ? _GEN_13221 : _GEN_11683; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13481 = _T_212 ? _GEN_13222 : _GEN_11684; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13482 = _T_212 ? _GEN_13223 : _GEN_11685; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13483 = _T_212 ? _GEN_13224 : _GEN_11686; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13484 = _T_212 ? _GEN_13225 : _GEN_11687; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13485 = _T_212 ? _GEN_13226 : _GEN_11688; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13486 = _T_212 ? _GEN_13227 : _GEN_11689; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13487 = _T_212 ? _GEN_13228 : _GEN_11690; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13488 = _T_212 ? _GEN_13229 : _GEN_11691; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13489 = _T_212 ? _GEN_13230 : _GEN_11692; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13490 = _T_212 ? _GEN_13231 : _GEN_11693; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13491 = _T_212 ? _GEN_13232 : _GEN_11694; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13492 = _T_212 ? _GEN_13233 : _GEN_11695; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13493 = _T_212 ? _GEN_13234 : _GEN_11696; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13494 = _T_212 ? _GEN_13235 : _GEN_11697; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13495 = _T_212 ? _GEN_13236 : _GEN_11698; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13496 = _T_212 ? _GEN_13237 : _GEN_11699; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13497 = _T_212 ? _GEN_13238 : _GEN_11700; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13498 = _T_212 ? _GEN_13239 : _GEN_11701; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13499 = _T_212 ? _GEN_13240 : _GEN_11702; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13500 = _T_212 ? _GEN_13241 : _GEN_11703; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13501 = _T_212 ? _GEN_13242 : _GEN_11704; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13502 = _T_212 ? _GEN_13243 : _GEN_11705; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13503 = _T_212 ? _GEN_13244 : _GEN_11706; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13504 = _T_212 ? _GEN_13245 : _GEN_11707; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13505 = _T_212 ? _GEN_13246 : _GEN_11708; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13506 = _T_212 ? _GEN_13247 : _GEN_11709; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13507 = _T_212 ? _GEN_13248 : _GEN_11710; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13508 = _T_212 ? _GEN_13249 : _GEN_11711; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13509 = _T_212 ? _GEN_13250 : _GEN_11712; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13510 = _T_212 ? _GEN_13251 : _GEN_11713; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13511 = _T_212 ? _GEN_13252 : _GEN_11714; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13512 = _T_212 ? _GEN_13253 : _GEN_11715; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13513 = _T_212 ? _GEN_13254 : _GEN_11716; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13514 = _T_212 ? _GEN_13255 : _GEN_11717; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13515 = _T_212 ? _GEN_13256 : _GEN_11718; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13516 = _T_212 ? _GEN_13257 : _GEN_11719; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13517 = _T_212 ? _GEN_13258 : _GEN_11720; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13518 = _T_212 ? _GEN_13259 : _GEN_11721; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13519 = _T_212 ? _GEN_13260 : _GEN_11722; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13520 = _T_212 ? _GEN_13261 : _GEN_11723; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13521 = _T_212 ? _GEN_13262 : _GEN_11724; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13522 = _T_212 ? _GEN_13263 : _GEN_11725; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13523 = _T_212 ? _GEN_13264 : _GEN_11726; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13524 = _T_212 ? _GEN_13265 : _GEN_11727; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13525 = _T_212 ? _GEN_13266 : _GEN_11728; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13526 = _T_212 ? _GEN_13267 : _GEN_11729; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13527 = _T_212 ? _GEN_13268 : _GEN_11730; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13528 = _T_212 ? _GEN_13269 : _GEN_11731; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13529 = _T_212 ? _GEN_13270 : _GEN_11732; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13530 = _T_212 ? _GEN_13271 : _GEN_11733; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13531 = _T_212 ? _GEN_13272 : _GEN_11734; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13532 = _T_212 ? _GEN_13273 : _GEN_11735; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13533 = _T_212 ? _GEN_13274 : _GEN_11736; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13534 = _T_212 ? _GEN_13275 : _GEN_11737; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13535 = _T_212 ? _GEN_13276 : _GEN_11738; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13536 = _T_212 ? _GEN_13277 : _GEN_11739; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13537 = _T_212 ? _GEN_13278 : _GEN_11740; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13538 = _T_212 ? _GEN_13279 : _GEN_11741; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13539 = _T_212 ? _GEN_13280 : _GEN_11742; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13540 = _T_212 ? _GEN_13281 : _GEN_11743; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13541 = _T_212 ? _GEN_13282 : _GEN_11744; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13542 = _T_212 ? _GEN_13283 : _GEN_11745; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13543 = _T_212 ? _GEN_13284 : _GEN_11746; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13544 = _T_212 ? _GEN_13285 : _GEN_11747; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13545 = _T_212 ? _GEN_13286 : _GEN_11748; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13546 = _T_212 ? _GEN_13287 : _GEN_11749; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13547 = _T_212 ? _GEN_13288 : _GEN_11750; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13548 = _T_212 ? _GEN_13289 : _GEN_11751; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13549 = _T_212 ? _GEN_13290 : _GEN_11752; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13550 = _T_212 ? _GEN_13291 : _GEN_11753; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13551 = _T_212 ? _GEN_13292 : _GEN_11754; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13552 = _T_212 ? _GEN_13293 : _GEN_11755; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13553 = _T_212 ? _GEN_13294 : _GEN_11756; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13554 = _T_212 ? _GEN_13295 : _GEN_11757; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13555 = _T_212 ? _GEN_13296 : _GEN_11758; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13556 = _T_212 ? _GEN_13297 : _GEN_11759; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13557 = _T_212 ? _GEN_13298 : _GEN_11760; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13558 = _T_212 ? _GEN_13299 : _GEN_11761; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13559 = _T_212 ? _GEN_13300 : _GEN_11762; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13560 = _T_212 ? _GEN_13301 : _GEN_11763; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13561 = _T_212 ? _GEN_13302 : _GEN_11764; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13562 = _T_212 ? _GEN_13303 : _GEN_11765; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13563 = _T_212 ? _GEN_13304 : _GEN_11766; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13564 = _T_212 ? _GEN_13305 : _GEN_11767; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13565 = _T_212 ? _GEN_13306 : _GEN_11768; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13566 = _T_212 ? _GEN_13307 : _GEN_11769; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13567 = _T_212 ? _GEN_13308 : _GEN_11770; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13568 = _T_212 ? _GEN_13309 : _GEN_11771; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13569 = _T_212 ? _GEN_13310 : _GEN_11772; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13570 = _T_212 ? _GEN_13311 : _GEN_11773; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13571 = _T_212 ? _GEN_13312 : _GEN_11774; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13572 = _T_212 ? _GEN_13313 : _GEN_11775; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13573 = _T_212 ? _GEN_13314 : _GEN_11776; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13574 = _T_212 ? _GEN_13315 : _GEN_11777; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13575 = _T_212 ? _GEN_13316 : _GEN_11778; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13576 = _T_212 ? _GEN_13317 : _GEN_11779; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13577 = _T_212 ? _GEN_13318 : _GEN_11780; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13578 = _T_212 ? _GEN_13319 : _GEN_11781; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13579 = _T_212 ? _GEN_13320 : _GEN_11782; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13580 = _T_212 ? _GEN_13321 : _GEN_11783; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13581 = _T_212 ? _GEN_13322 : _GEN_11784; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_13583 = _T_212 ? _GEN_13324 : {{9'd0}, packet_rob_idx_2}; // @[TestHarness.scala 199:26 197:29]
  wire [31:0] out_payload_3_tsc = io_from_noc_3_flit_bits_payload[63:32]; // @[TestHarness.scala 194:51]
  reg  packet_valid_3; // @[TestHarness.scala 196:31]
  reg [6:0] packet_rob_idx_3; // @[TestHarness.scala 197:29]
  wire [127:0] _T_217 = rob_valids >> out_payload_3_rob_idx; // @[TestHarness.scala 201:24]
  wire [31:0] _GEN_13585 = 7'h1 == out_payload_3_rob_idx[6:0] ? rob_payload_1_tsc : rob_payload_0_tsc; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13586 = 7'h2 == out_payload_3_rob_idx[6:0] ? rob_payload_2_tsc : _GEN_13585; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13587 = 7'h3 == out_payload_3_rob_idx[6:0] ? rob_payload_3_tsc : _GEN_13586; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13588 = 7'h4 == out_payload_3_rob_idx[6:0] ? rob_payload_4_tsc : _GEN_13587; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13589 = 7'h5 == out_payload_3_rob_idx[6:0] ? rob_payload_5_tsc : _GEN_13588; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13590 = 7'h6 == out_payload_3_rob_idx[6:0] ? rob_payload_6_tsc : _GEN_13589; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13591 = 7'h7 == out_payload_3_rob_idx[6:0] ? rob_payload_7_tsc : _GEN_13590; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13592 = 7'h8 == out_payload_3_rob_idx[6:0] ? rob_payload_8_tsc : _GEN_13591; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13593 = 7'h9 == out_payload_3_rob_idx[6:0] ? rob_payload_9_tsc : _GEN_13592; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13594 = 7'ha == out_payload_3_rob_idx[6:0] ? rob_payload_10_tsc : _GEN_13593; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13595 = 7'hb == out_payload_3_rob_idx[6:0] ? rob_payload_11_tsc : _GEN_13594; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13596 = 7'hc == out_payload_3_rob_idx[6:0] ? rob_payload_12_tsc : _GEN_13595; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13597 = 7'hd == out_payload_3_rob_idx[6:0] ? rob_payload_13_tsc : _GEN_13596; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13598 = 7'he == out_payload_3_rob_idx[6:0] ? rob_payload_14_tsc : _GEN_13597; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13599 = 7'hf == out_payload_3_rob_idx[6:0] ? rob_payload_15_tsc : _GEN_13598; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13600 = 7'h10 == out_payload_3_rob_idx[6:0] ? rob_payload_16_tsc : _GEN_13599; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13601 = 7'h11 == out_payload_3_rob_idx[6:0] ? rob_payload_17_tsc : _GEN_13600; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13602 = 7'h12 == out_payload_3_rob_idx[6:0] ? rob_payload_18_tsc : _GEN_13601; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13603 = 7'h13 == out_payload_3_rob_idx[6:0] ? rob_payload_19_tsc : _GEN_13602; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13604 = 7'h14 == out_payload_3_rob_idx[6:0] ? rob_payload_20_tsc : _GEN_13603; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13605 = 7'h15 == out_payload_3_rob_idx[6:0] ? rob_payload_21_tsc : _GEN_13604; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13606 = 7'h16 == out_payload_3_rob_idx[6:0] ? rob_payload_22_tsc : _GEN_13605; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13607 = 7'h17 == out_payload_3_rob_idx[6:0] ? rob_payload_23_tsc : _GEN_13606; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13608 = 7'h18 == out_payload_3_rob_idx[6:0] ? rob_payload_24_tsc : _GEN_13607; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13609 = 7'h19 == out_payload_3_rob_idx[6:0] ? rob_payload_25_tsc : _GEN_13608; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13610 = 7'h1a == out_payload_3_rob_idx[6:0] ? rob_payload_26_tsc : _GEN_13609; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13611 = 7'h1b == out_payload_3_rob_idx[6:0] ? rob_payload_27_tsc : _GEN_13610; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13612 = 7'h1c == out_payload_3_rob_idx[6:0] ? rob_payload_28_tsc : _GEN_13611; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13613 = 7'h1d == out_payload_3_rob_idx[6:0] ? rob_payload_29_tsc : _GEN_13612; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13614 = 7'h1e == out_payload_3_rob_idx[6:0] ? rob_payload_30_tsc : _GEN_13613; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13615 = 7'h1f == out_payload_3_rob_idx[6:0] ? rob_payload_31_tsc : _GEN_13614; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13616 = 7'h20 == out_payload_3_rob_idx[6:0] ? rob_payload_32_tsc : _GEN_13615; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13617 = 7'h21 == out_payload_3_rob_idx[6:0] ? rob_payload_33_tsc : _GEN_13616; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13618 = 7'h22 == out_payload_3_rob_idx[6:0] ? rob_payload_34_tsc : _GEN_13617; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13619 = 7'h23 == out_payload_3_rob_idx[6:0] ? rob_payload_35_tsc : _GEN_13618; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13620 = 7'h24 == out_payload_3_rob_idx[6:0] ? rob_payload_36_tsc : _GEN_13619; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13621 = 7'h25 == out_payload_3_rob_idx[6:0] ? rob_payload_37_tsc : _GEN_13620; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13622 = 7'h26 == out_payload_3_rob_idx[6:0] ? rob_payload_38_tsc : _GEN_13621; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13623 = 7'h27 == out_payload_3_rob_idx[6:0] ? rob_payload_39_tsc : _GEN_13622; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13624 = 7'h28 == out_payload_3_rob_idx[6:0] ? rob_payload_40_tsc : _GEN_13623; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13625 = 7'h29 == out_payload_3_rob_idx[6:0] ? rob_payload_41_tsc : _GEN_13624; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13626 = 7'h2a == out_payload_3_rob_idx[6:0] ? rob_payload_42_tsc : _GEN_13625; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13627 = 7'h2b == out_payload_3_rob_idx[6:0] ? rob_payload_43_tsc : _GEN_13626; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13628 = 7'h2c == out_payload_3_rob_idx[6:0] ? rob_payload_44_tsc : _GEN_13627; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13629 = 7'h2d == out_payload_3_rob_idx[6:0] ? rob_payload_45_tsc : _GEN_13628; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13630 = 7'h2e == out_payload_3_rob_idx[6:0] ? rob_payload_46_tsc : _GEN_13629; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13631 = 7'h2f == out_payload_3_rob_idx[6:0] ? rob_payload_47_tsc : _GEN_13630; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13632 = 7'h30 == out_payload_3_rob_idx[6:0] ? rob_payload_48_tsc : _GEN_13631; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13633 = 7'h31 == out_payload_3_rob_idx[6:0] ? rob_payload_49_tsc : _GEN_13632; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13634 = 7'h32 == out_payload_3_rob_idx[6:0] ? rob_payload_50_tsc : _GEN_13633; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13635 = 7'h33 == out_payload_3_rob_idx[6:0] ? rob_payload_51_tsc : _GEN_13634; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13636 = 7'h34 == out_payload_3_rob_idx[6:0] ? rob_payload_52_tsc : _GEN_13635; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13637 = 7'h35 == out_payload_3_rob_idx[6:0] ? rob_payload_53_tsc : _GEN_13636; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13638 = 7'h36 == out_payload_3_rob_idx[6:0] ? rob_payload_54_tsc : _GEN_13637; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13639 = 7'h37 == out_payload_3_rob_idx[6:0] ? rob_payload_55_tsc : _GEN_13638; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13640 = 7'h38 == out_payload_3_rob_idx[6:0] ? rob_payload_56_tsc : _GEN_13639; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13641 = 7'h39 == out_payload_3_rob_idx[6:0] ? rob_payload_57_tsc : _GEN_13640; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13642 = 7'h3a == out_payload_3_rob_idx[6:0] ? rob_payload_58_tsc : _GEN_13641; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13643 = 7'h3b == out_payload_3_rob_idx[6:0] ? rob_payload_59_tsc : _GEN_13642; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13644 = 7'h3c == out_payload_3_rob_idx[6:0] ? rob_payload_60_tsc : _GEN_13643; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13645 = 7'h3d == out_payload_3_rob_idx[6:0] ? rob_payload_61_tsc : _GEN_13644; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13646 = 7'h3e == out_payload_3_rob_idx[6:0] ? rob_payload_62_tsc : _GEN_13645; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13647 = 7'h3f == out_payload_3_rob_idx[6:0] ? rob_payload_63_tsc : _GEN_13646; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13648 = 7'h40 == out_payload_3_rob_idx[6:0] ? rob_payload_64_tsc : _GEN_13647; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13649 = 7'h41 == out_payload_3_rob_idx[6:0] ? rob_payload_65_tsc : _GEN_13648; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13650 = 7'h42 == out_payload_3_rob_idx[6:0] ? rob_payload_66_tsc : _GEN_13649; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13651 = 7'h43 == out_payload_3_rob_idx[6:0] ? rob_payload_67_tsc : _GEN_13650; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13652 = 7'h44 == out_payload_3_rob_idx[6:0] ? rob_payload_68_tsc : _GEN_13651; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13653 = 7'h45 == out_payload_3_rob_idx[6:0] ? rob_payload_69_tsc : _GEN_13652; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13654 = 7'h46 == out_payload_3_rob_idx[6:0] ? rob_payload_70_tsc : _GEN_13653; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13655 = 7'h47 == out_payload_3_rob_idx[6:0] ? rob_payload_71_tsc : _GEN_13654; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13656 = 7'h48 == out_payload_3_rob_idx[6:0] ? rob_payload_72_tsc : _GEN_13655; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13657 = 7'h49 == out_payload_3_rob_idx[6:0] ? rob_payload_73_tsc : _GEN_13656; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13658 = 7'h4a == out_payload_3_rob_idx[6:0] ? rob_payload_74_tsc : _GEN_13657; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13659 = 7'h4b == out_payload_3_rob_idx[6:0] ? rob_payload_75_tsc : _GEN_13658; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13660 = 7'h4c == out_payload_3_rob_idx[6:0] ? rob_payload_76_tsc : _GEN_13659; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13661 = 7'h4d == out_payload_3_rob_idx[6:0] ? rob_payload_77_tsc : _GEN_13660; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13662 = 7'h4e == out_payload_3_rob_idx[6:0] ? rob_payload_78_tsc : _GEN_13661; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13663 = 7'h4f == out_payload_3_rob_idx[6:0] ? rob_payload_79_tsc : _GEN_13662; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13664 = 7'h50 == out_payload_3_rob_idx[6:0] ? rob_payload_80_tsc : _GEN_13663; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13665 = 7'h51 == out_payload_3_rob_idx[6:0] ? rob_payload_81_tsc : _GEN_13664; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13666 = 7'h52 == out_payload_3_rob_idx[6:0] ? rob_payload_82_tsc : _GEN_13665; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13667 = 7'h53 == out_payload_3_rob_idx[6:0] ? rob_payload_83_tsc : _GEN_13666; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13668 = 7'h54 == out_payload_3_rob_idx[6:0] ? rob_payload_84_tsc : _GEN_13667; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13669 = 7'h55 == out_payload_3_rob_idx[6:0] ? rob_payload_85_tsc : _GEN_13668; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13670 = 7'h56 == out_payload_3_rob_idx[6:0] ? rob_payload_86_tsc : _GEN_13669; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13671 = 7'h57 == out_payload_3_rob_idx[6:0] ? rob_payload_87_tsc : _GEN_13670; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13672 = 7'h58 == out_payload_3_rob_idx[6:0] ? rob_payload_88_tsc : _GEN_13671; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13673 = 7'h59 == out_payload_3_rob_idx[6:0] ? rob_payload_89_tsc : _GEN_13672; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13674 = 7'h5a == out_payload_3_rob_idx[6:0] ? rob_payload_90_tsc : _GEN_13673; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13675 = 7'h5b == out_payload_3_rob_idx[6:0] ? rob_payload_91_tsc : _GEN_13674; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13676 = 7'h5c == out_payload_3_rob_idx[6:0] ? rob_payload_92_tsc : _GEN_13675; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13677 = 7'h5d == out_payload_3_rob_idx[6:0] ? rob_payload_93_tsc : _GEN_13676; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13678 = 7'h5e == out_payload_3_rob_idx[6:0] ? rob_payload_94_tsc : _GEN_13677; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13679 = 7'h5f == out_payload_3_rob_idx[6:0] ? rob_payload_95_tsc : _GEN_13678; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13680 = 7'h60 == out_payload_3_rob_idx[6:0] ? rob_payload_96_tsc : _GEN_13679; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13681 = 7'h61 == out_payload_3_rob_idx[6:0] ? rob_payload_97_tsc : _GEN_13680; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13682 = 7'h62 == out_payload_3_rob_idx[6:0] ? rob_payload_98_tsc : _GEN_13681; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13683 = 7'h63 == out_payload_3_rob_idx[6:0] ? rob_payload_99_tsc : _GEN_13682; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13684 = 7'h64 == out_payload_3_rob_idx[6:0] ? rob_payload_100_tsc : _GEN_13683; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13685 = 7'h65 == out_payload_3_rob_idx[6:0] ? rob_payload_101_tsc : _GEN_13684; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13686 = 7'h66 == out_payload_3_rob_idx[6:0] ? rob_payload_102_tsc : _GEN_13685; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13687 = 7'h67 == out_payload_3_rob_idx[6:0] ? rob_payload_103_tsc : _GEN_13686; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13688 = 7'h68 == out_payload_3_rob_idx[6:0] ? rob_payload_104_tsc : _GEN_13687; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13689 = 7'h69 == out_payload_3_rob_idx[6:0] ? rob_payload_105_tsc : _GEN_13688; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13690 = 7'h6a == out_payload_3_rob_idx[6:0] ? rob_payload_106_tsc : _GEN_13689; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13691 = 7'h6b == out_payload_3_rob_idx[6:0] ? rob_payload_107_tsc : _GEN_13690; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13692 = 7'h6c == out_payload_3_rob_idx[6:0] ? rob_payload_108_tsc : _GEN_13691; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13693 = 7'h6d == out_payload_3_rob_idx[6:0] ? rob_payload_109_tsc : _GEN_13692; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13694 = 7'h6e == out_payload_3_rob_idx[6:0] ? rob_payload_110_tsc : _GEN_13693; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13695 = 7'h6f == out_payload_3_rob_idx[6:0] ? rob_payload_111_tsc : _GEN_13694; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13696 = 7'h70 == out_payload_3_rob_idx[6:0] ? rob_payload_112_tsc : _GEN_13695; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13697 = 7'h71 == out_payload_3_rob_idx[6:0] ? rob_payload_113_tsc : _GEN_13696; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13698 = 7'h72 == out_payload_3_rob_idx[6:0] ? rob_payload_114_tsc : _GEN_13697; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13699 = 7'h73 == out_payload_3_rob_idx[6:0] ? rob_payload_115_tsc : _GEN_13698; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13700 = 7'h74 == out_payload_3_rob_idx[6:0] ? rob_payload_116_tsc : _GEN_13699; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13701 = 7'h75 == out_payload_3_rob_idx[6:0] ? rob_payload_117_tsc : _GEN_13700; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13702 = 7'h76 == out_payload_3_rob_idx[6:0] ? rob_payload_118_tsc : _GEN_13701; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13703 = 7'h77 == out_payload_3_rob_idx[6:0] ? rob_payload_119_tsc : _GEN_13702; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13704 = 7'h78 == out_payload_3_rob_idx[6:0] ? rob_payload_120_tsc : _GEN_13703; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13705 = 7'h79 == out_payload_3_rob_idx[6:0] ? rob_payload_121_tsc : _GEN_13704; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13706 = 7'h7a == out_payload_3_rob_idx[6:0] ? rob_payload_122_tsc : _GEN_13705; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13707 = 7'h7b == out_payload_3_rob_idx[6:0] ? rob_payload_123_tsc : _GEN_13706; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13708 = 7'h7c == out_payload_3_rob_idx[6:0] ? rob_payload_124_tsc : _GEN_13707; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13709 = 7'h7d == out_payload_3_rob_idx[6:0] ? rob_payload_125_tsc : _GEN_13708; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13710 = 7'h7e == out_payload_3_rob_idx[6:0] ? rob_payload_126_tsc : _GEN_13709; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_13711 = 7'h7f == out_payload_3_rob_idx[6:0] ? rob_payload_127_tsc : _GEN_13710; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13713 = 7'h1 == out_payload_3_rob_idx[6:0] ? rob_payload_1_rob_idx : rob_payload_0_rob_idx; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13714 = 7'h2 == out_payload_3_rob_idx[6:0] ? rob_payload_2_rob_idx : _GEN_13713; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13715 = 7'h3 == out_payload_3_rob_idx[6:0] ? rob_payload_3_rob_idx : _GEN_13714; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13716 = 7'h4 == out_payload_3_rob_idx[6:0] ? rob_payload_4_rob_idx : _GEN_13715; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13717 = 7'h5 == out_payload_3_rob_idx[6:0] ? rob_payload_5_rob_idx : _GEN_13716; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13718 = 7'h6 == out_payload_3_rob_idx[6:0] ? rob_payload_6_rob_idx : _GEN_13717; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13719 = 7'h7 == out_payload_3_rob_idx[6:0] ? rob_payload_7_rob_idx : _GEN_13718; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13720 = 7'h8 == out_payload_3_rob_idx[6:0] ? rob_payload_8_rob_idx : _GEN_13719; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13721 = 7'h9 == out_payload_3_rob_idx[6:0] ? rob_payload_9_rob_idx : _GEN_13720; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13722 = 7'ha == out_payload_3_rob_idx[6:0] ? rob_payload_10_rob_idx : _GEN_13721; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13723 = 7'hb == out_payload_3_rob_idx[6:0] ? rob_payload_11_rob_idx : _GEN_13722; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13724 = 7'hc == out_payload_3_rob_idx[6:0] ? rob_payload_12_rob_idx : _GEN_13723; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13725 = 7'hd == out_payload_3_rob_idx[6:0] ? rob_payload_13_rob_idx : _GEN_13724; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13726 = 7'he == out_payload_3_rob_idx[6:0] ? rob_payload_14_rob_idx : _GEN_13725; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13727 = 7'hf == out_payload_3_rob_idx[6:0] ? rob_payload_15_rob_idx : _GEN_13726; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13728 = 7'h10 == out_payload_3_rob_idx[6:0] ? rob_payload_16_rob_idx : _GEN_13727; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13729 = 7'h11 == out_payload_3_rob_idx[6:0] ? rob_payload_17_rob_idx : _GEN_13728; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13730 = 7'h12 == out_payload_3_rob_idx[6:0] ? rob_payload_18_rob_idx : _GEN_13729; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13731 = 7'h13 == out_payload_3_rob_idx[6:0] ? rob_payload_19_rob_idx : _GEN_13730; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13732 = 7'h14 == out_payload_3_rob_idx[6:0] ? rob_payload_20_rob_idx : _GEN_13731; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13733 = 7'h15 == out_payload_3_rob_idx[6:0] ? rob_payload_21_rob_idx : _GEN_13732; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13734 = 7'h16 == out_payload_3_rob_idx[6:0] ? rob_payload_22_rob_idx : _GEN_13733; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13735 = 7'h17 == out_payload_3_rob_idx[6:0] ? rob_payload_23_rob_idx : _GEN_13734; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13736 = 7'h18 == out_payload_3_rob_idx[6:0] ? rob_payload_24_rob_idx : _GEN_13735; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13737 = 7'h19 == out_payload_3_rob_idx[6:0] ? rob_payload_25_rob_idx : _GEN_13736; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13738 = 7'h1a == out_payload_3_rob_idx[6:0] ? rob_payload_26_rob_idx : _GEN_13737; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13739 = 7'h1b == out_payload_3_rob_idx[6:0] ? rob_payload_27_rob_idx : _GEN_13738; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13740 = 7'h1c == out_payload_3_rob_idx[6:0] ? rob_payload_28_rob_idx : _GEN_13739; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13741 = 7'h1d == out_payload_3_rob_idx[6:0] ? rob_payload_29_rob_idx : _GEN_13740; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13742 = 7'h1e == out_payload_3_rob_idx[6:0] ? rob_payload_30_rob_idx : _GEN_13741; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13743 = 7'h1f == out_payload_3_rob_idx[6:0] ? rob_payload_31_rob_idx : _GEN_13742; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13744 = 7'h20 == out_payload_3_rob_idx[6:0] ? rob_payload_32_rob_idx : _GEN_13743; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13745 = 7'h21 == out_payload_3_rob_idx[6:0] ? rob_payload_33_rob_idx : _GEN_13744; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13746 = 7'h22 == out_payload_3_rob_idx[6:0] ? rob_payload_34_rob_idx : _GEN_13745; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13747 = 7'h23 == out_payload_3_rob_idx[6:0] ? rob_payload_35_rob_idx : _GEN_13746; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13748 = 7'h24 == out_payload_3_rob_idx[6:0] ? rob_payload_36_rob_idx : _GEN_13747; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13749 = 7'h25 == out_payload_3_rob_idx[6:0] ? rob_payload_37_rob_idx : _GEN_13748; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13750 = 7'h26 == out_payload_3_rob_idx[6:0] ? rob_payload_38_rob_idx : _GEN_13749; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13751 = 7'h27 == out_payload_3_rob_idx[6:0] ? rob_payload_39_rob_idx : _GEN_13750; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13752 = 7'h28 == out_payload_3_rob_idx[6:0] ? rob_payload_40_rob_idx : _GEN_13751; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13753 = 7'h29 == out_payload_3_rob_idx[6:0] ? rob_payload_41_rob_idx : _GEN_13752; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13754 = 7'h2a == out_payload_3_rob_idx[6:0] ? rob_payload_42_rob_idx : _GEN_13753; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13755 = 7'h2b == out_payload_3_rob_idx[6:0] ? rob_payload_43_rob_idx : _GEN_13754; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13756 = 7'h2c == out_payload_3_rob_idx[6:0] ? rob_payload_44_rob_idx : _GEN_13755; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13757 = 7'h2d == out_payload_3_rob_idx[6:0] ? rob_payload_45_rob_idx : _GEN_13756; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13758 = 7'h2e == out_payload_3_rob_idx[6:0] ? rob_payload_46_rob_idx : _GEN_13757; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13759 = 7'h2f == out_payload_3_rob_idx[6:0] ? rob_payload_47_rob_idx : _GEN_13758; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13760 = 7'h30 == out_payload_3_rob_idx[6:0] ? rob_payload_48_rob_idx : _GEN_13759; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13761 = 7'h31 == out_payload_3_rob_idx[6:0] ? rob_payload_49_rob_idx : _GEN_13760; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13762 = 7'h32 == out_payload_3_rob_idx[6:0] ? rob_payload_50_rob_idx : _GEN_13761; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13763 = 7'h33 == out_payload_3_rob_idx[6:0] ? rob_payload_51_rob_idx : _GEN_13762; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13764 = 7'h34 == out_payload_3_rob_idx[6:0] ? rob_payload_52_rob_idx : _GEN_13763; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13765 = 7'h35 == out_payload_3_rob_idx[6:0] ? rob_payload_53_rob_idx : _GEN_13764; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13766 = 7'h36 == out_payload_3_rob_idx[6:0] ? rob_payload_54_rob_idx : _GEN_13765; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13767 = 7'h37 == out_payload_3_rob_idx[6:0] ? rob_payload_55_rob_idx : _GEN_13766; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13768 = 7'h38 == out_payload_3_rob_idx[6:0] ? rob_payload_56_rob_idx : _GEN_13767; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13769 = 7'h39 == out_payload_3_rob_idx[6:0] ? rob_payload_57_rob_idx : _GEN_13768; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13770 = 7'h3a == out_payload_3_rob_idx[6:0] ? rob_payload_58_rob_idx : _GEN_13769; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13771 = 7'h3b == out_payload_3_rob_idx[6:0] ? rob_payload_59_rob_idx : _GEN_13770; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13772 = 7'h3c == out_payload_3_rob_idx[6:0] ? rob_payload_60_rob_idx : _GEN_13771; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13773 = 7'h3d == out_payload_3_rob_idx[6:0] ? rob_payload_61_rob_idx : _GEN_13772; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13774 = 7'h3e == out_payload_3_rob_idx[6:0] ? rob_payload_62_rob_idx : _GEN_13773; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13775 = 7'h3f == out_payload_3_rob_idx[6:0] ? rob_payload_63_rob_idx : _GEN_13774; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13776 = 7'h40 == out_payload_3_rob_idx[6:0] ? rob_payload_64_rob_idx : _GEN_13775; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13777 = 7'h41 == out_payload_3_rob_idx[6:0] ? rob_payload_65_rob_idx : _GEN_13776; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13778 = 7'h42 == out_payload_3_rob_idx[6:0] ? rob_payload_66_rob_idx : _GEN_13777; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13779 = 7'h43 == out_payload_3_rob_idx[6:0] ? rob_payload_67_rob_idx : _GEN_13778; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13780 = 7'h44 == out_payload_3_rob_idx[6:0] ? rob_payload_68_rob_idx : _GEN_13779; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13781 = 7'h45 == out_payload_3_rob_idx[6:0] ? rob_payload_69_rob_idx : _GEN_13780; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13782 = 7'h46 == out_payload_3_rob_idx[6:0] ? rob_payload_70_rob_idx : _GEN_13781; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13783 = 7'h47 == out_payload_3_rob_idx[6:0] ? rob_payload_71_rob_idx : _GEN_13782; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13784 = 7'h48 == out_payload_3_rob_idx[6:0] ? rob_payload_72_rob_idx : _GEN_13783; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13785 = 7'h49 == out_payload_3_rob_idx[6:0] ? rob_payload_73_rob_idx : _GEN_13784; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13786 = 7'h4a == out_payload_3_rob_idx[6:0] ? rob_payload_74_rob_idx : _GEN_13785; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13787 = 7'h4b == out_payload_3_rob_idx[6:0] ? rob_payload_75_rob_idx : _GEN_13786; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13788 = 7'h4c == out_payload_3_rob_idx[6:0] ? rob_payload_76_rob_idx : _GEN_13787; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13789 = 7'h4d == out_payload_3_rob_idx[6:0] ? rob_payload_77_rob_idx : _GEN_13788; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13790 = 7'h4e == out_payload_3_rob_idx[6:0] ? rob_payload_78_rob_idx : _GEN_13789; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13791 = 7'h4f == out_payload_3_rob_idx[6:0] ? rob_payload_79_rob_idx : _GEN_13790; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13792 = 7'h50 == out_payload_3_rob_idx[6:0] ? rob_payload_80_rob_idx : _GEN_13791; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13793 = 7'h51 == out_payload_3_rob_idx[6:0] ? rob_payload_81_rob_idx : _GEN_13792; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13794 = 7'h52 == out_payload_3_rob_idx[6:0] ? rob_payload_82_rob_idx : _GEN_13793; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13795 = 7'h53 == out_payload_3_rob_idx[6:0] ? rob_payload_83_rob_idx : _GEN_13794; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13796 = 7'h54 == out_payload_3_rob_idx[6:0] ? rob_payload_84_rob_idx : _GEN_13795; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13797 = 7'h55 == out_payload_3_rob_idx[6:0] ? rob_payload_85_rob_idx : _GEN_13796; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13798 = 7'h56 == out_payload_3_rob_idx[6:0] ? rob_payload_86_rob_idx : _GEN_13797; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13799 = 7'h57 == out_payload_3_rob_idx[6:0] ? rob_payload_87_rob_idx : _GEN_13798; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13800 = 7'h58 == out_payload_3_rob_idx[6:0] ? rob_payload_88_rob_idx : _GEN_13799; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13801 = 7'h59 == out_payload_3_rob_idx[6:0] ? rob_payload_89_rob_idx : _GEN_13800; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13802 = 7'h5a == out_payload_3_rob_idx[6:0] ? rob_payload_90_rob_idx : _GEN_13801; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13803 = 7'h5b == out_payload_3_rob_idx[6:0] ? rob_payload_91_rob_idx : _GEN_13802; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13804 = 7'h5c == out_payload_3_rob_idx[6:0] ? rob_payload_92_rob_idx : _GEN_13803; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13805 = 7'h5d == out_payload_3_rob_idx[6:0] ? rob_payload_93_rob_idx : _GEN_13804; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13806 = 7'h5e == out_payload_3_rob_idx[6:0] ? rob_payload_94_rob_idx : _GEN_13805; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13807 = 7'h5f == out_payload_3_rob_idx[6:0] ? rob_payload_95_rob_idx : _GEN_13806; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13808 = 7'h60 == out_payload_3_rob_idx[6:0] ? rob_payload_96_rob_idx : _GEN_13807; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13809 = 7'h61 == out_payload_3_rob_idx[6:0] ? rob_payload_97_rob_idx : _GEN_13808; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13810 = 7'h62 == out_payload_3_rob_idx[6:0] ? rob_payload_98_rob_idx : _GEN_13809; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13811 = 7'h63 == out_payload_3_rob_idx[6:0] ? rob_payload_99_rob_idx : _GEN_13810; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13812 = 7'h64 == out_payload_3_rob_idx[6:0] ? rob_payload_100_rob_idx : _GEN_13811; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13813 = 7'h65 == out_payload_3_rob_idx[6:0] ? rob_payload_101_rob_idx : _GEN_13812; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13814 = 7'h66 == out_payload_3_rob_idx[6:0] ? rob_payload_102_rob_idx : _GEN_13813; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13815 = 7'h67 == out_payload_3_rob_idx[6:0] ? rob_payload_103_rob_idx : _GEN_13814; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13816 = 7'h68 == out_payload_3_rob_idx[6:0] ? rob_payload_104_rob_idx : _GEN_13815; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13817 = 7'h69 == out_payload_3_rob_idx[6:0] ? rob_payload_105_rob_idx : _GEN_13816; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13818 = 7'h6a == out_payload_3_rob_idx[6:0] ? rob_payload_106_rob_idx : _GEN_13817; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13819 = 7'h6b == out_payload_3_rob_idx[6:0] ? rob_payload_107_rob_idx : _GEN_13818; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13820 = 7'h6c == out_payload_3_rob_idx[6:0] ? rob_payload_108_rob_idx : _GEN_13819; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13821 = 7'h6d == out_payload_3_rob_idx[6:0] ? rob_payload_109_rob_idx : _GEN_13820; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13822 = 7'h6e == out_payload_3_rob_idx[6:0] ? rob_payload_110_rob_idx : _GEN_13821; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13823 = 7'h6f == out_payload_3_rob_idx[6:0] ? rob_payload_111_rob_idx : _GEN_13822; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13824 = 7'h70 == out_payload_3_rob_idx[6:0] ? rob_payload_112_rob_idx : _GEN_13823; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13825 = 7'h71 == out_payload_3_rob_idx[6:0] ? rob_payload_113_rob_idx : _GEN_13824; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13826 = 7'h72 == out_payload_3_rob_idx[6:0] ? rob_payload_114_rob_idx : _GEN_13825; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13827 = 7'h73 == out_payload_3_rob_idx[6:0] ? rob_payload_115_rob_idx : _GEN_13826; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13828 = 7'h74 == out_payload_3_rob_idx[6:0] ? rob_payload_116_rob_idx : _GEN_13827; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13829 = 7'h75 == out_payload_3_rob_idx[6:0] ? rob_payload_117_rob_idx : _GEN_13828; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13830 = 7'h76 == out_payload_3_rob_idx[6:0] ? rob_payload_118_rob_idx : _GEN_13829; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13831 = 7'h77 == out_payload_3_rob_idx[6:0] ? rob_payload_119_rob_idx : _GEN_13830; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13832 = 7'h78 == out_payload_3_rob_idx[6:0] ? rob_payload_120_rob_idx : _GEN_13831; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13833 = 7'h79 == out_payload_3_rob_idx[6:0] ? rob_payload_121_rob_idx : _GEN_13832; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13834 = 7'h7a == out_payload_3_rob_idx[6:0] ? rob_payload_122_rob_idx : _GEN_13833; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13835 = 7'h7b == out_payload_3_rob_idx[6:0] ? rob_payload_123_rob_idx : _GEN_13834; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13836 = 7'h7c == out_payload_3_rob_idx[6:0] ? rob_payload_124_rob_idx : _GEN_13835; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13837 = 7'h7d == out_payload_3_rob_idx[6:0] ? rob_payload_125_rob_idx : _GEN_13836; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13838 = 7'h7e == out_payload_3_rob_idx[6:0] ? rob_payload_126_rob_idx : _GEN_13837; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13839 = 7'h7f == out_payload_3_rob_idx[6:0] ? rob_payload_127_rob_idx : _GEN_13838; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13841 = 7'h1 == out_payload_3_rob_idx[6:0] ? rob_payload_1_flits_fired : rob_payload_0_flits_fired; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13842 = 7'h2 == out_payload_3_rob_idx[6:0] ? rob_payload_2_flits_fired : _GEN_13841; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13843 = 7'h3 == out_payload_3_rob_idx[6:0] ? rob_payload_3_flits_fired : _GEN_13842; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13844 = 7'h4 == out_payload_3_rob_idx[6:0] ? rob_payload_4_flits_fired : _GEN_13843; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13845 = 7'h5 == out_payload_3_rob_idx[6:0] ? rob_payload_5_flits_fired : _GEN_13844; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13846 = 7'h6 == out_payload_3_rob_idx[6:0] ? rob_payload_6_flits_fired : _GEN_13845; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13847 = 7'h7 == out_payload_3_rob_idx[6:0] ? rob_payload_7_flits_fired : _GEN_13846; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13848 = 7'h8 == out_payload_3_rob_idx[6:0] ? rob_payload_8_flits_fired : _GEN_13847; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13849 = 7'h9 == out_payload_3_rob_idx[6:0] ? rob_payload_9_flits_fired : _GEN_13848; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13850 = 7'ha == out_payload_3_rob_idx[6:0] ? rob_payload_10_flits_fired : _GEN_13849; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13851 = 7'hb == out_payload_3_rob_idx[6:0] ? rob_payload_11_flits_fired : _GEN_13850; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13852 = 7'hc == out_payload_3_rob_idx[6:0] ? rob_payload_12_flits_fired : _GEN_13851; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13853 = 7'hd == out_payload_3_rob_idx[6:0] ? rob_payload_13_flits_fired : _GEN_13852; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13854 = 7'he == out_payload_3_rob_idx[6:0] ? rob_payload_14_flits_fired : _GEN_13853; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13855 = 7'hf == out_payload_3_rob_idx[6:0] ? rob_payload_15_flits_fired : _GEN_13854; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13856 = 7'h10 == out_payload_3_rob_idx[6:0] ? rob_payload_16_flits_fired : _GEN_13855; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13857 = 7'h11 == out_payload_3_rob_idx[6:0] ? rob_payload_17_flits_fired : _GEN_13856; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13858 = 7'h12 == out_payload_3_rob_idx[6:0] ? rob_payload_18_flits_fired : _GEN_13857; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13859 = 7'h13 == out_payload_3_rob_idx[6:0] ? rob_payload_19_flits_fired : _GEN_13858; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13860 = 7'h14 == out_payload_3_rob_idx[6:0] ? rob_payload_20_flits_fired : _GEN_13859; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13861 = 7'h15 == out_payload_3_rob_idx[6:0] ? rob_payload_21_flits_fired : _GEN_13860; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13862 = 7'h16 == out_payload_3_rob_idx[6:0] ? rob_payload_22_flits_fired : _GEN_13861; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13863 = 7'h17 == out_payload_3_rob_idx[6:0] ? rob_payload_23_flits_fired : _GEN_13862; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13864 = 7'h18 == out_payload_3_rob_idx[6:0] ? rob_payload_24_flits_fired : _GEN_13863; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13865 = 7'h19 == out_payload_3_rob_idx[6:0] ? rob_payload_25_flits_fired : _GEN_13864; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13866 = 7'h1a == out_payload_3_rob_idx[6:0] ? rob_payload_26_flits_fired : _GEN_13865; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13867 = 7'h1b == out_payload_3_rob_idx[6:0] ? rob_payload_27_flits_fired : _GEN_13866; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13868 = 7'h1c == out_payload_3_rob_idx[6:0] ? rob_payload_28_flits_fired : _GEN_13867; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13869 = 7'h1d == out_payload_3_rob_idx[6:0] ? rob_payload_29_flits_fired : _GEN_13868; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13870 = 7'h1e == out_payload_3_rob_idx[6:0] ? rob_payload_30_flits_fired : _GEN_13869; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13871 = 7'h1f == out_payload_3_rob_idx[6:0] ? rob_payload_31_flits_fired : _GEN_13870; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13872 = 7'h20 == out_payload_3_rob_idx[6:0] ? rob_payload_32_flits_fired : _GEN_13871; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13873 = 7'h21 == out_payload_3_rob_idx[6:0] ? rob_payload_33_flits_fired : _GEN_13872; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13874 = 7'h22 == out_payload_3_rob_idx[6:0] ? rob_payload_34_flits_fired : _GEN_13873; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13875 = 7'h23 == out_payload_3_rob_idx[6:0] ? rob_payload_35_flits_fired : _GEN_13874; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13876 = 7'h24 == out_payload_3_rob_idx[6:0] ? rob_payload_36_flits_fired : _GEN_13875; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13877 = 7'h25 == out_payload_3_rob_idx[6:0] ? rob_payload_37_flits_fired : _GEN_13876; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13878 = 7'h26 == out_payload_3_rob_idx[6:0] ? rob_payload_38_flits_fired : _GEN_13877; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13879 = 7'h27 == out_payload_3_rob_idx[6:0] ? rob_payload_39_flits_fired : _GEN_13878; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13880 = 7'h28 == out_payload_3_rob_idx[6:0] ? rob_payload_40_flits_fired : _GEN_13879; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13881 = 7'h29 == out_payload_3_rob_idx[6:0] ? rob_payload_41_flits_fired : _GEN_13880; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13882 = 7'h2a == out_payload_3_rob_idx[6:0] ? rob_payload_42_flits_fired : _GEN_13881; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13883 = 7'h2b == out_payload_3_rob_idx[6:0] ? rob_payload_43_flits_fired : _GEN_13882; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13884 = 7'h2c == out_payload_3_rob_idx[6:0] ? rob_payload_44_flits_fired : _GEN_13883; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13885 = 7'h2d == out_payload_3_rob_idx[6:0] ? rob_payload_45_flits_fired : _GEN_13884; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13886 = 7'h2e == out_payload_3_rob_idx[6:0] ? rob_payload_46_flits_fired : _GEN_13885; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13887 = 7'h2f == out_payload_3_rob_idx[6:0] ? rob_payload_47_flits_fired : _GEN_13886; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13888 = 7'h30 == out_payload_3_rob_idx[6:0] ? rob_payload_48_flits_fired : _GEN_13887; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13889 = 7'h31 == out_payload_3_rob_idx[6:0] ? rob_payload_49_flits_fired : _GEN_13888; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13890 = 7'h32 == out_payload_3_rob_idx[6:0] ? rob_payload_50_flits_fired : _GEN_13889; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13891 = 7'h33 == out_payload_3_rob_idx[6:0] ? rob_payload_51_flits_fired : _GEN_13890; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13892 = 7'h34 == out_payload_3_rob_idx[6:0] ? rob_payload_52_flits_fired : _GEN_13891; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13893 = 7'h35 == out_payload_3_rob_idx[6:0] ? rob_payload_53_flits_fired : _GEN_13892; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13894 = 7'h36 == out_payload_3_rob_idx[6:0] ? rob_payload_54_flits_fired : _GEN_13893; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13895 = 7'h37 == out_payload_3_rob_idx[6:0] ? rob_payload_55_flits_fired : _GEN_13894; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13896 = 7'h38 == out_payload_3_rob_idx[6:0] ? rob_payload_56_flits_fired : _GEN_13895; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13897 = 7'h39 == out_payload_3_rob_idx[6:0] ? rob_payload_57_flits_fired : _GEN_13896; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13898 = 7'h3a == out_payload_3_rob_idx[6:0] ? rob_payload_58_flits_fired : _GEN_13897; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13899 = 7'h3b == out_payload_3_rob_idx[6:0] ? rob_payload_59_flits_fired : _GEN_13898; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13900 = 7'h3c == out_payload_3_rob_idx[6:0] ? rob_payload_60_flits_fired : _GEN_13899; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13901 = 7'h3d == out_payload_3_rob_idx[6:0] ? rob_payload_61_flits_fired : _GEN_13900; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13902 = 7'h3e == out_payload_3_rob_idx[6:0] ? rob_payload_62_flits_fired : _GEN_13901; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13903 = 7'h3f == out_payload_3_rob_idx[6:0] ? rob_payload_63_flits_fired : _GEN_13902; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13904 = 7'h40 == out_payload_3_rob_idx[6:0] ? rob_payload_64_flits_fired : _GEN_13903; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13905 = 7'h41 == out_payload_3_rob_idx[6:0] ? rob_payload_65_flits_fired : _GEN_13904; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13906 = 7'h42 == out_payload_3_rob_idx[6:0] ? rob_payload_66_flits_fired : _GEN_13905; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13907 = 7'h43 == out_payload_3_rob_idx[6:0] ? rob_payload_67_flits_fired : _GEN_13906; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13908 = 7'h44 == out_payload_3_rob_idx[6:0] ? rob_payload_68_flits_fired : _GEN_13907; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13909 = 7'h45 == out_payload_3_rob_idx[6:0] ? rob_payload_69_flits_fired : _GEN_13908; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13910 = 7'h46 == out_payload_3_rob_idx[6:0] ? rob_payload_70_flits_fired : _GEN_13909; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13911 = 7'h47 == out_payload_3_rob_idx[6:0] ? rob_payload_71_flits_fired : _GEN_13910; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13912 = 7'h48 == out_payload_3_rob_idx[6:0] ? rob_payload_72_flits_fired : _GEN_13911; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13913 = 7'h49 == out_payload_3_rob_idx[6:0] ? rob_payload_73_flits_fired : _GEN_13912; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13914 = 7'h4a == out_payload_3_rob_idx[6:0] ? rob_payload_74_flits_fired : _GEN_13913; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13915 = 7'h4b == out_payload_3_rob_idx[6:0] ? rob_payload_75_flits_fired : _GEN_13914; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13916 = 7'h4c == out_payload_3_rob_idx[6:0] ? rob_payload_76_flits_fired : _GEN_13915; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13917 = 7'h4d == out_payload_3_rob_idx[6:0] ? rob_payload_77_flits_fired : _GEN_13916; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13918 = 7'h4e == out_payload_3_rob_idx[6:0] ? rob_payload_78_flits_fired : _GEN_13917; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13919 = 7'h4f == out_payload_3_rob_idx[6:0] ? rob_payload_79_flits_fired : _GEN_13918; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13920 = 7'h50 == out_payload_3_rob_idx[6:0] ? rob_payload_80_flits_fired : _GEN_13919; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13921 = 7'h51 == out_payload_3_rob_idx[6:0] ? rob_payload_81_flits_fired : _GEN_13920; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13922 = 7'h52 == out_payload_3_rob_idx[6:0] ? rob_payload_82_flits_fired : _GEN_13921; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13923 = 7'h53 == out_payload_3_rob_idx[6:0] ? rob_payload_83_flits_fired : _GEN_13922; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13924 = 7'h54 == out_payload_3_rob_idx[6:0] ? rob_payload_84_flits_fired : _GEN_13923; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13925 = 7'h55 == out_payload_3_rob_idx[6:0] ? rob_payload_85_flits_fired : _GEN_13924; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13926 = 7'h56 == out_payload_3_rob_idx[6:0] ? rob_payload_86_flits_fired : _GEN_13925; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13927 = 7'h57 == out_payload_3_rob_idx[6:0] ? rob_payload_87_flits_fired : _GEN_13926; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13928 = 7'h58 == out_payload_3_rob_idx[6:0] ? rob_payload_88_flits_fired : _GEN_13927; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13929 = 7'h59 == out_payload_3_rob_idx[6:0] ? rob_payload_89_flits_fired : _GEN_13928; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13930 = 7'h5a == out_payload_3_rob_idx[6:0] ? rob_payload_90_flits_fired : _GEN_13929; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13931 = 7'h5b == out_payload_3_rob_idx[6:0] ? rob_payload_91_flits_fired : _GEN_13930; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13932 = 7'h5c == out_payload_3_rob_idx[6:0] ? rob_payload_92_flits_fired : _GEN_13931; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13933 = 7'h5d == out_payload_3_rob_idx[6:0] ? rob_payload_93_flits_fired : _GEN_13932; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13934 = 7'h5e == out_payload_3_rob_idx[6:0] ? rob_payload_94_flits_fired : _GEN_13933; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13935 = 7'h5f == out_payload_3_rob_idx[6:0] ? rob_payload_95_flits_fired : _GEN_13934; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13936 = 7'h60 == out_payload_3_rob_idx[6:0] ? rob_payload_96_flits_fired : _GEN_13935; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13937 = 7'h61 == out_payload_3_rob_idx[6:0] ? rob_payload_97_flits_fired : _GEN_13936; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13938 = 7'h62 == out_payload_3_rob_idx[6:0] ? rob_payload_98_flits_fired : _GEN_13937; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13939 = 7'h63 == out_payload_3_rob_idx[6:0] ? rob_payload_99_flits_fired : _GEN_13938; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13940 = 7'h64 == out_payload_3_rob_idx[6:0] ? rob_payload_100_flits_fired : _GEN_13939; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13941 = 7'h65 == out_payload_3_rob_idx[6:0] ? rob_payload_101_flits_fired : _GEN_13940; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13942 = 7'h66 == out_payload_3_rob_idx[6:0] ? rob_payload_102_flits_fired : _GEN_13941; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13943 = 7'h67 == out_payload_3_rob_idx[6:0] ? rob_payload_103_flits_fired : _GEN_13942; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13944 = 7'h68 == out_payload_3_rob_idx[6:0] ? rob_payload_104_flits_fired : _GEN_13943; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13945 = 7'h69 == out_payload_3_rob_idx[6:0] ? rob_payload_105_flits_fired : _GEN_13944; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13946 = 7'h6a == out_payload_3_rob_idx[6:0] ? rob_payload_106_flits_fired : _GEN_13945; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13947 = 7'h6b == out_payload_3_rob_idx[6:0] ? rob_payload_107_flits_fired : _GEN_13946; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13948 = 7'h6c == out_payload_3_rob_idx[6:0] ? rob_payload_108_flits_fired : _GEN_13947; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13949 = 7'h6d == out_payload_3_rob_idx[6:0] ? rob_payload_109_flits_fired : _GEN_13948; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13950 = 7'h6e == out_payload_3_rob_idx[6:0] ? rob_payload_110_flits_fired : _GEN_13949; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13951 = 7'h6f == out_payload_3_rob_idx[6:0] ? rob_payload_111_flits_fired : _GEN_13950; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13952 = 7'h70 == out_payload_3_rob_idx[6:0] ? rob_payload_112_flits_fired : _GEN_13951; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13953 = 7'h71 == out_payload_3_rob_idx[6:0] ? rob_payload_113_flits_fired : _GEN_13952; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13954 = 7'h72 == out_payload_3_rob_idx[6:0] ? rob_payload_114_flits_fired : _GEN_13953; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13955 = 7'h73 == out_payload_3_rob_idx[6:0] ? rob_payload_115_flits_fired : _GEN_13954; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13956 = 7'h74 == out_payload_3_rob_idx[6:0] ? rob_payload_116_flits_fired : _GEN_13955; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13957 = 7'h75 == out_payload_3_rob_idx[6:0] ? rob_payload_117_flits_fired : _GEN_13956; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13958 = 7'h76 == out_payload_3_rob_idx[6:0] ? rob_payload_118_flits_fired : _GEN_13957; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13959 = 7'h77 == out_payload_3_rob_idx[6:0] ? rob_payload_119_flits_fired : _GEN_13958; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13960 = 7'h78 == out_payload_3_rob_idx[6:0] ? rob_payload_120_flits_fired : _GEN_13959; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13961 = 7'h79 == out_payload_3_rob_idx[6:0] ? rob_payload_121_flits_fired : _GEN_13960; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13962 = 7'h7a == out_payload_3_rob_idx[6:0] ? rob_payload_122_flits_fired : _GEN_13961; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13963 = 7'h7b == out_payload_3_rob_idx[6:0] ? rob_payload_123_flits_fired : _GEN_13962; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13964 = 7'h7c == out_payload_3_rob_idx[6:0] ? rob_payload_124_flits_fired : _GEN_13963; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13965 = 7'h7d == out_payload_3_rob_idx[6:0] ? rob_payload_125_flits_fired : _GEN_13964; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13966 = 7'h7e == out_payload_3_rob_idx[6:0] ? rob_payload_126_flits_fired : _GEN_13965; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_13967 = 7'h7f == out_payload_3_rob_idx[6:0] ? rob_payload_127_flits_fired : _GEN_13966; // @[TestHarness.scala 202:{35,35}]
  wire [63:0] _T_223 = {_GEN_13711,_GEN_13839,_GEN_13967}; // @[TestHarness.scala 202:35]
  wire [1:0] _GEN_13969 = 7'h1 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_1 : rob_ingress_id_0; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_13970 = 7'h2 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_2 : _GEN_13969; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_13971 = 7'h3 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_3 : _GEN_13970; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_13972 = 7'h4 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_4 : _GEN_13971; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_13973 = 7'h5 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_5 : _GEN_13972; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_13974 = 7'h6 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_6 : _GEN_13973; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_13975 = 7'h7 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_7 : _GEN_13974; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_13976 = 7'h8 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_8 : _GEN_13975; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_13977 = 7'h9 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_9 : _GEN_13976; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_13978 = 7'ha == out_payload_3_rob_idx[6:0] ? rob_ingress_id_10 : _GEN_13977; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_13979 = 7'hb == out_payload_3_rob_idx[6:0] ? rob_ingress_id_11 : _GEN_13978; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_13980 = 7'hc == out_payload_3_rob_idx[6:0] ? rob_ingress_id_12 : _GEN_13979; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_13981 = 7'hd == out_payload_3_rob_idx[6:0] ? rob_ingress_id_13 : _GEN_13980; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_13982 = 7'he == out_payload_3_rob_idx[6:0] ? rob_ingress_id_14 : _GEN_13981; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_13983 = 7'hf == out_payload_3_rob_idx[6:0] ? rob_ingress_id_15 : _GEN_13982; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_13984 = 7'h10 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_16 : _GEN_13983; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_13985 = 7'h11 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_17 : _GEN_13984; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_13986 = 7'h12 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_18 : _GEN_13985; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_13987 = 7'h13 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_19 : _GEN_13986; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_13988 = 7'h14 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_20 : _GEN_13987; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_13989 = 7'h15 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_21 : _GEN_13988; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_13990 = 7'h16 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_22 : _GEN_13989; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_13991 = 7'h17 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_23 : _GEN_13990; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_13992 = 7'h18 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_24 : _GEN_13991; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_13993 = 7'h19 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_25 : _GEN_13992; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_13994 = 7'h1a == out_payload_3_rob_idx[6:0] ? rob_ingress_id_26 : _GEN_13993; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_13995 = 7'h1b == out_payload_3_rob_idx[6:0] ? rob_ingress_id_27 : _GEN_13994; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_13996 = 7'h1c == out_payload_3_rob_idx[6:0] ? rob_ingress_id_28 : _GEN_13995; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_13997 = 7'h1d == out_payload_3_rob_idx[6:0] ? rob_ingress_id_29 : _GEN_13996; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_13998 = 7'h1e == out_payload_3_rob_idx[6:0] ? rob_ingress_id_30 : _GEN_13997; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_13999 = 7'h1f == out_payload_3_rob_idx[6:0] ? rob_ingress_id_31 : _GEN_13998; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14000 = 7'h20 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_32 : _GEN_13999; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14001 = 7'h21 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_33 : _GEN_14000; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14002 = 7'h22 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_34 : _GEN_14001; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14003 = 7'h23 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_35 : _GEN_14002; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14004 = 7'h24 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_36 : _GEN_14003; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14005 = 7'h25 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_37 : _GEN_14004; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14006 = 7'h26 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_38 : _GEN_14005; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14007 = 7'h27 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_39 : _GEN_14006; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14008 = 7'h28 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_40 : _GEN_14007; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14009 = 7'h29 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_41 : _GEN_14008; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14010 = 7'h2a == out_payload_3_rob_idx[6:0] ? rob_ingress_id_42 : _GEN_14009; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14011 = 7'h2b == out_payload_3_rob_idx[6:0] ? rob_ingress_id_43 : _GEN_14010; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14012 = 7'h2c == out_payload_3_rob_idx[6:0] ? rob_ingress_id_44 : _GEN_14011; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14013 = 7'h2d == out_payload_3_rob_idx[6:0] ? rob_ingress_id_45 : _GEN_14012; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14014 = 7'h2e == out_payload_3_rob_idx[6:0] ? rob_ingress_id_46 : _GEN_14013; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14015 = 7'h2f == out_payload_3_rob_idx[6:0] ? rob_ingress_id_47 : _GEN_14014; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14016 = 7'h30 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_48 : _GEN_14015; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14017 = 7'h31 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_49 : _GEN_14016; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14018 = 7'h32 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_50 : _GEN_14017; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14019 = 7'h33 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_51 : _GEN_14018; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14020 = 7'h34 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_52 : _GEN_14019; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14021 = 7'h35 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_53 : _GEN_14020; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14022 = 7'h36 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_54 : _GEN_14021; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14023 = 7'h37 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_55 : _GEN_14022; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14024 = 7'h38 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_56 : _GEN_14023; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14025 = 7'h39 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_57 : _GEN_14024; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14026 = 7'h3a == out_payload_3_rob_idx[6:0] ? rob_ingress_id_58 : _GEN_14025; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14027 = 7'h3b == out_payload_3_rob_idx[6:0] ? rob_ingress_id_59 : _GEN_14026; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14028 = 7'h3c == out_payload_3_rob_idx[6:0] ? rob_ingress_id_60 : _GEN_14027; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14029 = 7'h3d == out_payload_3_rob_idx[6:0] ? rob_ingress_id_61 : _GEN_14028; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14030 = 7'h3e == out_payload_3_rob_idx[6:0] ? rob_ingress_id_62 : _GEN_14029; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14031 = 7'h3f == out_payload_3_rob_idx[6:0] ? rob_ingress_id_63 : _GEN_14030; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14032 = 7'h40 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_64 : _GEN_14031; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14033 = 7'h41 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_65 : _GEN_14032; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14034 = 7'h42 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_66 : _GEN_14033; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14035 = 7'h43 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_67 : _GEN_14034; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14036 = 7'h44 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_68 : _GEN_14035; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14037 = 7'h45 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_69 : _GEN_14036; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14038 = 7'h46 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_70 : _GEN_14037; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14039 = 7'h47 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_71 : _GEN_14038; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14040 = 7'h48 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_72 : _GEN_14039; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14041 = 7'h49 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_73 : _GEN_14040; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14042 = 7'h4a == out_payload_3_rob_idx[6:0] ? rob_ingress_id_74 : _GEN_14041; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14043 = 7'h4b == out_payload_3_rob_idx[6:0] ? rob_ingress_id_75 : _GEN_14042; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14044 = 7'h4c == out_payload_3_rob_idx[6:0] ? rob_ingress_id_76 : _GEN_14043; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14045 = 7'h4d == out_payload_3_rob_idx[6:0] ? rob_ingress_id_77 : _GEN_14044; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14046 = 7'h4e == out_payload_3_rob_idx[6:0] ? rob_ingress_id_78 : _GEN_14045; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14047 = 7'h4f == out_payload_3_rob_idx[6:0] ? rob_ingress_id_79 : _GEN_14046; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14048 = 7'h50 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_80 : _GEN_14047; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14049 = 7'h51 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_81 : _GEN_14048; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14050 = 7'h52 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_82 : _GEN_14049; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14051 = 7'h53 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_83 : _GEN_14050; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14052 = 7'h54 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_84 : _GEN_14051; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14053 = 7'h55 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_85 : _GEN_14052; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14054 = 7'h56 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_86 : _GEN_14053; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14055 = 7'h57 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_87 : _GEN_14054; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14056 = 7'h58 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_88 : _GEN_14055; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14057 = 7'h59 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_89 : _GEN_14056; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14058 = 7'h5a == out_payload_3_rob_idx[6:0] ? rob_ingress_id_90 : _GEN_14057; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14059 = 7'h5b == out_payload_3_rob_idx[6:0] ? rob_ingress_id_91 : _GEN_14058; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14060 = 7'h5c == out_payload_3_rob_idx[6:0] ? rob_ingress_id_92 : _GEN_14059; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14061 = 7'h5d == out_payload_3_rob_idx[6:0] ? rob_ingress_id_93 : _GEN_14060; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14062 = 7'h5e == out_payload_3_rob_idx[6:0] ? rob_ingress_id_94 : _GEN_14061; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14063 = 7'h5f == out_payload_3_rob_idx[6:0] ? rob_ingress_id_95 : _GEN_14062; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14064 = 7'h60 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_96 : _GEN_14063; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14065 = 7'h61 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_97 : _GEN_14064; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14066 = 7'h62 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_98 : _GEN_14065; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14067 = 7'h63 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_99 : _GEN_14066; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14068 = 7'h64 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_100 : _GEN_14067; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14069 = 7'h65 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_101 : _GEN_14068; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14070 = 7'h66 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_102 : _GEN_14069; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14071 = 7'h67 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_103 : _GEN_14070; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14072 = 7'h68 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_104 : _GEN_14071; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14073 = 7'h69 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_105 : _GEN_14072; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14074 = 7'h6a == out_payload_3_rob_idx[6:0] ? rob_ingress_id_106 : _GEN_14073; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14075 = 7'h6b == out_payload_3_rob_idx[6:0] ? rob_ingress_id_107 : _GEN_14074; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14076 = 7'h6c == out_payload_3_rob_idx[6:0] ? rob_ingress_id_108 : _GEN_14075; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14077 = 7'h6d == out_payload_3_rob_idx[6:0] ? rob_ingress_id_109 : _GEN_14076; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14078 = 7'h6e == out_payload_3_rob_idx[6:0] ? rob_ingress_id_110 : _GEN_14077; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14079 = 7'h6f == out_payload_3_rob_idx[6:0] ? rob_ingress_id_111 : _GEN_14078; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14080 = 7'h70 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_112 : _GEN_14079; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14081 = 7'h71 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_113 : _GEN_14080; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14082 = 7'h72 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_114 : _GEN_14081; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14083 = 7'h73 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_115 : _GEN_14082; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14084 = 7'h74 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_116 : _GEN_14083; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14085 = 7'h75 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_117 : _GEN_14084; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14086 = 7'h76 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_118 : _GEN_14085; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14087 = 7'h77 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_119 : _GEN_14086; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14088 = 7'h78 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_120 : _GEN_14087; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14089 = 7'h79 == out_payload_3_rob_idx[6:0] ? rob_ingress_id_121 : _GEN_14088; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14090 = 7'h7a == out_payload_3_rob_idx[6:0] ? rob_ingress_id_122 : _GEN_14089; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14091 = 7'h7b == out_payload_3_rob_idx[6:0] ? rob_ingress_id_123 : _GEN_14090; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14092 = 7'h7c == out_payload_3_rob_idx[6:0] ? rob_ingress_id_124 : _GEN_14091; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14093 = 7'h7d == out_payload_3_rob_idx[6:0] ? rob_ingress_id_125 : _GEN_14092; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14094 = 7'h7e == out_payload_3_rob_idx[6:0] ? rob_ingress_id_126 : _GEN_14093; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14095 = 7'h7f == out_payload_3_rob_idx[6:0] ? rob_ingress_id_127 : _GEN_14094; // @[TestHarness.scala 203:{37,37}]
  wire [1:0] _GEN_14097 = 7'h1 == out_payload_3_rob_idx[6:0] ? rob_egress_id_1 : rob_egress_id_0; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14098 = 7'h2 == out_payload_3_rob_idx[6:0] ? rob_egress_id_2 : _GEN_14097; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14099 = 7'h3 == out_payload_3_rob_idx[6:0] ? rob_egress_id_3 : _GEN_14098; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14100 = 7'h4 == out_payload_3_rob_idx[6:0] ? rob_egress_id_4 : _GEN_14099; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14101 = 7'h5 == out_payload_3_rob_idx[6:0] ? rob_egress_id_5 : _GEN_14100; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14102 = 7'h6 == out_payload_3_rob_idx[6:0] ? rob_egress_id_6 : _GEN_14101; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14103 = 7'h7 == out_payload_3_rob_idx[6:0] ? rob_egress_id_7 : _GEN_14102; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14104 = 7'h8 == out_payload_3_rob_idx[6:0] ? rob_egress_id_8 : _GEN_14103; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14105 = 7'h9 == out_payload_3_rob_idx[6:0] ? rob_egress_id_9 : _GEN_14104; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14106 = 7'ha == out_payload_3_rob_idx[6:0] ? rob_egress_id_10 : _GEN_14105; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14107 = 7'hb == out_payload_3_rob_idx[6:0] ? rob_egress_id_11 : _GEN_14106; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14108 = 7'hc == out_payload_3_rob_idx[6:0] ? rob_egress_id_12 : _GEN_14107; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14109 = 7'hd == out_payload_3_rob_idx[6:0] ? rob_egress_id_13 : _GEN_14108; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14110 = 7'he == out_payload_3_rob_idx[6:0] ? rob_egress_id_14 : _GEN_14109; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14111 = 7'hf == out_payload_3_rob_idx[6:0] ? rob_egress_id_15 : _GEN_14110; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14112 = 7'h10 == out_payload_3_rob_idx[6:0] ? rob_egress_id_16 : _GEN_14111; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14113 = 7'h11 == out_payload_3_rob_idx[6:0] ? rob_egress_id_17 : _GEN_14112; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14114 = 7'h12 == out_payload_3_rob_idx[6:0] ? rob_egress_id_18 : _GEN_14113; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14115 = 7'h13 == out_payload_3_rob_idx[6:0] ? rob_egress_id_19 : _GEN_14114; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14116 = 7'h14 == out_payload_3_rob_idx[6:0] ? rob_egress_id_20 : _GEN_14115; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14117 = 7'h15 == out_payload_3_rob_idx[6:0] ? rob_egress_id_21 : _GEN_14116; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14118 = 7'h16 == out_payload_3_rob_idx[6:0] ? rob_egress_id_22 : _GEN_14117; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14119 = 7'h17 == out_payload_3_rob_idx[6:0] ? rob_egress_id_23 : _GEN_14118; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14120 = 7'h18 == out_payload_3_rob_idx[6:0] ? rob_egress_id_24 : _GEN_14119; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14121 = 7'h19 == out_payload_3_rob_idx[6:0] ? rob_egress_id_25 : _GEN_14120; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14122 = 7'h1a == out_payload_3_rob_idx[6:0] ? rob_egress_id_26 : _GEN_14121; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14123 = 7'h1b == out_payload_3_rob_idx[6:0] ? rob_egress_id_27 : _GEN_14122; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14124 = 7'h1c == out_payload_3_rob_idx[6:0] ? rob_egress_id_28 : _GEN_14123; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14125 = 7'h1d == out_payload_3_rob_idx[6:0] ? rob_egress_id_29 : _GEN_14124; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14126 = 7'h1e == out_payload_3_rob_idx[6:0] ? rob_egress_id_30 : _GEN_14125; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14127 = 7'h1f == out_payload_3_rob_idx[6:0] ? rob_egress_id_31 : _GEN_14126; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14128 = 7'h20 == out_payload_3_rob_idx[6:0] ? rob_egress_id_32 : _GEN_14127; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14129 = 7'h21 == out_payload_3_rob_idx[6:0] ? rob_egress_id_33 : _GEN_14128; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14130 = 7'h22 == out_payload_3_rob_idx[6:0] ? rob_egress_id_34 : _GEN_14129; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14131 = 7'h23 == out_payload_3_rob_idx[6:0] ? rob_egress_id_35 : _GEN_14130; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14132 = 7'h24 == out_payload_3_rob_idx[6:0] ? rob_egress_id_36 : _GEN_14131; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14133 = 7'h25 == out_payload_3_rob_idx[6:0] ? rob_egress_id_37 : _GEN_14132; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14134 = 7'h26 == out_payload_3_rob_idx[6:0] ? rob_egress_id_38 : _GEN_14133; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14135 = 7'h27 == out_payload_3_rob_idx[6:0] ? rob_egress_id_39 : _GEN_14134; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14136 = 7'h28 == out_payload_3_rob_idx[6:0] ? rob_egress_id_40 : _GEN_14135; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14137 = 7'h29 == out_payload_3_rob_idx[6:0] ? rob_egress_id_41 : _GEN_14136; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14138 = 7'h2a == out_payload_3_rob_idx[6:0] ? rob_egress_id_42 : _GEN_14137; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14139 = 7'h2b == out_payload_3_rob_idx[6:0] ? rob_egress_id_43 : _GEN_14138; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14140 = 7'h2c == out_payload_3_rob_idx[6:0] ? rob_egress_id_44 : _GEN_14139; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14141 = 7'h2d == out_payload_3_rob_idx[6:0] ? rob_egress_id_45 : _GEN_14140; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14142 = 7'h2e == out_payload_3_rob_idx[6:0] ? rob_egress_id_46 : _GEN_14141; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14143 = 7'h2f == out_payload_3_rob_idx[6:0] ? rob_egress_id_47 : _GEN_14142; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14144 = 7'h30 == out_payload_3_rob_idx[6:0] ? rob_egress_id_48 : _GEN_14143; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14145 = 7'h31 == out_payload_3_rob_idx[6:0] ? rob_egress_id_49 : _GEN_14144; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14146 = 7'h32 == out_payload_3_rob_idx[6:0] ? rob_egress_id_50 : _GEN_14145; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14147 = 7'h33 == out_payload_3_rob_idx[6:0] ? rob_egress_id_51 : _GEN_14146; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14148 = 7'h34 == out_payload_3_rob_idx[6:0] ? rob_egress_id_52 : _GEN_14147; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14149 = 7'h35 == out_payload_3_rob_idx[6:0] ? rob_egress_id_53 : _GEN_14148; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14150 = 7'h36 == out_payload_3_rob_idx[6:0] ? rob_egress_id_54 : _GEN_14149; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14151 = 7'h37 == out_payload_3_rob_idx[6:0] ? rob_egress_id_55 : _GEN_14150; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14152 = 7'h38 == out_payload_3_rob_idx[6:0] ? rob_egress_id_56 : _GEN_14151; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14153 = 7'h39 == out_payload_3_rob_idx[6:0] ? rob_egress_id_57 : _GEN_14152; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14154 = 7'h3a == out_payload_3_rob_idx[6:0] ? rob_egress_id_58 : _GEN_14153; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14155 = 7'h3b == out_payload_3_rob_idx[6:0] ? rob_egress_id_59 : _GEN_14154; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14156 = 7'h3c == out_payload_3_rob_idx[6:0] ? rob_egress_id_60 : _GEN_14155; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14157 = 7'h3d == out_payload_3_rob_idx[6:0] ? rob_egress_id_61 : _GEN_14156; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14158 = 7'h3e == out_payload_3_rob_idx[6:0] ? rob_egress_id_62 : _GEN_14157; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14159 = 7'h3f == out_payload_3_rob_idx[6:0] ? rob_egress_id_63 : _GEN_14158; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14160 = 7'h40 == out_payload_3_rob_idx[6:0] ? rob_egress_id_64 : _GEN_14159; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14161 = 7'h41 == out_payload_3_rob_idx[6:0] ? rob_egress_id_65 : _GEN_14160; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14162 = 7'h42 == out_payload_3_rob_idx[6:0] ? rob_egress_id_66 : _GEN_14161; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14163 = 7'h43 == out_payload_3_rob_idx[6:0] ? rob_egress_id_67 : _GEN_14162; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14164 = 7'h44 == out_payload_3_rob_idx[6:0] ? rob_egress_id_68 : _GEN_14163; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14165 = 7'h45 == out_payload_3_rob_idx[6:0] ? rob_egress_id_69 : _GEN_14164; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14166 = 7'h46 == out_payload_3_rob_idx[6:0] ? rob_egress_id_70 : _GEN_14165; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14167 = 7'h47 == out_payload_3_rob_idx[6:0] ? rob_egress_id_71 : _GEN_14166; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14168 = 7'h48 == out_payload_3_rob_idx[6:0] ? rob_egress_id_72 : _GEN_14167; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14169 = 7'h49 == out_payload_3_rob_idx[6:0] ? rob_egress_id_73 : _GEN_14168; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14170 = 7'h4a == out_payload_3_rob_idx[6:0] ? rob_egress_id_74 : _GEN_14169; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14171 = 7'h4b == out_payload_3_rob_idx[6:0] ? rob_egress_id_75 : _GEN_14170; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14172 = 7'h4c == out_payload_3_rob_idx[6:0] ? rob_egress_id_76 : _GEN_14171; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14173 = 7'h4d == out_payload_3_rob_idx[6:0] ? rob_egress_id_77 : _GEN_14172; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14174 = 7'h4e == out_payload_3_rob_idx[6:0] ? rob_egress_id_78 : _GEN_14173; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14175 = 7'h4f == out_payload_3_rob_idx[6:0] ? rob_egress_id_79 : _GEN_14174; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14176 = 7'h50 == out_payload_3_rob_idx[6:0] ? rob_egress_id_80 : _GEN_14175; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14177 = 7'h51 == out_payload_3_rob_idx[6:0] ? rob_egress_id_81 : _GEN_14176; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14178 = 7'h52 == out_payload_3_rob_idx[6:0] ? rob_egress_id_82 : _GEN_14177; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14179 = 7'h53 == out_payload_3_rob_idx[6:0] ? rob_egress_id_83 : _GEN_14178; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14180 = 7'h54 == out_payload_3_rob_idx[6:0] ? rob_egress_id_84 : _GEN_14179; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14181 = 7'h55 == out_payload_3_rob_idx[6:0] ? rob_egress_id_85 : _GEN_14180; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14182 = 7'h56 == out_payload_3_rob_idx[6:0] ? rob_egress_id_86 : _GEN_14181; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14183 = 7'h57 == out_payload_3_rob_idx[6:0] ? rob_egress_id_87 : _GEN_14182; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14184 = 7'h58 == out_payload_3_rob_idx[6:0] ? rob_egress_id_88 : _GEN_14183; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14185 = 7'h59 == out_payload_3_rob_idx[6:0] ? rob_egress_id_89 : _GEN_14184; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14186 = 7'h5a == out_payload_3_rob_idx[6:0] ? rob_egress_id_90 : _GEN_14185; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14187 = 7'h5b == out_payload_3_rob_idx[6:0] ? rob_egress_id_91 : _GEN_14186; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14188 = 7'h5c == out_payload_3_rob_idx[6:0] ? rob_egress_id_92 : _GEN_14187; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14189 = 7'h5d == out_payload_3_rob_idx[6:0] ? rob_egress_id_93 : _GEN_14188; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14190 = 7'h5e == out_payload_3_rob_idx[6:0] ? rob_egress_id_94 : _GEN_14189; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14191 = 7'h5f == out_payload_3_rob_idx[6:0] ? rob_egress_id_95 : _GEN_14190; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14192 = 7'h60 == out_payload_3_rob_idx[6:0] ? rob_egress_id_96 : _GEN_14191; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14193 = 7'h61 == out_payload_3_rob_idx[6:0] ? rob_egress_id_97 : _GEN_14192; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14194 = 7'h62 == out_payload_3_rob_idx[6:0] ? rob_egress_id_98 : _GEN_14193; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14195 = 7'h63 == out_payload_3_rob_idx[6:0] ? rob_egress_id_99 : _GEN_14194; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14196 = 7'h64 == out_payload_3_rob_idx[6:0] ? rob_egress_id_100 : _GEN_14195; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14197 = 7'h65 == out_payload_3_rob_idx[6:0] ? rob_egress_id_101 : _GEN_14196; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14198 = 7'h66 == out_payload_3_rob_idx[6:0] ? rob_egress_id_102 : _GEN_14197; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14199 = 7'h67 == out_payload_3_rob_idx[6:0] ? rob_egress_id_103 : _GEN_14198; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14200 = 7'h68 == out_payload_3_rob_idx[6:0] ? rob_egress_id_104 : _GEN_14199; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14201 = 7'h69 == out_payload_3_rob_idx[6:0] ? rob_egress_id_105 : _GEN_14200; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14202 = 7'h6a == out_payload_3_rob_idx[6:0] ? rob_egress_id_106 : _GEN_14201; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14203 = 7'h6b == out_payload_3_rob_idx[6:0] ? rob_egress_id_107 : _GEN_14202; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14204 = 7'h6c == out_payload_3_rob_idx[6:0] ? rob_egress_id_108 : _GEN_14203; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14205 = 7'h6d == out_payload_3_rob_idx[6:0] ? rob_egress_id_109 : _GEN_14204; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14206 = 7'h6e == out_payload_3_rob_idx[6:0] ? rob_egress_id_110 : _GEN_14205; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14207 = 7'h6f == out_payload_3_rob_idx[6:0] ? rob_egress_id_111 : _GEN_14206; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14208 = 7'h70 == out_payload_3_rob_idx[6:0] ? rob_egress_id_112 : _GEN_14207; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14209 = 7'h71 == out_payload_3_rob_idx[6:0] ? rob_egress_id_113 : _GEN_14208; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14210 = 7'h72 == out_payload_3_rob_idx[6:0] ? rob_egress_id_114 : _GEN_14209; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14211 = 7'h73 == out_payload_3_rob_idx[6:0] ? rob_egress_id_115 : _GEN_14210; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14212 = 7'h74 == out_payload_3_rob_idx[6:0] ? rob_egress_id_116 : _GEN_14211; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14213 = 7'h75 == out_payload_3_rob_idx[6:0] ? rob_egress_id_117 : _GEN_14212; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14214 = 7'h76 == out_payload_3_rob_idx[6:0] ? rob_egress_id_118 : _GEN_14213; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14215 = 7'h77 == out_payload_3_rob_idx[6:0] ? rob_egress_id_119 : _GEN_14214; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14216 = 7'h78 == out_payload_3_rob_idx[6:0] ? rob_egress_id_120 : _GEN_14215; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14217 = 7'h79 == out_payload_3_rob_idx[6:0] ? rob_egress_id_121 : _GEN_14216; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14218 = 7'h7a == out_payload_3_rob_idx[6:0] ? rob_egress_id_122 : _GEN_14217; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14219 = 7'h7b == out_payload_3_rob_idx[6:0] ? rob_egress_id_123 : _GEN_14218; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14220 = 7'h7c == out_payload_3_rob_idx[6:0] ? rob_egress_id_124 : _GEN_14219; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14221 = 7'h7d == out_payload_3_rob_idx[6:0] ? rob_egress_id_125 : _GEN_14220; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14222 = 7'h7e == out_payload_3_rob_idx[6:0] ? rob_egress_id_126 : _GEN_14221; // @[TestHarness.scala 204:{18,18}]
  wire [1:0] _GEN_14223 = 7'h7f == out_payload_3_rob_idx[6:0] ? rob_egress_id_127 : _GEN_14222; // @[TestHarness.scala 204:{18,18}]
  wire [3:0] _GEN_14225 = 7'h1 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_1 : rob_flits_returned_0; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14226 = 7'h2 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_2 : _GEN_14225; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14227 = 7'h3 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_3 : _GEN_14226; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14228 = 7'h4 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_4 : _GEN_14227; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14229 = 7'h5 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_5 : _GEN_14228; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14230 = 7'h6 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_6 : _GEN_14229; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14231 = 7'h7 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_7 : _GEN_14230; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14232 = 7'h8 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_8 : _GEN_14231; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14233 = 7'h9 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_9 : _GEN_14232; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14234 = 7'ha == out_payload_3_rob_idx[6:0] ? rob_flits_returned_10 : _GEN_14233; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14235 = 7'hb == out_payload_3_rob_idx[6:0] ? rob_flits_returned_11 : _GEN_14234; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14236 = 7'hc == out_payload_3_rob_idx[6:0] ? rob_flits_returned_12 : _GEN_14235; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14237 = 7'hd == out_payload_3_rob_idx[6:0] ? rob_flits_returned_13 : _GEN_14236; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14238 = 7'he == out_payload_3_rob_idx[6:0] ? rob_flits_returned_14 : _GEN_14237; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14239 = 7'hf == out_payload_3_rob_idx[6:0] ? rob_flits_returned_15 : _GEN_14238; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14240 = 7'h10 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_16 : _GEN_14239; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14241 = 7'h11 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_17 : _GEN_14240; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14242 = 7'h12 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_18 : _GEN_14241; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14243 = 7'h13 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_19 : _GEN_14242; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14244 = 7'h14 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_20 : _GEN_14243; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14245 = 7'h15 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_21 : _GEN_14244; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14246 = 7'h16 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_22 : _GEN_14245; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14247 = 7'h17 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_23 : _GEN_14246; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14248 = 7'h18 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_24 : _GEN_14247; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14249 = 7'h19 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_25 : _GEN_14248; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14250 = 7'h1a == out_payload_3_rob_idx[6:0] ? rob_flits_returned_26 : _GEN_14249; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14251 = 7'h1b == out_payload_3_rob_idx[6:0] ? rob_flits_returned_27 : _GEN_14250; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14252 = 7'h1c == out_payload_3_rob_idx[6:0] ? rob_flits_returned_28 : _GEN_14251; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14253 = 7'h1d == out_payload_3_rob_idx[6:0] ? rob_flits_returned_29 : _GEN_14252; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14254 = 7'h1e == out_payload_3_rob_idx[6:0] ? rob_flits_returned_30 : _GEN_14253; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14255 = 7'h1f == out_payload_3_rob_idx[6:0] ? rob_flits_returned_31 : _GEN_14254; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14256 = 7'h20 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_32 : _GEN_14255; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14257 = 7'h21 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_33 : _GEN_14256; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14258 = 7'h22 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_34 : _GEN_14257; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14259 = 7'h23 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_35 : _GEN_14258; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14260 = 7'h24 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_36 : _GEN_14259; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14261 = 7'h25 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_37 : _GEN_14260; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14262 = 7'h26 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_38 : _GEN_14261; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14263 = 7'h27 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_39 : _GEN_14262; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14264 = 7'h28 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_40 : _GEN_14263; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14265 = 7'h29 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_41 : _GEN_14264; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14266 = 7'h2a == out_payload_3_rob_idx[6:0] ? rob_flits_returned_42 : _GEN_14265; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14267 = 7'h2b == out_payload_3_rob_idx[6:0] ? rob_flits_returned_43 : _GEN_14266; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14268 = 7'h2c == out_payload_3_rob_idx[6:0] ? rob_flits_returned_44 : _GEN_14267; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14269 = 7'h2d == out_payload_3_rob_idx[6:0] ? rob_flits_returned_45 : _GEN_14268; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14270 = 7'h2e == out_payload_3_rob_idx[6:0] ? rob_flits_returned_46 : _GEN_14269; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14271 = 7'h2f == out_payload_3_rob_idx[6:0] ? rob_flits_returned_47 : _GEN_14270; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14272 = 7'h30 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_48 : _GEN_14271; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14273 = 7'h31 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_49 : _GEN_14272; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14274 = 7'h32 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_50 : _GEN_14273; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14275 = 7'h33 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_51 : _GEN_14274; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14276 = 7'h34 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_52 : _GEN_14275; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14277 = 7'h35 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_53 : _GEN_14276; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14278 = 7'h36 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_54 : _GEN_14277; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14279 = 7'h37 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_55 : _GEN_14278; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14280 = 7'h38 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_56 : _GEN_14279; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14281 = 7'h39 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_57 : _GEN_14280; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14282 = 7'h3a == out_payload_3_rob_idx[6:0] ? rob_flits_returned_58 : _GEN_14281; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14283 = 7'h3b == out_payload_3_rob_idx[6:0] ? rob_flits_returned_59 : _GEN_14282; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14284 = 7'h3c == out_payload_3_rob_idx[6:0] ? rob_flits_returned_60 : _GEN_14283; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14285 = 7'h3d == out_payload_3_rob_idx[6:0] ? rob_flits_returned_61 : _GEN_14284; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14286 = 7'h3e == out_payload_3_rob_idx[6:0] ? rob_flits_returned_62 : _GEN_14285; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14287 = 7'h3f == out_payload_3_rob_idx[6:0] ? rob_flits_returned_63 : _GEN_14286; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14288 = 7'h40 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_64 : _GEN_14287; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14289 = 7'h41 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_65 : _GEN_14288; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14290 = 7'h42 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_66 : _GEN_14289; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14291 = 7'h43 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_67 : _GEN_14290; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14292 = 7'h44 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_68 : _GEN_14291; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14293 = 7'h45 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_69 : _GEN_14292; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14294 = 7'h46 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_70 : _GEN_14293; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14295 = 7'h47 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_71 : _GEN_14294; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14296 = 7'h48 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_72 : _GEN_14295; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14297 = 7'h49 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_73 : _GEN_14296; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14298 = 7'h4a == out_payload_3_rob_idx[6:0] ? rob_flits_returned_74 : _GEN_14297; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14299 = 7'h4b == out_payload_3_rob_idx[6:0] ? rob_flits_returned_75 : _GEN_14298; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14300 = 7'h4c == out_payload_3_rob_idx[6:0] ? rob_flits_returned_76 : _GEN_14299; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14301 = 7'h4d == out_payload_3_rob_idx[6:0] ? rob_flits_returned_77 : _GEN_14300; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14302 = 7'h4e == out_payload_3_rob_idx[6:0] ? rob_flits_returned_78 : _GEN_14301; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14303 = 7'h4f == out_payload_3_rob_idx[6:0] ? rob_flits_returned_79 : _GEN_14302; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14304 = 7'h50 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_80 : _GEN_14303; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14305 = 7'h51 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_81 : _GEN_14304; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14306 = 7'h52 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_82 : _GEN_14305; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14307 = 7'h53 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_83 : _GEN_14306; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14308 = 7'h54 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_84 : _GEN_14307; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14309 = 7'h55 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_85 : _GEN_14308; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14310 = 7'h56 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_86 : _GEN_14309; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14311 = 7'h57 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_87 : _GEN_14310; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14312 = 7'h58 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_88 : _GEN_14311; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14313 = 7'h59 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_89 : _GEN_14312; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14314 = 7'h5a == out_payload_3_rob_idx[6:0] ? rob_flits_returned_90 : _GEN_14313; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14315 = 7'h5b == out_payload_3_rob_idx[6:0] ? rob_flits_returned_91 : _GEN_14314; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14316 = 7'h5c == out_payload_3_rob_idx[6:0] ? rob_flits_returned_92 : _GEN_14315; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14317 = 7'h5d == out_payload_3_rob_idx[6:0] ? rob_flits_returned_93 : _GEN_14316; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14318 = 7'h5e == out_payload_3_rob_idx[6:0] ? rob_flits_returned_94 : _GEN_14317; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14319 = 7'h5f == out_payload_3_rob_idx[6:0] ? rob_flits_returned_95 : _GEN_14318; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14320 = 7'h60 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_96 : _GEN_14319; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14321 = 7'h61 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_97 : _GEN_14320; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14322 = 7'h62 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_98 : _GEN_14321; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14323 = 7'h63 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_99 : _GEN_14322; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14324 = 7'h64 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_100 : _GEN_14323; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14325 = 7'h65 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_101 : _GEN_14324; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14326 = 7'h66 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_102 : _GEN_14325; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14327 = 7'h67 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_103 : _GEN_14326; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14328 = 7'h68 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_104 : _GEN_14327; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14329 = 7'h69 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_105 : _GEN_14328; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14330 = 7'h6a == out_payload_3_rob_idx[6:0] ? rob_flits_returned_106 : _GEN_14329; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14331 = 7'h6b == out_payload_3_rob_idx[6:0] ? rob_flits_returned_107 : _GEN_14330; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14332 = 7'h6c == out_payload_3_rob_idx[6:0] ? rob_flits_returned_108 : _GEN_14331; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14333 = 7'h6d == out_payload_3_rob_idx[6:0] ? rob_flits_returned_109 : _GEN_14332; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14334 = 7'h6e == out_payload_3_rob_idx[6:0] ? rob_flits_returned_110 : _GEN_14333; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14335 = 7'h6f == out_payload_3_rob_idx[6:0] ? rob_flits_returned_111 : _GEN_14334; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14336 = 7'h70 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_112 : _GEN_14335; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14337 = 7'h71 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_113 : _GEN_14336; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14338 = 7'h72 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_114 : _GEN_14337; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14339 = 7'h73 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_115 : _GEN_14338; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14340 = 7'h74 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_116 : _GEN_14339; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14341 = 7'h75 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_117 : _GEN_14340; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14342 = 7'h76 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_118 : _GEN_14341; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14343 = 7'h77 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_119 : _GEN_14342; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14344 = 7'h78 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_120 : _GEN_14343; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14345 = 7'h79 == out_payload_3_rob_idx[6:0] ? rob_flits_returned_121 : _GEN_14344; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14346 = 7'h7a == out_payload_3_rob_idx[6:0] ? rob_flits_returned_122 : _GEN_14345; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14347 = 7'h7b == out_payload_3_rob_idx[6:0] ? rob_flits_returned_123 : _GEN_14346; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14348 = 7'h7c == out_payload_3_rob_idx[6:0] ? rob_flits_returned_124 : _GEN_14347; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14349 = 7'h7d == out_payload_3_rob_idx[6:0] ? rob_flits_returned_125 : _GEN_14348; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14350 = 7'h7e == out_payload_3_rob_idx[6:0] ? rob_flits_returned_126 : _GEN_14349; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14351 = 7'h7f == out_payload_3_rob_idx[6:0] ? rob_flits_returned_127 : _GEN_14350; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14353 = 7'h1 == out_payload_3_rob_idx[6:0] ? rob_n_flits_1 : rob_n_flits_0; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14354 = 7'h2 == out_payload_3_rob_idx[6:0] ? rob_n_flits_2 : _GEN_14353; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14355 = 7'h3 == out_payload_3_rob_idx[6:0] ? rob_n_flits_3 : _GEN_14354; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14356 = 7'h4 == out_payload_3_rob_idx[6:0] ? rob_n_flits_4 : _GEN_14355; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14357 = 7'h5 == out_payload_3_rob_idx[6:0] ? rob_n_flits_5 : _GEN_14356; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14358 = 7'h6 == out_payload_3_rob_idx[6:0] ? rob_n_flits_6 : _GEN_14357; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14359 = 7'h7 == out_payload_3_rob_idx[6:0] ? rob_n_flits_7 : _GEN_14358; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14360 = 7'h8 == out_payload_3_rob_idx[6:0] ? rob_n_flits_8 : _GEN_14359; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14361 = 7'h9 == out_payload_3_rob_idx[6:0] ? rob_n_flits_9 : _GEN_14360; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14362 = 7'ha == out_payload_3_rob_idx[6:0] ? rob_n_flits_10 : _GEN_14361; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14363 = 7'hb == out_payload_3_rob_idx[6:0] ? rob_n_flits_11 : _GEN_14362; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14364 = 7'hc == out_payload_3_rob_idx[6:0] ? rob_n_flits_12 : _GEN_14363; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14365 = 7'hd == out_payload_3_rob_idx[6:0] ? rob_n_flits_13 : _GEN_14364; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14366 = 7'he == out_payload_3_rob_idx[6:0] ? rob_n_flits_14 : _GEN_14365; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14367 = 7'hf == out_payload_3_rob_idx[6:0] ? rob_n_flits_15 : _GEN_14366; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14368 = 7'h10 == out_payload_3_rob_idx[6:0] ? rob_n_flits_16 : _GEN_14367; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14369 = 7'h11 == out_payload_3_rob_idx[6:0] ? rob_n_flits_17 : _GEN_14368; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14370 = 7'h12 == out_payload_3_rob_idx[6:0] ? rob_n_flits_18 : _GEN_14369; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14371 = 7'h13 == out_payload_3_rob_idx[6:0] ? rob_n_flits_19 : _GEN_14370; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14372 = 7'h14 == out_payload_3_rob_idx[6:0] ? rob_n_flits_20 : _GEN_14371; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14373 = 7'h15 == out_payload_3_rob_idx[6:0] ? rob_n_flits_21 : _GEN_14372; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14374 = 7'h16 == out_payload_3_rob_idx[6:0] ? rob_n_flits_22 : _GEN_14373; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14375 = 7'h17 == out_payload_3_rob_idx[6:0] ? rob_n_flits_23 : _GEN_14374; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14376 = 7'h18 == out_payload_3_rob_idx[6:0] ? rob_n_flits_24 : _GEN_14375; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14377 = 7'h19 == out_payload_3_rob_idx[6:0] ? rob_n_flits_25 : _GEN_14376; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14378 = 7'h1a == out_payload_3_rob_idx[6:0] ? rob_n_flits_26 : _GEN_14377; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14379 = 7'h1b == out_payload_3_rob_idx[6:0] ? rob_n_flits_27 : _GEN_14378; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14380 = 7'h1c == out_payload_3_rob_idx[6:0] ? rob_n_flits_28 : _GEN_14379; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14381 = 7'h1d == out_payload_3_rob_idx[6:0] ? rob_n_flits_29 : _GEN_14380; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14382 = 7'h1e == out_payload_3_rob_idx[6:0] ? rob_n_flits_30 : _GEN_14381; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14383 = 7'h1f == out_payload_3_rob_idx[6:0] ? rob_n_flits_31 : _GEN_14382; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14384 = 7'h20 == out_payload_3_rob_idx[6:0] ? rob_n_flits_32 : _GEN_14383; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14385 = 7'h21 == out_payload_3_rob_idx[6:0] ? rob_n_flits_33 : _GEN_14384; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14386 = 7'h22 == out_payload_3_rob_idx[6:0] ? rob_n_flits_34 : _GEN_14385; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14387 = 7'h23 == out_payload_3_rob_idx[6:0] ? rob_n_flits_35 : _GEN_14386; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14388 = 7'h24 == out_payload_3_rob_idx[6:0] ? rob_n_flits_36 : _GEN_14387; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14389 = 7'h25 == out_payload_3_rob_idx[6:0] ? rob_n_flits_37 : _GEN_14388; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14390 = 7'h26 == out_payload_3_rob_idx[6:0] ? rob_n_flits_38 : _GEN_14389; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14391 = 7'h27 == out_payload_3_rob_idx[6:0] ? rob_n_flits_39 : _GEN_14390; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14392 = 7'h28 == out_payload_3_rob_idx[6:0] ? rob_n_flits_40 : _GEN_14391; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14393 = 7'h29 == out_payload_3_rob_idx[6:0] ? rob_n_flits_41 : _GEN_14392; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14394 = 7'h2a == out_payload_3_rob_idx[6:0] ? rob_n_flits_42 : _GEN_14393; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14395 = 7'h2b == out_payload_3_rob_idx[6:0] ? rob_n_flits_43 : _GEN_14394; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14396 = 7'h2c == out_payload_3_rob_idx[6:0] ? rob_n_flits_44 : _GEN_14395; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14397 = 7'h2d == out_payload_3_rob_idx[6:0] ? rob_n_flits_45 : _GEN_14396; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14398 = 7'h2e == out_payload_3_rob_idx[6:0] ? rob_n_flits_46 : _GEN_14397; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14399 = 7'h2f == out_payload_3_rob_idx[6:0] ? rob_n_flits_47 : _GEN_14398; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14400 = 7'h30 == out_payload_3_rob_idx[6:0] ? rob_n_flits_48 : _GEN_14399; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14401 = 7'h31 == out_payload_3_rob_idx[6:0] ? rob_n_flits_49 : _GEN_14400; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14402 = 7'h32 == out_payload_3_rob_idx[6:0] ? rob_n_flits_50 : _GEN_14401; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14403 = 7'h33 == out_payload_3_rob_idx[6:0] ? rob_n_flits_51 : _GEN_14402; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14404 = 7'h34 == out_payload_3_rob_idx[6:0] ? rob_n_flits_52 : _GEN_14403; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14405 = 7'h35 == out_payload_3_rob_idx[6:0] ? rob_n_flits_53 : _GEN_14404; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14406 = 7'h36 == out_payload_3_rob_idx[6:0] ? rob_n_flits_54 : _GEN_14405; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14407 = 7'h37 == out_payload_3_rob_idx[6:0] ? rob_n_flits_55 : _GEN_14406; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14408 = 7'h38 == out_payload_3_rob_idx[6:0] ? rob_n_flits_56 : _GEN_14407; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14409 = 7'h39 == out_payload_3_rob_idx[6:0] ? rob_n_flits_57 : _GEN_14408; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14410 = 7'h3a == out_payload_3_rob_idx[6:0] ? rob_n_flits_58 : _GEN_14409; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14411 = 7'h3b == out_payload_3_rob_idx[6:0] ? rob_n_flits_59 : _GEN_14410; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14412 = 7'h3c == out_payload_3_rob_idx[6:0] ? rob_n_flits_60 : _GEN_14411; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14413 = 7'h3d == out_payload_3_rob_idx[6:0] ? rob_n_flits_61 : _GEN_14412; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14414 = 7'h3e == out_payload_3_rob_idx[6:0] ? rob_n_flits_62 : _GEN_14413; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14415 = 7'h3f == out_payload_3_rob_idx[6:0] ? rob_n_flits_63 : _GEN_14414; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14416 = 7'h40 == out_payload_3_rob_idx[6:0] ? rob_n_flits_64 : _GEN_14415; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14417 = 7'h41 == out_payload_3_rob_idx[6:0] ? rob_n_flits_65 : _GEN_14416; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14418 = 7'h42 == out_payload_3_rob_idx[6:0] ? rob_n_flits_66 : _GEN_14417; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14419 = 7'h43 == out_payload_3_rob_idx[6:0] ? rob_n_flits_67 : _GEN_14418; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14420 = 7'h44 == out_payload_3_rob_idx[6:0] ? rob_n_flits_68 : _GEN_14419; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14421 = 7'h45 == out_payload_3_rob_idx[6:0] ? rob_n_flits_69 : _GEN_14420; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14422 = 7'h46 == out_payload_3_rob_idx[6:0] ? rob_n_flits_70 : _GEN_14421; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14423 = 7'h47 == out_payload_3_rob_idx[6:0] ? rob_n_flits_71 : _GEN_14422; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14424 = 7'h48 == out_payload_3_rob_idx[6:0] ? rob_n_flits_72 : _GEN_14423; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14425 = 7'h49 == out_payload_3_rob_idx[6:0] ? rob_n_flits_73 : _GEN_14424; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14426 = 7'h4a == out_payload_3_rob_idx[6:0] ? rob_n_flits_74 : _GEN_14425; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14427 = 7'h4b == out_payload_3_rob_idx[6:0] ? rob_n_flits_75 : _GEN_14426; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14428 = 7'h4c == out_payload_3_rob_idx[6:0] ? rob_n_flits_76 : _GEN_14427; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14429 = 7'h4d == out_payload_3_rob_idx[6:0] ? rob_n_flits_77 : _GEN_14428; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14430 = 7'h4e == out_payload_3_rob_idx[6:0] ? rob_n_flits_78 : _GEN_14429; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14431 = 7'h4f == out_payload_3_rob_idx[6:0] ? rob_n_flits_79 : _GEN_14430; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14432 = 7'h50 == out_payload_3_rob_idx[6:0] ? rob_n_flits_80 : _GEN_14431; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14433 = 7'h51 == out_payload_3_rob_idx[6:0] ? rob_n_flits_81 : _GEN_14432; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14434 = 7'h52 == out_payload_3_rob_idx[6:0] ? rob_n_flits_82 : _GEN_14433; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14435 = 7'h53 == out_payload_3_rob_idx[6:0] ? rob_n_flits_83 : _GEN_14434; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14436 = 7'h54 == out_payload_3_rob_idx[6:0] ? rob_n_flits_84 : _GEN_14435; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14437 = 7'h55 == out_payload_3_rob_idx[6:0] ? rob_n_flits_85 : _GEN_14436; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14438 = 7'h56 == out_payload_3_rob_idx[6:0] ? rob_n_flits_86 : _GEN_14437; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14439 = 7'h57 == out_payload_3_rob_idx[6:0] ? rob_n_flits_87 : _GEN_14438; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14440 = 7'h58 == out_payload_3_rob_idx[6:0] ? rob_n_flits_88 : _GEN_14439; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14441 = 7'h59 == out_payload_3_rob_idx[6:0] ? rob_n_flits_89 : _GEN_14440; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14442 = 7'h5a == out_payload_3_rob_idx[6:0] ? rob_n_flits_90 : _GEN_14441; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14443 = 7'h5b == out_payload_3_rob_idx[6:0] ? rob_n_flits_91 : _GEN_14442; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14444 = 7'h5c == out_payload_3_rob_idx[6:0] ? rob_n_flits_92 : _GEN_14443; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14445 = 7'h5d == out_payload_3_rob_idx[6:0] ? rob_n_flits_93 : _GEN_14444; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14446 = 7'h5e == out_payload_3_rob_idx[6:0] ? rob_n_flits_94 : _GEN_14445; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14447 = 7'h5f == out_payload_3_rob_idx[6:0] ? rob_n_flits_95 : _GEN_14446; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14448 = 7'h60 == out_payload_3_rob_idx[6:0] ? rob_n_flits_96 : _GEN_14447; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14449 = 7'h61 == out_payload_3_rob_idx[6:0] ? rob_n_flits_97 : _GEN_14448; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14450 = 7'h62 == out_payload_3_rob_idx[6:0] ? rob_n_flits_98 : _GEN_14449; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14451 = 7'h63 == out_payload_3_rob_idx[6:0] ? rob_n_flits_99 : _GEN_14450; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14452 = 7'h64 == out_payload_3_rob_idx[6:0] ? rob_n_flits_100 : _GEN_14451; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14453 = 7'h65 == out_payload_3_rob_idx[6:0] ? rob_n_flits_101 : _GEN_14452; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14454 = 7'h66 == out_payload_3_rob_idx[6:0] ? rob_n_flits_102 : _GEN_14453; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14455 = 7'h67 == out_payload_3_rob_idx[6:0] ? rob_n_flits_103 : _GEN_14454; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14456 = 7'h68 == out_payload_3_rob_idx[6:0] ? rob_n_flits_104 : _GEN_14455; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14457 = 7'h69 == out_payload_3_rob_idx[6:0] ? rob_n_flits_105 : _GEN_14456; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14458 = 7'h6a == out_payload_3_rob_idx[6:0] ? rob_n_flits_106 : _GEN_14457; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14459 = 7'h6b == out_payload_3_rob_idx[6:0] ? rob_n_flits_107 : _GEN_14458; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14460 = 7'h6c == out_payload_3_rob_idx[6:0] ? rob_n_flits_108 : _GEN_14459; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14461 = 7'h6d == out_payload_3_rob_idx[6:0] ? rob_n_flits_109 : _GEN_14460; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14462 = 7'h6e == out_payload_3_rob_idx[6:0] ? rob_n_flits_110 : _GEN_14461; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14463 = 7'h6f == out_payload_3_rob_idx[6:0] ? rob_n_flits_111 : _GEN_14462; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14464 = 7'h70 == out_payload_3_rob_idx[6:0] ? rob_n_flits_112 : _GEN_14463; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14465 = 7'h71 == out_payload_3_rob_idx[6:0] ? rob_n_flits_113 : _GEN_14464; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14466 = 7'h72 == out_payload_3_rob_idx[6:0] ? rob_n_flits_114 : _GEN_14465; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14467 = 7'h73 == out_payload_3_rob_idx[6:0] ? rob_n_flits_115 : _GEN_14466; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14468 = 7'h74 == out_payload_3_rob_idx[6:0] ? rob_n_flits_116 : _GEN_14467; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14469 = 7'h75 == out_payload_3_rob_idx[6:0] ? rob_n_flits_117 : _GEN_14468; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14470 = 7'h76 == out_payload_3_rob_idx[6:0] ? rob_n_flits_118 : _GEN_14469; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14471 = 7'h77 == out_payload_3_rob_idx[6:0] ? rob_n_flits_119 : _GEN_14470; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14472 = 7'h78 == out_payload_3_rob_idx[6:0] ? rob_n_flits_120 : _GEN_14471; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14473 = 7'h79 == out_payload_3_rob_idx[6:0] ? rob_n_flits_121 : _GEN_14472; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14474 = 7'h7a == out_payload_3_rob_idx[6:0] ? rob_n_flits_122 : _GEN_14473; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14475 = 7'h7b == out_payload_3_rob_idx[6:0] ? rob_n_flits_123 : _GEN_14474; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14476 = 7'h7c == out_payload_3_rob_idx[6:0] ? rob_n_flits_124 : _GEN_14475; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14477 = 7'h7d == out_payload_3_rob_idx[6:0] ? rob_n_flits_125 : _GEN_14476; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14478 = 7'h7e == out_payload_3_rob_idx[6:0] ? rob_n_flits_126 : _GEN_14477; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_14479 = 7'h7f == out_payload_3_rob_idx[6:0] ? rob_n_flits_127 : _GEN_14478; // @[TestHarness.scala 205:{42,42}]
  wire [15:0] _GEN_15384 = {{9'd0}, packet_rob_idx_3}; // @[TestHarness.scala 206:61]
  wire  _T_251 = io_from_noc_3_flit_bits_head & enable_print_latency; // @[TestHarness.scala 208:30]
  wire [3:0] _rob_flits_returned_T_11 = _GEN_14351 + 4'h1; // @[TestHarness.scala 213:66]
  wire [15:0] _rob_payload_flits_fired_T_11 = _GEN_13967 + 16'h1; // @[TestHarness.scala 214:76]
  wire  _GEN_15120 = io_from_noc_3_flit_bits_head | packet_valid_3; // @[TestHarness.scala 196:31 215:{31,46}]
  wire [15:0] _GEN_15121 = io_from_noc_3_flit_bits_head ? out_payload_3_rob_idx : {{9'd0}, packet_rob_idx_3}; // @[TestHarness.scala 197:29 215:{31,72}]
  wire [15:0] _GEN_15380 = _T_259 ? _GEN_15121 : {{9'd0}, packet_rob_idx_3}; // @[TestHarness.scala 199:26 197:29]
  wire [127:0] _rob_valids_T = rob_valids | rob_allocs; // @[TestHarness.scala 222:29]
  wire [65535:0] _rob_valids_T_1 = ~rob_frees; // @[TestHarness.scala 222:45]
  wire [65535:0] _GEN_15385 = {{65408'd0}, _rob_valids_T}; // @[TestHarness.scala 222:43]
  wire [65535:0] _rob_valids_T_2 = _GEN_15385 & _rob_valids_T_1; // @[TestHarness.scala 222:43]
  wire [1:0] _flits_T_4 = _T_118 + _T_165; // @[TestHarness.scala 224:66]
  wire [1:0] _GEN_15386 = {{1'd0}, _T_212}; // @[TestHarness.scala 224:66]
  wire [2:0] _flits_T_5 = _flits_T_4 + _GEN_15386; // @[TestHarness.scala 224:66]
  wire [2:0] _GEN_15387 = {{2'd0}, _T_259}; // @[TestHarness.scala 224:66]
  wire [3:0] _flits_T_6 = _flits_T_5 + _GEN_15387; // @[TestHarness.scala 224:66]
  wire [31:0] _GEN_15388 = {{28'd0}, _flits_T_6}; // @[TestHarness.scala 224:18]
  wire [31:0] _flits_T_8 = flits + _GEN_15388; // @[TestHarness.scala 224:18]
  wire  tx_fire_0 = igen_io_fire; // @[TestHarness.scala 169:21 186:18]
  wire  tx_fire_1 = igen_1_io_fire; // @[TestHarness.scala 169:21 186:18]
  wire [1:0] _txs_T = tx_fire_0 + tx_fire_1; // @[Bitwise.scala 51:90]
  wire  tx_fire_2 = igen_2_io_fire; // @[TestHarness.scala 169:21 186:18]
  wire  tx_fire_3 = igen_3_io_fire; // @[TestHarness.scala 169:21 186:18]
  wire [1:0] _txs_T_2 = tx_fire_2 + tx_fire_3; // @[Bitwise.scala 51:90]
  wire [2:0] _txs_T_4 = _txs_T + _txs_T_2; // @[Bitwise.scala 51:90]
  wire [31:0] _GEN_15389 = {{29'd0}, _txs_T_4}; // @[TestHarness.scala 225:14]
  wire [31:0] _txs_T_7 = txs + _GEN_15389; // @[TestHarness.scala 225:14]
  wire [63:0] _T_264 = _rob_tscs_T_31 - rob_tscs_0; // @[TestHarness.scala 229:18]
  wire [63:0] _T_271 = _rob_tscs_T_31 - rob_tscs_1; // @[TestHarness.scala 229:18]
  wire [63:0] _T_278 = _rob_tscs_T_31 - rob_tscs_2; // @[TestHarness.scala 229:18]
  wire [63:0] _T_285 = _rob_tscs_T_31 - rob_tscs_3; // @[TestHarness.scala 229:18]
  wire [63:0] _T_292 = _rob_tscs_T_31 - rob_tscs_4; // @[TestHarness.scala 229:18]
  wire [63:0] _T_299 = _rob_tscs_T_31 - rob_tscs_5; // @[TestHarness.scala 229:18]
  wire [63:0] _T_306 = _rob_tscs_T_31 - rob_tscs_6; // @[TestHarness.scala 229:18]
  wire [63:0] _T_313 = _rob_tscs_T_31 - rob_tscs_7; // @[TestHarness.scala 229:18]
  wire [63:0] _T_320 = _rob_tscs_T_31 - rob_tscs_8; // @[TestHarness.scala 229:18]
  wire [63:0] _T_327 = _rob_tscs_T_31 - rob_tscs_9; // @[TestHarness.scala 229:18]
  wire [63:0] _T_334 = _rob_tscs_T_31 - rob_tscs_10; // @[TestHarness.scala 229:18]
  wire [63:0] _T_341 = _rob_tscs_T_31 - rob_tscs_11; // @[TestHarness.scala 229:18]
  wire [63:0] _T_348 = _rob_tscs_T_31 - rob_tscs_12; // @[TestHarness.scala 229:18]
  wire [63:0] _T_355 = _rob_tscs_T_31 - rob_tscs_13; // @[TestHarness.scala 229:18]
  wire [63:0] _T_362 = _rob_tscs_T_31 - rob_tscs_14; // @[TestHarness.scala 229:18]
  wire [63:0] _T_369 = _rob_tscs_T_31 - rob_tscs_15; // @[TestHarness.scala 229:18]
  wire [63:0] _T_376 = _rob_tscs_T_31 - rob_tscs_16; // @[TestHarness.scala 229:18]
  wire [63:0] _T_383 = _rob_tscs_T_31 - rob_tscs_17; // @[TestHarness.scala 229:18]
  wire [63:0] _T_390 = _rob_tscs_T_31 - rob_tscs_18; // @[TestHarness.scala 229:18]
  wire [63:0] _T_397 = _rob_tscs_T_31 - rob_tscs_19; // @[TestHarness.scala 229:18]
  wire [63:0] _T_404 = _rob_tscs_T_31 - rob_tscs_20; // @[TestHarness.scala 229:18]
  wire [63:0] _T_411 = _rob_tscs_T_31 - rob_tscs_21; // @[TestHarness.scala 229:18]
  wire [63:0] _T_418 = _rob_tscs_T_31 - rob_tscs_22; // @[TestHarness.scala 229:18]
  wire [63:0] _T_425 = _rob_tscs_T_31 - rob_tscs_23; // @[TestHarness.scala 229:18]
  wire [63:0] _T_432 = _rob_tscs_T_31 - rob_tscs_24; // @[TestHarness.scala 229:18]
  wire [63:0] _T_439 = _rob_tscs_T_31 - rob_tscs_25; // @[TestHarness.scala 229:18]
  wire [63:0] _T_446 = _rob_tscs_T_31 - rob_tscs_26; // @[TestHarness.scala 229:18]
  wire [63:0] _T_453 = _rob_tscs_T_31 - rob_tscs_27; // @[TestHarness.scala 229:18]
  wire [63:0] _T_460 = _rob_tscs_T_31 - rob_tscs_28; // @[TestHarness.scala 229:18]
  wire [63:0] _T_467 = _rob_tscs_T_31 - rob_tscs_29; // @[TestHarness.scala 229:18]
  wire [63:0] _T_474 = _rob_tscs_T_31 - rob_tscs_30; // @[TestHarness.scala 229:18]
  wire [63:0] _T_481 = _rob_tscs_T_31 - rob_tscs_31; // @[TestHarness.scala 229:18]
  wire [63:0] _T_488 = _rob_tscs_T_31 - rob_tscs_32; // @[TestHarness.scala 229:18]
  wire [63:0] _T_495 = _rob_tscs_T_31 - rob_tscs_33; // @[TestHarness.scala 229:18]
  wire [63:0] _T_502 = _rob_tscs_T_31 - rob_tscs_34; // @[TestHarness.scala 229:18]
  wire [63:0] _T_509 = _rob_tscs_T_31 - rob_tscs_35; // @[TestHarness.scala 229:18]
  wire [63:0] _T_516 = _rob_tscs_T_31 - rob_tscs_36; // @[TestHarness.scala 229:18]
  wire [63:0] _T_523 = _rob_tscs_T_31 - rob_tscs_37; // @[TestHarness.scala 229:18]
  wire [63:0] _T_530 = _rob_tscs_T_31 - rob_tscs_38; // @[TestHarness.scala 229:18]
  wire [63:0] _T_537 = _rob_tscs_T_31 - rob_tscs_39; // @[TestHarness.scala 229:18]
  wire [63:0] _T_544 = _rob_tscs_T_31 - rob_tscs_40; // @[TestHarness.scala 229:18]
  wire [63:0] _T_551 = _rob_tscs_T_31 - rob_tscs_41; // @[TestHarness.scala 229:18]
  wire [63:0] _T_558 = _rob_tscs_T_31 - rob_tscs_42; // @[TestHarness.scala 229:18]
  wire [63:0] _T_565 = _rob_tscs_T_31 - rob_tscs_43; // @[TestHarness.scala 229:18]
  wire [63:0] _T_572 = _rob_tscs_T_31 - rob_tscs_44; // @[TestHarness.scala 229:18]
  wire [63:0] _T_579 = _rob_tscs_T_31 - rob_tscs_45; // @[TestHarness.scala 229:18]
  wire [63:0] _T_586 = _rob_tscs_T_31 - rob_tscs_46; // @[TestHarness.scala 229:18]
  wire [63:0] _T_593 = _rob_tscs_T_31 - rob_tscs_47; // @[TestHarness.scala 229:18]
  wire [63:0] _T_600 = _rob_tscs_T_31 - rob_tscs_48; // @[TestHarness.scala 229:18]
  wire [63:0] _T_607 = _rob_tscs_T_31 - rob_tscs_49; // @[TestHarness.scala 229:18]
  wire [63:0] _T_614 = _rob_tscs_T_31 - rob_tscs_50; // @[TestHarness.scala 229:18]
  wire [63:0] _T_621 = _rob_tscs_T_31 - rob_tscs_51; // @[TestHarness.scala 229:18]
  wire [63:0] _T_628 = _rob_tscs_T_31 - rob_tscs_52; // @[TestHarness.scala 229:18]
  wire [63:0] _T_635 = _rob_tscs_T_31 - rob_tscs_53; // @[TestHarness.scala 229:18]
  wire [63:0] _T_642 = _rob_tscs_T_31 - rob_tscs_54; // @[TestHarness.scala 229:18]
  wire [63:0] _T_649 = _rob_tscs_T_31 - rob_tscs_55; // @[TestHarness.scala 229:18]
  wire [63:0] _T_656 = _rob_tscs_T_31 - rob_tscs_56; // @[TestHarness.scala 229:18]
  wire [63:0] _T_663 = _rob_tscs_T_31 - rob_tscs_57; // @[TestHarness.scala 229:18]
  wire [63:0] _T_670 = _rob_tscs_T_31 - rob_tscs_58; // @[TestHarness.scala 229:18]
  wire [63:0] _T_677 = _rob_tscs_T_31 - rob_tscs_59; // @[TestHarness.scala 229:18]
  wire [63:0] _T_684 = _rob_tscs_T_31 - rob_tscs_60; // @[TestHarness.scala 229:18]
  wire [63:0] _T_691 = _rob_tscs_T_31 - rob_tscs_61; // @[TestHarness.scala 229:18]
  wire [63:0] _T_698 = _rob_tscs_T_31 - rob_tscs_62; // @[TestHarness.scala 229:18]
  wire [63:0] _T_705 = _rob_tscs_T_31 - rob_tscs_63; // @[TestHarness.scala 229:18]
  wire [63:0] _T_712 = _rob_tscs_T_31 - rob_tscs_64; // @[TestHarness.scala 229:18]
  wire [63:0] _T_719 = _rob_tscs_T_31 - rob_tscs_65; // @[TestHarness.scala 229:18]
  wire [63:0] _T_726 = _rob_tscs_T_31 - rob_tscs_66; // @[TestHarness.scala 229:18]
  wire [63:0] _T_733 = _rob_tscs_T_31 - rob_tscs_67; // @[TestHarness.scala 229:18]
  wire [63:0] _T_740 = _rob_tscs_T_31 - rob_tscs_68; // @[TestHarness.scala 229:18]
  wire [63:0] _T_747 = _rob_tscs_T_31 - rob_tscs_69; // @[TestHarness.scala 229:18]
  wire [63:0] _T_754 = _rob_tscs_T_31 - rob_tscs_70; // @[TestHarness.scala 229:18]
  wire [63:0] _T_761 = _rob_tscs_T_31 - rob_tscs_71; // @[TestHarness.scala 229:18]
  wire [63:0] _T_768 = _rob_tscs_T_31 - rob_tscs_72; // @[TestHarness.scala 229:18]
  wire [63:0] _T_775 = _rob_tscs_T_31 - rob_tscs_73; // @[TestHarness.scala 229:18]
  wire [63:0] _T_782 = _rob_tscs_T_31 - rob_tscs_74; // @[TestHarness.scala 229:18]
  wire [63:0] _T_789 = _rob_tscs_T_31 - rob_tscs_75; // @[TestHarness.scala 229:18]
  wire [63:0] _T_796 = _rob_tscs_T_31 - rob_tscs_76; // @[TestHarness.scala 229:18]
  wire [63:0] _T_803 = _rob_tscs_T_31 - rob_tscs_77; // @[TestHarness.scala 229:18]
  wire [63:0] _T_810 = _rob_tscs_T_31 - rob_tscs_78; // @[TestHarness.scala 229:18]
  wire [63:0] _T_817 = _rob_tscs_T_31 - rob_tscs_79; // @[TestHarness.scala 229:18]
  wire [63:0] _T_824 = _rob_tscs_T_31 - rob_tscs_80; // @[TestHarness.scala 229:18]
  wire [63:0] _T_831 = _rob_tscs_T_31 - rob_tscs_81; // @[TestHarness.scala 229:18]
  wire [63:0] _T_838 = _rob_tscs_T_31 - rob_tscs_82; // @[TestHarness.scala 229:18]
  wire [63:0] _T_845 = _rob_tscs_T_31 - rob_tscs_83; // @[TestHarness.scala 229:18]
  wire [63:0] _T_852 = _rob_tscs_T_31 - rob_tscs_84; // @[TestHarness.scala 229:18]
  wire [63:0] _T_859 = _rob_tscs_T_31 - rob_tscs_85; // @[TestHarness.scala 229:18]
  wire [63:0] _T_866 = _rob_tscs_T_31 - rob_tscs_86; // @[TestHarness.scala 229:18]
  wire [63:0] _T_873 = _rob_tscs_T_31 - rob_tscs_87; // @[TestHarness.scala 229:18]
  wire [63:0] _T_880 = _rob_tscs_T_31 - rob_tscs_88; // @[TestHarness.scala 229:18]
  wire [63:0] _T_887 = _rob_tscs_T_31 - rob_tscs_89; // @[TestHarness.scala 229:18]
  wire [63:0] _T_894 = _rob_tscs_T_31 - rob_tscs_90; // @[TestHarness.scala 229:18]
  wire [63:0] _T_901 = _rob_tscs_T_31 - rob_tscs_91; // @[TestHarness.scala 229:18]
  wire [63:0] _T_908 = _rob_tscs_T_31 - rob_tscs_92; // @[TestHarness.scala 229:18]
  wire [63:0] _T_915 = _rob_tscs_T_31 - rob_tscs_93; // @[TestHarness.scala 229:18]
  wire [63:0] _T_922 = _rob_tscs_T_31 - rob_tscs_94; // @[TestHarness.scala 229:18]
  wire [63:0] _T_929 = _rob_tscs_T_31 - rob_tscs_95; // @[TestHarness.scala 229:18]
  wire [63:0] _T_936 = _rob_tscs_T_31 - rob_tscs_96; // @[TestHarness.scala 229:18]
  wire [63:0] _T_943 = _rob_tscs_T_31 - rob_tscs_97; // @[TestHarness.scala 229:18]
  wire [63:0] _T_950 = _rob_tscs_T_31 - rob_tscs_98; // @[TestHarness.scala 229:18]
  wire [63:0] _T_957 = _rob_tscs_T_31 - rob_tscs_99; // @[TestHarness.scala 229:18]
  wire [63:0] _T_964 = _rob_tscs_T_31 - rob_tscs_100; // @[TestHarness.scala 229:18]
  wire [63:0] _T_971 = _rob_tscs_T_31 - rob_tscs_101; // @[TestHarness.scala 229:18]
  wire [63:0] _T_978 = _rob_tscs_T_31 - rob_tscs_102; // @[TestHarness.scala 229:18]
  wire [63:0] _T_985 = _rob_tscs_T_31 - rob_tscs_103; // @[TestHarness.scala 229:18]
  wire [63:0] _T_992 = _rob_tscs_T_31 - rob_tscs_104; // @[TestHarness.scala 229:18]
  wire [63:0] _T_999 = _rob_tscs_T_31 - rob_tscs_105; // @[TestHarness.scala 229:18]
  wire [63:0] _T_1006 = _rob_tscs_T_31 - rob_tscs_106; // @[TestHarness.scala 229:18]
  wire [63:0] _T_1013 = _rob_tscs_T_31 - rob_tscs_107; // @[TestHarness.scala 229:18]
  wire [63:0] _T_1020 = _rob_tscs_T_31 - rob_tscs_108; // @[TestHarness.scala 229:18]
  wire [63:0] _T_1027 = _rob_tscs_T_31 - rob_tscs_109; // @[TestHarness.scala 229:18]
  wire [63:0] _T_1034 = _rob_tscs_T_31 - rob_tscs_110; // @[TestHarness.scala 229:18]
  wire [63:0] _T_1041 = _rob_tscs_T_31 - rob_tscs_111; // @[TestHarness.scala 229:18]
  wire [63:0] _T_1048 = _rob_tscs_T_31 - rob_tscs_112; // @[TestHarness.scala 229:18]
  wire [63:0] _T_1055 = _rob_tscs_T_31 - rob_tscs_113; // @[TestHarness.scala 229:18]
  wire [63:0] _T_1062 = _rob_tscs_T_31 - rob_tscs_114; // @[TestHarness.scala 229:18]
  wire [63:0] _T_1069 = _rob_tscs_T_31 - rob_tscs_115; // @[TestHarness.scala 229:18]
  wire [63:0] _T_1076 = _rob_tscs_T_31 - rob_tscs_116; // @[TestHarness.scala 229:18]
  wire [63:0] _T_1083 = _rob_tscs_T_31 - rob_tscs_117; // @[TestHarness.scala 229:18]
  wire [63:0] _T_1090 = _rob_tscs_T_31 - rob_tscs_118; // @[TestHarness.scala 229:18]
  wire [63:0] _T_1097 = _rob_tscs_T_31 - rob_tscs_119; // @[TestHarness.scala 229:18]
  wire [63:0] _T_1104 = _rob_tscs_T_31 - rob_tscs_120; // @[TestHarness.scala 229:18]
  wire [63:0] _T_1111 = _rob_tscs_T_31 - rob_tscs_121; // @[TestHarness.scala 229:18]
  wire [63:0] _T_1118 = _rob_tscs_T_31 - rob_tscs_122; // @[TestHarness.scala 229:18]
  wire [63:0] _T_1125 = _rob_tscs_T_31 - rob_tscs_123; // @[TestHarness.scala 229:18]
  wire [63:0] _T_1132 = _rob_tscs_T_31 - rob_tscs_124; // @[TestHarness.scala 229:18]
  wire [63:0] _T_1139 = _rob_tscs_T_31 - rob_tscs_125; // @[TestHarness.scala 229:18]
  wire [63:0] _T_1146 = _rob_tscs_T_31 - rob_tscs_126; // @[TestHarness.scala 229:18]
  wire [63:0] _T_1153 = _rob_tscs_T_31 - rob_tscs_127; // @[TestHarness.scala 229:18]
  wire [65535:0] _GEN_15518 = reset ? 65536'h0 : _rob_valids_T_2; // @[TestHarness.scala 156:{27,27} 222:14]
  wire  _GEN_15519 = _T_118 & _T_3; // @[TestHarness.scala 201:13]
  wire  _GEN_15526 = _T_165 & _T_3; // @[TestHarness.scala 201:13]
  wire  _GEN_15533 = _T_212 & _T_3; // @[TestHarness.scala 201:13]
  wire  _GEN_15540 = _T_259 & _T_3; // @[TestHarness.scala 201:13]
  InputGen igen ( // @[TestHarness.scala 171:22]
    .clock(igen_clock),
    .reset(igen_reset),
    .io_out_ready(igen_io_out_ready),
    .io_out_valid(igen_io_out_valid),
    .io_out_bits_head(igen_io_out_bits_head),
    .io_out_bits_tail(igen_io_out_bits_tail),
    .io_out_bits_payload(igen_io_out_bits_payload),
    .io_out_bits_egress_id(igen_io_out_bits_egress_id),
    .io_rob_ready(igen_io_rob_ready),
    .io_rob_idx(igen_io_rob_idx),
    .io_tsc(igen_io_tsc),
    .io_fire(igen_io_fire),
    .io_n_flits(igen_io_n_flits)
  );
  Queue_52 io_to_noc_0_flit_q ( // @[Decoupled.scala 375:21]
    .clock(io_to_noc_0_flit_q_clock),
    .reset(io_to_noc_0_flit_q_reset),
    .io_enq_ready(io_to_noc_0_flit_q_io_enq_ready),
    .io_enq_valid(io_to_noc_0_flit_q_io_enq_valid),
    .io_enq_bits_head(io_to_noc_0_flit_q_io_enq_bits_head),
    .io_enq_bits_tail(io_to_noc_0_flit_q_io_enq_bits_tail),
    .io_enq_bits_payload(io_to_noc_0_flit_q_io_enq_bits_payload),
    .io_enq_bits_egress_id(io_to_noc_0_flit_q_io_enq_bits_egress_id),
    .io_deq_ready(io_to_noc_0_flit_q_io_deq_ready),
    .io_deq_valid(io_to_noc_0_flit_q_io_deq_valid),
    .io_deq_bits_head(io_to_noc_0_flit_q_io_deq_bits_head),
    .io_deq_bits_tail(io_to_noc_0_flit_q_io_deq_bits_tail),
    .io_deq_bits_payload(io_to_noc_0_flit_q_io_deq_bits_payload),
    .io_deq_bits_egress_id(io_to_noc_0_flit_q_io_deq_bits_egress_id)
  );
  InputGen igen_1 ( // @[TestHarness.scala 171:22]
    .clock(igen_1_clock),
    .reset(igen_1_reset),
    .io_out_ready(igen_1_io_out_ready),
    .io_out_valid(igen_1_io_out_valid),
    .io_out_bits_head(igen_1_io_out_bits_head),
    .io_out_bits_tail(igen_1_io_out_bits_tail),
    .io_out_bits_payload(igen_1_io_out_bits_payload),
    .io_out_bits_egress_id(igen_1_io_out_bits_egress_id),
    .io_rob_ready(igen_1_io_rob_ready),
    .io_rob_idx(igen_1_io_rob_idx),
    .io_tsc(igen_1_io_tsc),
    .io_fire(igen_1_io_fire),
    .io_n_flits(igen_1_io_n_flits)
  );
  Queue_52 io_to_noc_1_flit_q ( // @[Decoupled.scala 375:21]
    .clock(io_to_noc_1_flit_q_clock),
    .reset(io_to_noc_1_flit_q_reset),
    .io_enq_ready(io_to_noc_1_flit_q_io_enq_ready),
    .io_enq_valid(io_to_noc_1_flit_q_io_enq_valid),
    .io_enq_bits_head(io_to_noc_1_flit_q_io_enq_bits_head),
    .io_enq_bits_tail(io_to_noc_1_flit_q_io_enq_bits_tail),
    .io_enq_bits_payload(io_to_noc_1_flit_q_io_enq_bits_payload),
    .io_enq_bits_egress_id(io_to_noc_1_flit_q_io_enq_bits_egress_id),
    .io_deq_ready(io_to_noc_1_flit_q_io_deq_ready),
    .io_deq_valid(io_to_noc_1_flit_q_io_deq_valid),
    .io_deq_bits_head(io_to_noc_1_flit_q_io_deq_bits_head),
    .io_deq_bits_tail(io_to_noc_1_flit_q_io_deq_bits_tail),
    .io_deq_bits_payload(io_to_noc_1_flit_q_io_deq_bits_payload),
    .io_deq_bits_egress_id(io_to_noc_1_flit_q_io_deq_bits_egress_id)
  );
  InputGen igen_2 ( // @[TestHarness.scala 171:22]
    .clock(igen_2_clock),
    .reset(igen_2_reset),
    .io_out_ready(igen_2_io_out_ready),
    .io_out_valid(igen_2_io_out_valid),
    .io_out_bits_head(igen_2_io_out_bits_head),
    .io_out_bits_tail(igen_2_io_out_bits_tail),
    .io_out_bits_payload(igen_2_io_out_bits_payload),
    .io_out_bits_egress_id(igen_2_io_out_bits_egress_id),
    .io_rob_ready(igen_2_io_rob_ready),
    .io_rob_idx(igen_2_io_rob_idx),
    .io_tsc(igen_2_io_tsc),
    .io_fire(igen_2_io_fire),
    .io_n_flits(igen_2_io_n_flits)
  );
  Queue_52 io_to_noc_2_flit_q ( // @[Decoupled.scala 375:21]
    .clock(io_to_noc_2_flit_q_clock),
    .reset(io_to_noc_2_flit_q_reset),
    .io_enq_ready(io_to_noc_2_flit_q_io_enq_ready),
    .io_enq_valid(io_to_noc_2_flit_q_io_enq_valid),
    .io_enq_bits_head(io_to_noc_2_flit_q_io_enq_bits_head),
    .io_enq_bits_tail(io_to_noc_2_flit_q_io_enq_bits_tail),
    .io_enq_bits_payload(io_to_noc_2_flit_q_io_enq_bits_payload),
    .io_enq_bits_egress_id(io_to_noc_2_flit_q_io_enq_bits_egress_id),
    .io_deq_ready(io_to_noc_2_flit_q_io_deq_ready),
    .io_deq_valid(io_to_noc_2_flit_q_io_deq_valid),
    .io_deq_bits_head(io_to_noc_2_flit_q_io_deq_bits_head),
    .io_deq_bits_tail(io_to_noc_2_flit_q_io_deq_bits_tail),
    .io_deq_bits_payload(io_to_noc_2_flit_q_io_deq_bits_payload),
    .io_deq_bits_egress_id(io_to_noc_2_flit_q_io_deq_bits_egress_id)
  );
  InputGen igen_3 ( // @[TestHarness.scala 171:22]
    .clock(igen_3_clock),
    .reset(igen_3_reset),
    .io_out_ready(igen_3_io_out_ready),
    .io_out_valid(igen_3_io_out_valid),
    .io_out_bits_head(igen_3_io_out_bits_head),
    .io_out_bits_tail(igen_3_io_out_bits_tail),
    .io_out_bits_payload(igen_3_io_out_bits_payload),
    .io_out_bits_egress_id(igen_3_io_out_bits_egress_id),
    .io_rob_ready(igen_3_io_rob_ready),
    .io_rob_idx(igen_3_io_rob_idx),
    .io_tsc(igen_3_io_tsc),
    .io_fire(igen_3_io_fire),
    .io_n_flits(igen_3_io_n_flits)
  );
  Queue_52 io_to_noc_3_flit_q ( // @[Decoupled.scala 375:21]
    .clock(io_to_noc_3_flit_q_clock),
    .reset(io_to_noc_3_flit_q_reset),
    .io_enq_ready(io_to_noc_3_flit_q_io_enq_ready),
    .io_enq_valid(io_to_noc_3_flit_q_io_enq_valid),
    .io_enq_bits_head(io_to_noc_3_flit_q_io_enq_bits_head),
    .io_enq_bits_tail(io_to_noc_3_flit_q_io_enq_bits_tail),
    .io_enq_bits_payload(io_to_noc_3_flit_q_io_enq_bits_payload),
    .io_enq_bits_egress_id(io_to_noc_3_flit_q_io_enq_bits_egress_id),
    .io_deq_ready(io_to_noc_3_flit_q_io_deq_ready),
    .io_deq_valid(io_to_noc_3_flit_q_io_deq_valid),
    .io_deq_bits_head(io_to_noc_3_flit_q_io_deq_bits_head),
    .io_deq_bits_tail(io_to_noc_3_flit_q_io_deq_bits_tail),
    .io_deq_bits_payload(io_to_noc_3_flit_q_io_deq_bits_payload),
    .io_deq_bits_egress_id(io_to_noc_3_flit_q_io_deq_bits_egress_id)
  );
  plusarg_reader #(.FORMAT("noctest_enable_print=%d"), .DEFAULT(0), .WIDTH(1)) plusarg_reader ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_out)
  );
  MaxPeriodFibonacciLFSR io_from_noc_0_flit_ready_prng ( // @[PRNG.scala 91:22]
    .clock(io_from_noc_0_flit_ready_prng_clock),
    .reset(io_from_noc_0_flit_ready_prng_reset),
    .io_out_0(io_from_noc_0_flit_ready_prng_io_out_0),
    .io_out_1(io_from_noc_0_flit_ready_prng_io_out_1),
    .io_out_2(io_from_noc_0_flit_ready_prng_io_out_2),
    .io_out_3(io_from_noc_0_flit_ready_prng_io_out_3),
    .io_out_4(io_from_noc_0_flit_ready_prng_io_out_4),
    .io_out_5(io_from_noc_0_flit_ready_prng_io_out_5),
    .io_out_6(io_from_noc_0_flit_ready_prng_io_out_6),
    .io_out_7(io_from_noc_0_flit_ready_prng_io_out_7),
    .io_out_8(io_from_noc_0_flit_ready_prng_io_out_8),
    .io_out_9(io_from_noc_0_flit_ready_prng_io_out_9),
    .io_out_10(io_from_noc_0_flit_ready_prng_io_out_10),
    .io_out_11(io_from_noc_0_flit_ready_prng_io_out_11),
    .io_out_12(io_from_noc_0_flit_ready_prng_io_out_12),
    .io_out_13(io_from_noc_0_flit_ready_prng_io_out_13),
    .io_out_14(io_from_noc_0_flit_ready_prng_io_out_14),
    .io_out_15(io_from_noc_0_flit_ready_prng_io_out_15),
    .io_out_16(io_from_noc_0_flit_ready_prng_io_out_16),
    .io_out_17(io_from_noc_0_flit_ready_prng_io_out_17),
    .io_out_18(io_from_noc_0_flit_ready_prng_io_out_18),
    .io_out_19(io_from_noc_0_flit_ready_prng_io_out_19)
  );
  MaxPeriodFibonacciLFSR io_from_noc_1_flit_ready_prng ( // @[PRNG.scala 91:22]
    .clock(io_from_noc_1_flit_ready_prng_clock),
    .reset(io_from_noc_1_flit_ready_prng_reset),
    .io_out_0(io_from_noc_1_flit_ready_prng_io_out_0),
    .io_out_1(io_from_noc_1_flit_ready_prng_io_out_1),
    .io_out_2(io_from_noc_1_flit_ready_prng_io_out_2),
    .io_out_3(io_from_noc_1_flit_ready_prng_io_out_3),
    .io_out_4(io_from_noc_1_flit_ready_prng_io_out_4),
    .io_out_5(io_from_noc_1_flit_ready_prng_io_out_5),
    .io_out_6(io_from_noc_1_flit_ready_prng_io_out_6),
    .io_out_7(io_from_noc_1_flit_ready_prng_io_out_7),
    .io_out_8(io_from_noc_1_flit_ready_prng_io_out_8),
    .io_out_9(io_from_noc_1_flit_ready_prng_io_out_9),
    .io_out_10(io_from_noc_1_flit_ready_prng_io_out_10),
    .io_out_11(io_from_noc_1_flit_ready_prng_io_out_11),
    .io_out_12(io_from_noc_1_flit_ready_prng_io_out_12),
    .io_out_13(io_from_noc_1_flit_ready_prng_io_out_13),
    .io_out_14(io_from_noc_1_flit_ready_prng_io_out_14),
    .io_out_15(io_from_noc_1_flit_ready_prng_io_out_15),
    .io_out_16(io_from_noc_1_flit_ready_prng_io_out_16),
    .io_out_17(io_from_noc_1_flit_ready_prng_io_out_17),
    .io_out_18(io_from_noc_1_flit_ready_prng_io_out_18),
    .io_out_19(io_from_noc_1_flit_ready_prng_io_out_19)
  );
  MaxPeriodFibonacciLFSR io_from_noc_2_flit_ready_prng ( // @[PRNG.scala 91:22]
    .clock(io_from_noc_2_flit_ready_prng_clock),
    .reset(io_from_noc_2_flit_ready_prng_reset),
    .io_out_0(io_from_noc_2_flit_ready_prng_io_out_0),
    .io_out_1(io_from_noc_2_flit_ready_prng_io_out_1),
    .io_out_2(io_from_noc_2_flit_ready_prng_io_out_2),
    .io_out_3(io_from_noc_2_flit_ready_prng_io_out_3),
    .io_out_4(io_from_noc_2_flit_ready_prng_io_out_4),
    .io_out_5(io_from_noc_2_flit_ready_prng_io_out_5),
    .io_out_6(io_from_noc_2_flit_ready_prng_io_out_6),
    .io_out_7(io_from_noc_2_flit_ready_prng_io_out_7),
    .io_out_8(io_from_noc_2_flit_ready_prng_io_out_8),
    .io_out_9(io_from_noc_2_flit_ready_prng_io_out_9),
    .io_out_10(io_from_noc_2_flit_ready_prng_io_out_10),
    .io_out_11(io_from_noc_2_flit_ready_prng_io_out_11),
    .io_out_12(io_from_noc_2_flit_ready_prng_io_out_12),
    .io_out_13(io_from_noc_2_flit_ready_prng_io_out_13),
    .io_out_14(io_from_noc_2_flit_ready_prng_io_out_14),
    .io_out_15(io_from_noc_2_flit_ready_prng_io_out_15),
    .io_out_16(io_from_noc_2_flit_ready_prng_io_out_16),
    .io_out_17(io_from_noc_2_flit_ready_prng_io_out_17),
    .io_out_18(io_from_noc_2_flit_ready_prng_io_out_18),
    .io_out_19(io_from_noc_2_flit_ready_prng_io_out_19)
  );
  MaxPeriodFibonacciLFSR io_from_noc_3_flit_ready_prng ( // @[PRNG.scala 91:22]
    .clock(io_from_noc_3_flit_ready_prng_clock),
    .reset(io_from_noc_3_flit_ready_prng_reset),
    .io_out_0(io_from_noc_3_flit_ready_prng_io_out_0),
    .io_out_1(io_from_noc_3_flit_ready_prng_io_out_1),
    .io_out_2(io_from_noc_3_flit_ready_prng_io_out_2),
    .io_out_3(io_from_noc_3_flit_ready_prng_io_out_3),
    .io_out_4(io_from_noc_3_flit_ready_prng_io_out_4),
    .io_out_5(io_from_noc_3_flit_ready_prng_io_out_5),
    .io_out_6(io_from_noc_3_flit_ready_prng_io_out_6),
    .io_out_7(io_from_noc_3_flit_ready_prng_io_out_7),
    .io_out_8(io_from_noc_3_flit_ready_prng_io_out_8),
    .io_out_9(io_from_noc_3_flit_ready_prng_io_out_9),
    .io_out_10(io_from_noc_3_flit_ready_prng_io_out_10),
    .io_out_11(io_from_noc_3_flit_ready_prng_io_out_11),
    .io_out_12(io_from_noc_3_flit_ready_prng_io_out_12),
    .io_out_13(io_from_noc_3_flit_ready_prng_io_out_13),
    .io_out_14(io_from_noc_3_flit_ready_prng_io_out_14),
    .io_out_15(io_from_noc_3_flit_ready_prng_io_out_15),
    .io_out_16(io_from_noc_3_flit_ready_prng_io_out_16),
    .io_out_17(io_from_noc_3_flit_ready_prng_io_out_17),
    .io_out_18(io_from_noc_3_flit_ready_prng_io_out_18),
    .io_out_19(io_from_noc_3_flit_ready_prng_io_out_19)
  );
  assign io_to_noc_3_flit_valid = io_to_noc_3_flit_q_io_deq_valid; // @[TestHarness.scala 177:12]
  assign io_to_noc_3_flit_bits_head = io_to_noc_3_flit_q_io_deq_bits_head; // @[TestHarness.scala 177:12]
  assign io_to_noc_3_flit_bits_tail = io_to_noc_3_flit_q_io_deq_bits_tail; // @[TestHarness.scala 177:12]
  assign io_to_noc_3_flit_bits_payload = io_to_noc_3_flit_q_io_deq_bits_payload; // @[TestHarness.scala 177:12]
  assign io_to_noc_3_flit_bits_egress_id = io_to_noc_3_flit_q_io_deq_bits_egress_id; // @[TestHarness.scala 177:12]
  assign io_to_noc_2_flit_valid = io_to_noc_2_flit_q_io_deq_valid; // @[TestHarness.scala 177:12]
  assign io_to_noc_2_flit_bits_head = io_to_noc_2_flit_q_io_deq_bits_head; // @[TestHarness.scala 177:12]
  assign io_to_noc_2_flit_bits_tail = io_to_noc_2_flit_q_io_deq_bits_tail; // @[TestHarness.scala 177:12]
  assign io_to_noc_2_flit_bits_payload = io_to_noc_2_flit_q_io_deq_bits_payload; // @[TestHarness.scala 177:12]
  assign io_to_noc_2_flit_bits_egress_id = io_to_noc_2_flit_q_io_deq_bits_egress_id; // @[TestHarness.scala 177:12]
  assign io_to_noc_1_flit_valid = io_to_noc_1_flit_q_io_deq_valid; // @[TestHarness.scala 177:12]
  assign io_to_noc_1_flit_bits_head = io_to_noc_1_flit_q_io_deq_bits_head; // @[TestHarness.scala 177:12]
  assign io_to_noc_1_flit_bits_tail = io_to_noc_1_flit_q_io_deq_bits_tail; // @[TestHarness.scala 177:12]
  assign io_to_noc_1_flit_bits_payload = io_to_noc_1_flit_q_io_deq_bits_payload; // @[TestHarness.scala 177:12]
  assign io_to_noc_1_flit_bits_egress_id = io_to_noc_1_flit_q_io_deq_bits_egress_id; // @[TestHarness.scala 177:12]
  assign io_to_noc_0_flit_valid = io_to_noc_0_flit_q_io_deq_valid; // @[TestHarness.scala 177:12]
  assign io_to_noc_0_flit_bits_head = io_to_noc_0_flit_q_io_deq_bits_head; // @[TestHarness.scala 177:12]
  assign io_to_noc_0_flit_bits_tail = io_to_noc_0_flit_q_io_deq_bits_tail; // @[TestHarness.scala 177:12]
  assign io_to_noc_0_flit_bits_payload = io_to_noc_0_flit_q_io_deq_bits_payload; // @[TestHarness.scala 177:12]
  assign io_to_noc_0_flit_bits_egress_id = io_to_noc_0_flit_q_io_deq_bits_egress_id; // @[TestHarness.scala 177:12]
  assign io_from_noc_3_flit_ready = 1'h1; // @[TestHarness.scala 193:30]
  assign io_from_noc_2_flit_ready = 1'h1; // @[TestHarness.scala 193:30]
  assign io_from_noc_1_flit_ready = 1'h1; // @[TestHarness.scala 193:30]
  assign io_from_noc_0_flit_ready = 1'h1; // @[TestHarness.scala 193:30]
  assign io_success = io_success_REG; // @[TestHarness.scala 164:14]
  assign igen_clock = clock;
  assign igen_reset = reset;
  assign igen_io_out_ready = io_to_noc_0_flit_q_io_enq_ready; // @[Decoupled.scala 379:17]
  assign igen_io_rob_ready = _igen_io_rob_ready_T_2 & txs < 32'hc350; // @[TestHarness.scala 175:19]
  assign igen_io_rob_idx = _T_5[0] ? 7'h0 : _sels_0_T_253; // @[Mux.scala 47:70]
  assign igen_io_tsc = tsc; // @[TestHarness.scala 176:17]
  assign io_to_noc_0_flit_q_clock = clock;
  assign io_to_noc_0_flit_q_reset = reset;
  assign io_to_noc_0_flit_q_io_enq_valid = igen_io_out_valid; // @[Decoupled.scala 377:22]
  assign io_to_noc_0_flit_q_io_enq_bits_head = igen_io_out_bits_head; // @[Decoupled.scala 378:21]
  assign io_to_noc_0_flit_q_io_enq_bits_tail = igen_io_out_bits_tail; // @[Decoupled.scala 378:21]
  assign io_to_noc_0_flit_q_io_enq_bits_payload = igen_io_out_bits_payload; // @[Decoupled.scala 378:21]
  assign io_to_noc_0_flit_q_io_enq_bits_egress_id = igen_io_out_bits_egress_id; // @[Decoupled.scala 378:21]
  assign io_to_noc_0_flit_q_io_deq_ready = io_to_noc_0_flit_ready; // @[TestHarness.scala 177:12]
  assign igen_1_clock = clock;
  assign igen_1_reset = reset;
  assign igen_1_io_out_ready = io_to_noc_1_flit_q_io_enq_ready; // @[Decoupled.scala 379:17]
  assign igen_1_io_rob_ready = _igen_io_rob_ready_T_7 & txs < 32'hc350; // @[TestHarness.scala 175:19]
  assign igen_1_io_rob_idx = _T_8[0] ? 7'h0 : _sels_1_T_253; // @[Mux.scala 47:70]
  assign igen_1_io_tsc = tsc; // @[TestHarness.scala 176:17]
  assign io_to_noc_1_flit_q_clock = clock;
  assign io_to_noc_1_flit_q_reset = reset;
  assign io_to_noc_1_flit_q_io_enq_valid = igen_1_io_out_valid; // @[Decoupled.scala 377:22]
  assign io_to_noc_1_flit_q_io_enq_bits_head = igen_1_io_out_bits_head; // @[Decoupled.scala 378:21]
  assign io_to_noc_1_flit_q_io_enq_bits_tail = igen_1_io_out_bits_tail; // @[Decoupled.scala 378:21]
  assign io_to_noc_1_flit_q_io_enq_bits_payload = igen_1_io_out_bits_payload; // @[Decoupled.scala 378:21]
  assign io_to_noc_1_flit_q_io_enq_bits_egress_id = igen_1_io_out_bits_egress_id; // @[Decoupled.scala 378:21]
  assign io_to_noc_1_flit_q_io_deq_ready = io_to_noc_1_flit_ready; // @[TestHarness.scala 177:12]
  assign igen_2_clock = clock;
  assign igen_2_reset = reset;
  assign igen_2_io_out_ready = io_to_noc_2_flit_q_io_enq_ready; // @[Decoupled.scala 379:17]
  assign igen_2_io_rob_ready = _igen_io_rob_ready_T_12 & txs < 32'hc350; // @[TestHarness.scala 175:19]
  assign igen_2_io_rob_idx = _T_11[0] ? 7'h0 : _sels_2_T_253; // @[Mux.scala 47:70]
  assign igen_2_io_tsc = tsc; // @[TestHarness.scala 176:17]
  assign io_to_noc_2_flit_q_clock = clock;
  assign io_to_noc_2_flit_q_reset = reset;
  assign io_to_noc_2_flit_q_io_enq_valid = igen_2_io_out_valid; // @[Decoupled.scala 377:22]
  assign io_to_noc_2_flit_q_io_enq_bits_head = igen_2_io_out_bits_head; // @[Decoupled.scala 378:21]
  assign io_to_noc_2_flit_q_io_enq_bits_tail = igen_2_io_out_bits_tail; // @[Decoupled.scala 378:21]
  assign io_to_noc_2_flit_q_io_enq_bits_payload = igen_2_io_out_bits_payload; // @[Decoupled.scala 378:21]
  assign io_to_noc_2_flit_q_io_enq_bits_egress_id = igen_2_io_out_bits_egress_id; // @[Decoupled.scala 378:21]
  assign io_to_noc_2_flit_q_io_deq_ready = io_to_noc_2_flit_ready; // @[TestHarness.scala 177:12]
  assign igen_3_clock = clock;
  assign igen_3_reset = reset;
  assign igen_3_io_out_ready = io_to_noc_3_flit_q_io_enq_ready; // @[Decoupled.scala 379:17]
  assign igen_3_io_rob_ready = _igen_io_rob_ready_T_17 & txs < 32'hc350; // @[TestHarness.scala 175:19]
  assign igen_3_io_rob_idx = _T_14[0] ? 7'h0 : _sels_3_T_253; // @[Mux.scala 47:70]
  assign igen_3_io_tsc = tsc; // @[TestHarness.scala 176:17]
  assign io_to_noc_3_flit_q_clock = clock;
  assign io_to_noc_3_flit_q_reset = reset;
  assign io_to_noc_3_flit_q_io_enq_valid = igen_3_io_out_valid; // @[Decoupled.scala 377:22]
  assign io_to_noc_3_flit_q_io_enq_bits_head = igen_3_io_out_bits_head; // @[Decoupled.scala 378:21]
  assign io_to_noc_3_flit_q_io_enq_bits_tail = igen_3_io_out_bits_tail; // @[Decoupled.scala 378:21]
  assign io_to_noc_3_flit_q_io_enq_bits_payload = igen_3_io_out_bits_payload; // @[Decoupled.scala 378:21]
  assign io_to_noc_3_flit_q_io_enq_bits_egress_id = igen_3_io_out_bits_egress_id; // @[Decoupled.scala 378:21]
  assign io_to_noc_3_flit_q_io_deq_ready = io_to_noc_3_flit_ready; // @[TestHarness.scala 177:12]
  assign io_from_noc_0_flit_ready_prng_clock = clock;
  assign io_from_noc_0_flit_ready_prng_reset = reset;
  assign io_from_noc_1_flit_ready_prng_clock = clock;
  assign io_from_noc_1_flit_ready_prng_reset = reset;
  assign io_from_noc_2_flit_ready_prng_clock = clock;
  assign io_from_noc_2_flit_ready_prng_reset = reset;
  assign io_from_noc_3_flit_ready_prng_clock = clock;
  assign io_from_noc_3_flit_ready_prng_reset = reset;
  always @(posedge clock) begin
    if (reset) begin // @[TestHarness.scala 136:20]
      txs <= 32'h0; // @[TestHarness.scala 136:20]
    end else begin
      txs <= _txs_T_7; // @[TestHarness.scala 225:7]
    end
    if (reset) begin // @[TestHarness.scala 137:22]
      flits <= 32'h0; // @[TestHarness.scala 137:22]
    end else begin
      flits <= _flits_T_8; // @[TestHarness.scala 224:9]
    end
    if (reset) begin // @[TestHarness.scala 141:20]
      tsc <= 32'h0; // @[TestHarness.scala 141:20]
    end else begin
      tsc <= _tsc_T_1; // @[TestHarness.scala 142:7]
    end
    if (reset) begin // @[TestHarness.scala 144:29]
      idle_counter <= 11'h0; // @[TestHarness.scala 144:29]
    end else if (idle) begin // @[TestHarness.scala 146:15]
      idle_counter <= _idle_counter_T_1; // @[TestHarness.scala 146:30]
    end else begin
      idle_counter <= 11'h0; // @[TestHarness.scala 147:31]
    end
    rob_valids <= _GEN_15518[127:0]; // @[TestHarness.scala 156:{27,27} 222:14]
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h0 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_0_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_0_tsc <= _GEN_5121;
      end
    end else begin
      rob_payload_0_tsc <= _GEN_5121;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h0 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_0_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_0_rob_idx <= _GEN_5249;
      end
    end else begin
      rob_payload_0_rob_idx <= _GEN_5249;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h0 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_0_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_0_flits_fired <= _GEN_13454;
      end
    end else begin
      rob_payload_0_flits_fired <= _GEN_13454;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_1_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_1_tsc <= _GEN_5122;
      end
    end else begin
      rob_payload_1_tsc <= _GEN_5122;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_1_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_1_rob_idx <= _GEN_5250;
      end
    end else begin
      rob_payload_1_rob_idx <= _GEN_5250;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h1 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_1_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_1_flits_fired <= _GEN_13455;
      end
    end else begin
      rob_payload_1_flits_fired <= _GEN_13455;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_2_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_2_tsc <= _GEN_5123;
      end
    end else begin
      rob_payload_2_tsc <= _GEN_5123;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_2_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_2_rob_idx <= _GEN_5251;
      end
    end else begin
      rob_payload_2_rob_idx <= _GEN_5251;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h2 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_2_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_2_flits_fired <= _GEN_13456;
      end
    end else begin
      rob_payload_2_flits_fired <= _GEN_13456;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_3_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_3_tsc <= _GEN_5124;
      end
    end else begin
      rob_payload_3_tsc <= _GEN_5124;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_3_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_3_rob_idx <= _GEN_5252;
      end
    end else begin
      rob_payload_3_rob_idx <= _GEN_5252;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h3 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_3_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_3_flits_fired <= _GEN_13457;
      end
    end else begin
      rob_payload_3_flits_fired <= _GEN_13457;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_4_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_4_tsc <= _GEN_5125;
      end
    end else begin
      rob_payload_4_tsc <= _GEN_5125;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_4_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_4_rob_idx <= _GEN_5253;
      end
    end else begin
      rob_payload_4_rob_idx <= _GEN_5253;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h4 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_4_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_4_flits_fired <= _GEN_13458;
      end
    end else begin
      rob_payload_4_flits_fired <= _GEN_13458;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_5_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_5_tsc <= _GEN_5126;
      end
    end else begin
      rob_payload_5_tsc <= _GEN_5126;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_5_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_5_rob_idx <= _GEN_5254;
      end
    end else begin
      rob_payload_5_rob_idx <= _GEN_5254;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h5 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_5_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_5_flits_fired <= _GEN_13459;
      end
    end else begin
      rob_payload_5_flits_fired <= _GEN_13459;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_6_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_6_tsc <= _GEN_5127;
      end
    end else begin
      rob_payload_6_tsc <= _GEN_5127;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_6_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_6_rob_idx <= _GEN_5255;
      end
    end else begin
      rob_payload_6_rob_idx <= _GEN_5255;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h6 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_6_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_6_flits_fired <= _GEN_13460;
      end
    end else begin
      rob_payload_6_flits_fired <= _GEN_13460;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_7_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_7_tsc <= _GEN_5128;
      end
    end else begin
      rob_payload_7_tsc <= _GEN_5128;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_7_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_7_rob_idx <= _GEN_5256;
      end
    end else begin
      rob_payload_7_rob_idx <= _GEN_5256;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h7 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_7_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_7_flits_fired <= _GEN_13461;
      end
    end else begin
      rob_payload_7_flits_fired <= _GEN_13461;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h8 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_8_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_8_tsc <= _GEN_5129;
      end
    end else begin
      rob_payload_8_tsc <= _GEN_5129;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h8 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_8_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_8_rob_idx <= _GEN_5257;
      end
    end else begin
      rob_payload_8_rob_idx <= _GEN_5257;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h8 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_8_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_8_flits_fired <= _GEN_13462;
      end
    end else begin
      rob_payload_8_flits_fired <= _GEN_13462;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h9 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_9_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_9_tsc <= _GEN_5130;
      end
    end else begin
      rob_payload_9_tsc <= _GEN_5130;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h9 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_9_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_9_rob_idx <= _GEN_5258;
      end
    end else begin
      rob_payload_9_rob_idx <= _GEN_5258;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h9 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_9_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_9_flits_fired <= _GEN_13463;
      end
    end else begin
      rob_payload_9_flits_fired <= _GEN_13463;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'ha == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_10_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_10_tsc <= _GEN_5131;
      end
    end else begin
      rob_payload_10_tsc <= _GEN_5131;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'ha == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_10_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_10_rob_idx <= _GEN_5259;
      end
    end else begin
      rob_payload_10_rob_idx <= _GEN_5259;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'ha == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_10_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_10_flits_fired <= _GEN_13464;
      end
    end else begin
      rob_payload_10_flits_fired <= _GEN_13464;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hb == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_11_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_11_tsc <= _GEN_5132;
      end
    end else begin
      rob_payload_11_tsc <= _GEN_5132;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hb == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_11_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_11_rob_idx <= _GEN_5260;
      end
    end else begin
      rob_payload_11_rob_idx <= _GEN_5260;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'hb == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_11_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_11_flits_fired <= _GEN_13465;
      end
    end else begin
      rob_payload_11_flits_fired <= _GEN_13465;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hc == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_12_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_12_tsc <= _GEN_5133;
      end
    end else begin
      rob_payload_12_tsc <= _GEN_5133;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hc == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_12_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_12_rob_idx <= _GEN_5261;
      end
    end else begin
      rob_payload_12_rob_idx <= _GEN_5261;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'hc == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_12_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_12_flits_fired <= _GEN_13466;
      end
    end else begin
      rob_payload_12_flits_fired <= _GEN_13466;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hd == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_13_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_13_tsc <= _GEN_5134;
      end
    end else begin
      rob_payload_13_tsc <= _GEN_5134;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hd == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_13_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_13_rob_idx <= _GEN_5262;
      end
    end else begin
      rob_payload_13_rob_idx <= _GEN_5262;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'hd == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_13_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_13_flits_fired <= _GEN_13467;
      end
    end else begin
      rob_payload_13_flits_fired <= _GEN_13467;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'he == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_14_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_14_tsc <= _GEN_5135;
      end
    end else begin
      rob_payload_14_tsc <= _GEN_5135;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'he == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_14_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_14_rob_idx <= _GEN_5263;
      end
    end else begin
      rob_payload_14_rob_idx <= _GEN_5263;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'he == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_14_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_14_flits_fired <= _GEN_13468;
      end
    end else begin
      rob_payload_14_flits_fired <= _GEN_13468;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hf == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_15_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_15_tsc <= _GEN_5136;
      end
    end else begin
      rob_payload_15_tsc <= _GEN_5136;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hf == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_15_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_15_rob_idx <= _GEN_5264;
      end
    end else begin
      rob_payload_15_rob_idx <= _GEN_5264;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'hf == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_15_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_15_flits_fired <= _GEN_13469;
      end
    end else begin
      rob_payload_15_flits_fired <= _GEN_13469;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h10 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_16_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_16_tsc <= _GEN_5137;
      end
    end else begin
      rob_payload_16_tsc <= _GEN_5137;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h10 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_16_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_16_rob_idx <= _GEN_5265;
      end
    end else begin
      rob_payload_16_rob_idx <= _GEN_5265;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h10 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_16_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_16_flits_fired <= _GEN_13470;
      end
    end else begin
      rob_payload_16_flits_fired <= _GEN_13470;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h11 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_17_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_17_tsc <= _GEN_5138;
      end
    end else begin
      rob_payload_17_tsc <= _GEN_5138;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h11 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_17_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_17_rob_idx <= _GEN_5266;
      end
    end else begin
      rob_payload_17_rob_idx <= _GEN_5266;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h11 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_17_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_17_flits_fired <= _GEN_13471;
      end
    end else begin
      rob_payload_17_flits_fired <= _GEN_13471;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h12 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_18_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_18_tsc <= _GEN_5139;
      end
    end else begin
      rob_payload_18_tsc <= _GEN_5139;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h12 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_18_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_18_rob_idx <= _GEN_5267;
      end
    end else begin
      rob_payload_18_rob_idx <= _GEN_5267;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h12 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_18_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_18_flits_fired <= _GEN_13472;
      end
    end else begin
      rob_payload_18_flits_fired <= _GEN_13472;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h13 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_19_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_19_tsc <= _GEN_5140;
      end
    end else begin
      rob_payload_19_tsc <= _GEN_5140;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h13 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_19_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_19_rob_idx <= _GEN_5268;
      end
    end else begin
      rob_payload_19_rob_idx <= _GEN_5268;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h13 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_19_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_19_flits_fired <= _GEN_13473;
      end
    end else begin
      rob_payload_19_flits_fired <= _GEN_13473;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h14 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_20_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_20_tsc <= _GEN_5141;
      end
    end else begin
      rob_payload_20_tsc <= _GEN_5141;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h14 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_20_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_20_rob_idx <= _GEN_5269;
      end
    end else begin
      rob_payload_20_rob_idx <= _GEN_5269;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h14 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_20_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_20_flits_fired <= _GEN_13474;
      end
    end else begin
      rob_payload_20_flits_fired <= _GEN_13474;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h15 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_21_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_21_tsc <= _GEN_5142;
      end
    end else begin
      rob_payload_21_tsc <= _GEN_5142;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h15 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_21_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_21_rob_idx <= _GEN_5270;
      end
    end else begin
      rob_payload_21_rob_idx <= _GEN_5270;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h15 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_21_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_21_flits_fired <= _GEN_13475;
      end
    end else begin
      rob_payload_21_flits_fired <= _GEN_13475;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h16 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_22_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_22_tsc <= _GEN_5143;
      end
    end else begin
      rob_payload_22_tsc <= _GEN_5143;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h16 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_22_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_22_rob_idx <= _GEN_5271;
      end
    end else begin
      rob_payload_22_rob_idx <= _GEN_5271;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h16 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_22_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_22_flits_fired <= _GEN_13476;
      end
    end else begin
      rob_payload_22_flits_fired <= _GEN_13476;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h17 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_23_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_23_tsc <= _GEN_5144;
      end
    end else begin
      rob_payload_23_tsc <= _GEN_5144;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h17 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_23_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_23_rob_idx <= _GEN_5272;
      end
    end else begin
      rob_payload_23_rob_idx <= _GEN_5272;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h17 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_23_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_23_flits_fired <= _GEN_13477;
      end
    end else begin
      rob_payload_23_flits_fired <= _GEN_13477;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h18 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_24_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_24_tsc <= _GEN_5145;
      end
    end else begin
      rob_payload_24_tsc <= _GEN_5145;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h18 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_24_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_24_rob_idx <= _GEN_5273;
      end
    end else begin
      rob_payload_24_rob_idx <= _GEN_5273;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h18 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_24_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_24_flits_fired <= _GEN_13478;
      end
    end else begin
      rob_payload_24_flits_fired <= _GEN_13478;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h19 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_25_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_25_tsc <= _GEN_5146;
      end
    end else begin
      rob_payload_25_tsc <= _GEN_5146;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h19 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_25_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_25_rob_idx <= _GEN_5274;
      end
    end else begin
      rob_payload_25_rob_idx <= _GEN_5274;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h19 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_25_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_25_flits_fired <= _GEN_13479;
      end
    end else begin
      rob_payload_25_flits_fired <= _GEN_13479;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1a == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_26_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_26_tsc <= _GEN_5147;
      end
    end else begin
      rob_payload_26_tsc <= _GEN_5147;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1a == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_26_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_26_rob_idx <= _GEN_5275;
      end
    end else begin
      rob_payload_26_rob_idx <= _GEN_5275;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h1a == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_26_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_26_flits_fired <= _GEN_13480;
      end
    end else begin
      rob_payload_26_flits_fired <= _GEN_13480;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1b == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_27_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_27_tsc <= _GEN_5148;
      end
    end else begin
      rob_payload_27_tsc <= _GEN_5148;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1b == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_27_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_27_rob_idx <= _GEN_5276;
      end
    end else begin
      rob_payload_27_rob_idx <= _GEN_5276;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h1b == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_27_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_27_flits_fired <= _GEN_13481;
      end
    end else begin
      rob_payload_27_flits_fired <= _GEN_13481;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1c == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_28_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_28_tsc <= _GEN_5149;
      end
    end else begin
      rob_payload_28_tsc <= _GEN_5149;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1c == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_28_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_28_rob_idx <= _GEN_5277;
      end
    end else begin
      rob_payload_28_rob_idx <= _GEN_5277;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h1c == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_28_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_28_flits_fired <= _GEN_13482;
      end
    end else begin
      rob_payload_28_flits_fired <= _GEN_13482;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1d == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_29_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_29_tsc <= _GEN_5150;
      end
    end else begin
      rob_payload_29_tsc <= _GEN_5150;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1d == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_29_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_29_rob_idx <= _GEN_5278;
      end
    end else begin
      rob_payload_29_rob_idx <= _GEN_5278;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h1d == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_29_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_29_flits_fired <= _GEN_13483;
      end
    end else begin
      rob_payload_29_flits_fired <= _GEN_13483;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1e == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_30_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_30_tsc <= _GEN_5151;
      end
    end else begin
      rob_payload_30_tsc <= _GEN_5151;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1e == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_30_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_30_rob_idx <= _GEN_5279;
      end
    end else begin
      rob_payload_30_rob_idx <= _GEN_5279;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h1e == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_30_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_30_flits_fired <= _GEN_13484;
      end
    end else begin
      rob_payload_30_flits_fired <= _GEN_13484;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1f == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_31_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_31_tsc <= _GEN_5152;
      end
    end else begin
      rob_payload_31_tsc <= _GEN_5152;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1f == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_31_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_31_rob_idx <= _GEN_5280;
      end
    end else begin
      rob_payload_31_rob_idx <= _GEN_5280;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h1f == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_31_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_31_flits_fired <= _GEN_13485;
      end
    end else begin
      rob_payload_31_flits_fired <= _GEN_13485;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h20 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_32_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_32_tsc <= _GEN_5153;
      end
    end else begin
      rob_payload_32_tsc <= _GEN_5153;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h20 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_32_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_32_rob_idx <= _GEN_5281;
      end
    end else begin
      rob_payload_32_rob_idx <= _GEN_5281;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h20 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_32_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_32_flits_fired <= _GEN_13486;
      end
    end else begin
      rob_payload_32_flits_fired <= _GEN_13486;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h21 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_33_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_33_tsc <= _GEN_5154;
      end
    end else begin
      rob_payload_33_tsc <= _GEN_5154;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h21 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_33_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_33_rob_idx <= _GEN_5282;
      end
    end else begin
      rob_payload_33_rob_idx <= _GEN_5282;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h21 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_33_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_33_flits_fired <= _GEN_13487;
      end
    end else begin
      rob_payload_33_flits_fired <= _GEN_13487;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h22 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_34_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_34_tsc <= _GEN_5155;
      end
    end else begin
      rob_payload_34_tsc <= _GEN_5155;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h22 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_34_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_34_rob_idx <= _GEN_5283;
      end
    end else begin
      rob_payload_34_rob_idx <= _GEN_5283;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h22 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_34_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_34_flits_fired <= _GEN_13488;
      end
    end else begin
      rob_payload_34_flits_fired <= _GEN_13488;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h23 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_35_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_35_tsc <= _GEN_5156;
      end
    end else begin
      rob_payload_35_tsc <= _GEN_5156;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h23 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_35_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_35_rob_idx <= _GEN_5284;
      end
    end else begin
      rob_payload_35_rob_idx <= _GEN_5284;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h23 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_35_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_35_flits_fired <= _GEN_13489;
      end
    end else begin
      rob_payload_35_flits_fired <= _GEN_13489;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h24 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_36_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_36_tsc <= _GEN_5157;
      end
    end else begin
      rob_payload_36_tsc <= _GEN_5157;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h24 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_36_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_36_rob_idx <= _GEN_5285;
      end
    end else begin
      rob_payload_36_rob_idx <= _GEN_5285;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h24 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_36_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_36_flits_fired <= _GEN_13490;
      end
    end else begin
      rob_payload_36_flits_fired <= _GEN_13490;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h25 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_37_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_37_tsc <= _GEN_5158;
      end
    end else begin
      rob_payload_37_tsc <= _GEN_5158;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h25 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_37_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_37_rob_idx <= _GEN_5286;
      end
    end else begin
      rob_payload_37_rob_idx <= _GEN_5286;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h25 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_37_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_37_flits_fired <= _GEN_13491;
      end
    end else begin
      rob_payload_37_flits_fired <= _GEN_13491;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h26 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_38_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_38_tsc <= _GEN_5159;
      end
    end else begin
      rob_payload_38_tsc <= _GEN_5159;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h26 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_38_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_38_rob_idx <= _GEN_5287;
      end
    end else begin
      rob_payload_38_rob_idx <= _GEN_5287;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h26 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_38_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_38_flits_fired <= _GEN_13492;
      end
    end else begin
      rob_payload_38_flits_fired <= _GEN_13492;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h27 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_39_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_39_tsc <= _GEN_5160;
      end
    end else begin
      rob_payload_39_tsc <= _GEN_5160;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h27 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_39_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_39_rob_idx <= _GEN_5288;
      end
    end else begin
      rob_payload_39_rob_idx <= _GEN_5288;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h27 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_39_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_39_flits_fired <= _GEN_13493;
      end
    end else begin
      rob_payload_39_flits_fired <= _GEN_13493;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h28 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_40_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_40_tsc <= _GEN_5161;
      end
    end else begin
      rob_payload_40_tsc <= _GEN_5161;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h28 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_40_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_40_rob_idx <= _GEN_5289;
      end
    end else begin
      rob_payload_40_rob_idx <= _GEN_5289;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h28 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_40_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_40_flits_fired <= _GEN_13494;
      end
    end else begin
      rob_payload_40_flits_fired <= _GEN_13494;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h29 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_41_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_41_tsc <= _GEN_5162;
      end
    end else begin
      rob_payload_41_tsc <= _GEN_5162;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h29 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_41_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_41_rob_idx <= _GEN_5290;
      end
    end else begin
      rob_payload_41_rob_idx <= _GEN_5290;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h29 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_41_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_41_flits_fired <= _GEN_13495;
      end
    end else begin
      rob_payload_41_flits_fired <= _GEN_13495;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2a == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_42_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_42_tsc <= _GEN_5163;
      end
    end else begin
      rob_payload_42_tsc <= _GEN_5163;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2a == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_42_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_42_rob_idx <= _GEN_5291;
      end
    end else begin
      rob_payload_42_rob_idx <= _GEN_5291;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h2a == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_42_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_42_flits_fired <= _GEN_13496;
      end
    end else begin
      rob_payload_42_flits_fired <= _GEN_13496;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2b == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_43_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_43_tsc <= _GEN_5164;
      end
    end else begin
      rob_payload_43_tsc <= _GEN_5164;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2b == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_43_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_43_rob_idx <= _GEN_5292;
      end
    end else begin
      rob_payload_43_rob_idx <= _GEN_5292;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h2b == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_43_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_43_flits_fired <= _GEN_13497;
      end
    end else begin
      rob_payload_43_flits_fired <= _GEN_13497;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2c == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_44_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_44_tsc <= _GEN_5165;
      end
    end else begin
      rob_payload_44_tsc <= _GEN_5165;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2c == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_44_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_44_rob_idx <= _GEN_5293;
      end
    end else begin
      rob_payload_44_rob_idx <= _GEN_5293;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h2c == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_44_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_44_flits_fired <= _GEN_13498;
      end
    end else begin
      rob_payload_44_flits_fired <= _GEN_13498;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2d == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_45_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_45_tsc <= _GEN_5166;
      end
    end else begin
      rob_payload_45_tsc <= _GEN_5166;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2d == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_45_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_45_rob_idx <= _GEN_5294;
      end
    end else begin
      rob_payload_45_rob_idx <= _GEN_5294;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h2d == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_45_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_45_flits_fired <= _GEN_13499;
      end
    end else begin
      rob_payload_45_flits_fired <= _GEN_13499;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2e == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_46_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_46_tsc <= _GEN_5167;
      end
    end else begin
      rob_payload_46_tsc <= _GEN_5167;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2e == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_46_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_46_rob_idx <= _GEN_5295;
      end
    end else begin
      rob_payload_46_rob_idx <= _GEN_5295;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h2e == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_46_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_46_flits_fired <= _GEN_13500;
      end
    end else begin
      rob_payload_46_flits_fired <= _GEN_13500;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2f == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_47_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_47_tsc <= _GEN_5168;
      end
    end else begin
      rob_payload_47_tsc <= _GEN_5168;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2f == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_47_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_47_rob_idx <= _GEN_5296;
      end
    end else begin
      rob_payload_47_rob_idx <= _GEN_5296;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h2f == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_47_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_47_flits_fired <= _GEN_13501;
      end
    end else begin
      rob_payload_47_flits_fired <= _GEN_13501;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h30 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_48_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_48_tsc <= _GEN_5169;
      end
    end else begin
      rob_payload_48_tsc <= _GEN_5169;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h30 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_48_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_48_rob_idx <= _GEN_5297;
      end
    end else begin
      rob_payload_48_rob_idx <= _GEN_5297;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h30 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_48_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_48_flits_fired <= _GEN_13502;
      end
    end else begin
      rob_payload_48_flits_fired <= _GEN_13502;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h31 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_49_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_49_tsc <= _GEN_5170;
      end
    end else begin
      rob_payload_49_tsc <= _GEN_5170;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h31 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_49_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_49_rob_idx <= _GEN_5298;
      end
    end else begin
      rob_payload_49_rob_idx <= _GEN_5298;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h31 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_49_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_49_flits_fired <= _GEN_13503;
      end
    end else begin
      rob_payload_49_flits_fired <= _GEN_13503;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h32 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_50_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_50_tsc <= _GEN_5171;
      end
    end else begin
      rob_payload_50_tsc <= _GEN_5171;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h32 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_50_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_50_rob_idx <= _GEN_5299;
      end
    end else begin
      rob_payload_50_rob_idx <= _GEN_5299;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h32 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_50_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_50_flits_fired <= _GEN_13504;
      end
    end else begin
      rob_payload_50_flits_fired <= _GEN_13504;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h33 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_51_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_51_tsc <= _GEN_5172;
      end
    end else begin
      rob_payload_51_tsc <= _GEN_5172;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h33 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_51_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_51_rob_idx <= _GEN_5300;
      end
    end else begin
      rob_payload_51_rob_idx <= _GEN_5300;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h33 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_51_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_51_flits_fired <= _GEN_13505;
      end
    end else begin
      rob_payload_51_flits_fired <= _GEN_13505;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h34 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_52_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_52_tsc <= _GEN_5173;
      end
    end else begin
      rob_payload_52_tsc <= _GEN_5173;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h34 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_52_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_52_rob_idx <= _GEN_5301;
      end
    end else begin
      rob_payload_52_rob_idx <= _GEN_5301;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h34 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_52_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_52_flits_fired <= _GEN_13506;
      end
    end else begin
      rob_payload_52_flits_fired <= _GEN_13506;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h35 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_53_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_53_tsc <= _GEN_5174;
      end
    end else begin
      rob_payload_53_tsc <= _GEN_5174;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h35 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_53_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_53_rob_idx <= _GEN_5302;
      end
    end else begin
      rob_payload_53_rob_idx <= _GEN_5302;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h35 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_53_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_53_flits_fired <= _GEN_13507;
      end
    end else begin
      rob_payload_53_flits_fired <= _GEN_13507;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h36 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_54_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_54_tsc <= _GEN_5175;
      end
    end else begin
      rob_payload_54_tsc <= _GEN_5175;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h36 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_54_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_54_rob_idx <= _GEN_5303;
      end
    end else begin
      rob_payload_54_rob_idx <= _GEN_5303;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h36 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_54_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_54_flits_fired <= _GEN_13508;
      end
    end else begin
      rob_payload_54_flits_fired <= _GEN_13508;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h37 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_55_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_55_tsc <= _GEN_5176;
      end
    end else begin
      rob_payload_55_tsc <= _GEN_5176;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h37 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_55_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_55_rob_idx <= _GEN_5304;
      end
    end else begin
      rob_payload_55_rob_idx <= _GEN_5304;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h37 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_55_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_55_flits_fired <= _GEN_13509;
      end
    end else begin
      rob_payload_55_flits_fired <= _GEN_13509;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h38 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_56_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_56_tsc <= _GEN_5177;
      end
    end else begin
      rob_payload_56_tsc <= _GEN_5177;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h38 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_56_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_56_rob_idx <= _GEN_5305;
      end
    end else begin
      rob_payload_56_rob_idx <= _GEN_5305;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h38 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_56_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_56_flits_fired <= _GEN_13510;
      end
    end else begin
      rob_payload_56_flits_fired <= _GEN_13510;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h39 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_57_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_57_tsc <= _GEN_5178;
      end
    end else begin
      rob_payload_57_tsc <= _GEN_5178;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h39 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_57_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_57_rob_idx <= _GEN_5306;
      end
    end else begin
      rob_payload_57_rob_idx <= _GEN_5306;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h39 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_57_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_57_flits_fired <= _GEN_13511;
      end
    end else begin
      rob_payload_57_flits_fired <= _GEN_13511;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3a == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_58_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_58_tsc <= _GEN_5179;
      end
    end else begin
      rob_payload_58_tsc <= _GEN_5179;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3a == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_58_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_58_rob_idx <= _GEN_5307;
      end
    end else begin
      rob_payload_58_rob_idx <= _GEN_5307;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h3a == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_58_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_58_flits_fired <= _GEN_13512;
      end
    end else begin
      rob_payload_58_flits_fired <= _GEN_13512;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3b == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_59_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_59_tsc <= _GEN_5180;
      end
    end else begin
      rob_payload_59_tsc <= _GEN_5180;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3b == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_59_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_59_rob_idx <= _GEN_5308;
      end
    end else begin
      rob_payload_59_rob_idx <= _GEN_5308;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h3b == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_59_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_59_flits_fired <= _GEN_13513;
      end
    end else begin
      rob_payload_59_flits_fired <= _GEN_13513;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3c == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_60_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_60_tsc <= _GEN_5181;
      end
    end else begin
      rob_payload_60_tsc <= _GEN_5181;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3c == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_60_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_60_rob_idx <= _GEN_5309;
      end
    end else begin
      rob_payload_60_rob_idx <= _GEN_5309;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h3c == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_60_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_60_flits_fired <= _GEN_13514;
      end
    end else begin
      rob_payload_60_flits_fired <= _GEN_13514;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3d == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_61_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_61_tsc <= _GEN_5182;
      end
    end else begin
      rob_payload_61_tsc <= _GEN_5182;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3d == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_61_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_61_rob_idx <= _GEN_5310;
      end
    end else begin
      rob_payload_61_rob_idx <= _GEN_5310;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h3d == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_61_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_61_flits_fired <= _GEN_13515;
      end
    end else begin
      rob_payload_61_flits_fired <= _GEN_13515;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3e == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_62_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_62_tsc <= _GEN_5183;
      end
    end else begin
      rob_payload_62_tsc <= _GEN_5183;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3e == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_62_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_62_rob_idx <= _GEN_5311;
      end
    end else begin
      rob_payload_62_rob_idx <= _GEN_5311;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h3e == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_62_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_62_flits_fired <= _GEN_13516;
      end
    end else begin
      rob_payload_62_flits_fired <= _GEN_13516;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3f == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_63_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_63_tsc <= _GEN_5184;
      end
    end else begin
      rob_payload_63_tsc <= _GEN_5184;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3f == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_63_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_63_rob_idx <= _GEN_5312;
      end
    end else begin
      rob_payload_63_rob_idx <= _GEN_5312;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h3f == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_63_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_63_flits_fired <= _GEN_13517;
      end
    end else begin
      rob_payload_63_flits_fired <= _GEN_13517;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h40 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_64_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_64_tsc <= _GEN_5185;
      end
    end else begin
      rob_payload_64_tsc <= _GEN_5185;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h40 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_64_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_64_rob_idx <= _GEN_5313;
      end
    end else begin
      rob_payload_64_rob_idx <= _GEN_5313;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h40 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_64_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_64_flits_fired <= _GEN_13518;
      end
    end else begin
      rob_payload_64_flits_fired <= _GEN_13518;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h41 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_65_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_65_tsc <= _GEN_5186;
      end
    end else begin
      rob_payload_65_tsc <= _GEN_5186;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h41 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_65_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_65_rob_idx <= _GEN_5314;
      end
    end else begin
      rob_payload_65_rob_idx <= _GEN_5314;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h41 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_65_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_65_flits_fired <= _GEN_13519;
      end
    end else begin
      rob_payload_65_flits_fired <= _GEN_13519;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h42 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_66_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_66_tsc <= _GEN_5187;
      end
    end else begin
      rob_payload_66_tsc <= _GEN_5187;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h42 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_66_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_66_rob_idx <= _GEN_5315;
      end
    end else begin
      rob_payload_66_rob_idx <= _GEN_5315;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h42 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_66_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_66_flits_fired <= _GEN_13520;
      end
    end else begin
      rob_payload_66_flits_fired <= _GEN_13520;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h43 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_67_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_67_tsc <= _GEN_5188;
      end
    end else begin
      rob_payload_67_tsc <= _GEN_5188;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h43 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_67_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_67_rob_idx <= _GEN_5316;
      end
    end else begin
      rob_payload_67_rob_idx <= _GEN_5316;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h43 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_67_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_67_flits_fired <= _GEN_13521;
      end
    end else begin
      rob_payload_67_flits_fired <= _GEN_13521;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h44 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_68_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_68_tsc <= _GEN_5189;
      end
    end else begin
      rob_payload_68_tsc <= _GEN_5189;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h44 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_68_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_68_rob_idx <= _GEN_5317;
      end
    end else begin
      rob_payload_68_rob_idx <= _GEN_5317;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h44 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_68_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_68_flits_fired <= _GEN_13522;
      end
    end else begin
      rob_payload_68_flits_fired <= _GEN_13522;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h45 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_69_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_69_tsc <= _GEN_5190;
      end
    end else begin
      rob_payload_69_tsc <= _GEN_5190;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h45 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_69_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_69_rob_idx <= _GEN_5318;
      end
    end else begin
      rob_payload_69_rob_idx <= _GEN_5318;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h45 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_69_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_69_flits_fired <= _GEN_13523;
      end
    end else begin
      rob_payload_69_flits_fired <= _GEN_13523;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h46 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_70_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_70_tsc <= _GEN_5191;
      end
    end else begin
      rob_payload_70_tsc <= _GEN_5191;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h46 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_70_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_70_rob_idx <= _GEN_5319;
      end
    end else begin
      rob_payload_70_rob_idx <= _GEN_5319;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h46 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_70_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_70_flits_fired <= _GEN_13524;
      end
    end else begin
      rob_payload_70_flits_fired <= _GEN_13524;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h47 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_71_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_71_tsc <= _GEN_5192;
      end
    end else begin
      rob_payload_71_tsc <= _GEN_5192;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h47 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_71_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_71_rob_idx <= _GEN_5320;
      end
    end else begin
      rob_payload_71_rob_idx <= _GEN_5320;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h47 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_71_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_71_flits_fired <= _GEN_13525;
      end
    end else begin
      rob_payload_71_flits_fired <= _GEN_13525;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h48 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_72_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_72_tsc <= _GEN_5193;
      end
    end else begin
      rob_payload_72_tsc <= _GEN_5193;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h48 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_72_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_72_rob_idx <= _GEN_5321;
      end
    end else begin
      rob_payload_72_rob_idx <= _GEN_5321;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h48 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_72_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_72_flits_fired <= _GEN_13526;
      end
    end else begin
      rob_payload_72_flits_fired <= _GEN_13526;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h49 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_73_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_73_tsc <= _GEN_5194;
      end
    end else begin
      rob_payload_73_tsc <= _GEN_5194;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h49 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_73_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_73_rob_idx <= _GEN_5322;
      end
    end else begin
      rob_payload_73_rob_idx <= _GEN_5322;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h49 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_73_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_73_flits_fired <= _GEN_13527;
      end
    end else begin
      rob_payload_73_flits_fired <= _GEN_13527;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4a == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_74_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_74_tsc <= _GEN_5195;
      end
    end else begin
      rob_payload_74_tsc <= _GEN_5195;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4a == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_74_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_74_rob_idx <= _GEN_5323;
      end
    end else begin
      rob_payload_74_rob_idx <= _GEN_5323;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h4a == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_74_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_74_flits_fired <= _GEN_13528;
      end
    end else begin
      rob_payload_74_flits_fired <= _GEN_13528;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4b == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_75_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_75_tsc <= _GEN_5196;
      end
    end else begin
      rob_payload_75_tsc <= _GEN_5196;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4b == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_75_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_75_rob_idx <= _GEN_5324;
      end
    end else begin
      rob_payload_75_rob_idx <= _GEN_5324;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h4b == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_75_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_75_flits_fired <= _GEN_13529;
      end
    end else begin
      rob_payload_75_flits_fired <= _GEN_13529;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4c == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_76_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_76_tsc <= _GEN_5197;
      end
    end else begin
      rob_payload_76_tsc <= _GEN_5197;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4c == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_76_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_76_rob_idx <= _GEN_5325;
      end
    end else begin
      rob_payload_76_rob_idx <= _GEN_5325;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h4c == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_76_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_76_flits_fired <= _GEN_13530;
      end
    end else begin
      rob_payload_76_flits_fired <= _GEN_13530;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4d == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_77_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_77_tsc <= _GEN_5198;
      end
    end else begin
      rob_payload_77_tsc <= _GEN_5198;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4d == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_77_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_77_rob_idx <= _GEN_5326;
      end
    end else begin
      rob_payload_77_rob_idx <= _GEN_5326;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h4d == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_77_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_77_flits_fired <= _GEN_13531;
      end
    end else begin
      rob_payload_77_flits_fired <= _GEN_13531;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4e == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_78_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_78_tsc <= _GEN_5199;
      end
    end else begin
      rob_payload_78_tsc <= _GEN_5199;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4e == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_78_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_78_rob_idx <= _GEN_5327;
      end
    end else begin
      rob_payload_78_rob_idx <= _GEN_5327;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h4e == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_78_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_78_flits_fired <= _GEN_13532;
      end
    end else begin
      rob_payload_78_flits_fired <= _GEN_13532;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4f == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_79_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_79_tsc <= _GEN_5200;
      end
    end else begin
      rob_payload_79_tsc <= _GEN_5200;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4f == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_79_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_79_rob_idx <= _GEN_5328;
      end
    end else begin
      rob_payload_79_rob_idx <= _GEN_5328;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h4f == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_79_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_79_flits_fired <= _GEN_13533;
      end
    end else begin
      rob_payload_79_flits_fired <= _GEN_13533;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h50 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_80_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_80_tsc <= _GEN_5201;
      end
    end else begin
      rob_payload_80_tsc <= _GEN_5201;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h50 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_80_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_80_rob_idx <= _GEN_5329;
      end
    end else begin
      rob_payload_80_rob_idx <= _GEN_5329;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h50 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_80_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_80_flits_fired <= _GEN_13534;
      end
    end else begin
      rob_payload_80_flits_fired <= _GEN_13534;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h51 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_81_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_81_tsc <= _GEN_5202;
      end
    end else begin
      rob_payload_81_tsc <= _GEN_5202;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h51 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_81_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_81_rob_idx <= _GEN_5330;
      end
    end else begin
      rob_payload_81_rob_idx <= _GEN_5330;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h51 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_81_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_81_flits_fired <= _GEN_13535;
      end
    end else begin
      rob_payload_81_flits_fired <= _GEN_13535;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h52 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_82_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_82_tsc <= _GEN_5203;
      end
    end else begin
      rob_payload_82_tsc <= _GEN_5203;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h52 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_82_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_82_rob_idx <= _GEN_5331;
      end
    end else begin
      rob_payload_82_rob_idx <= _GEN_5331;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h52 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_82_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_82_flits_fired <= _GEN_13536;
      end
    end else begin
      rob_payload_82_flits_fired <= _GEN_13536;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h53 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_83_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_83_tsc <= _GEN_5204;
      end
    end else begin
      rob_payload_83_tsc <= _GEN_5204;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h53 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_83_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_83_rob_idx <= _GEN_5332;
      end
    end else begin
      rob_payload_83_rob_idx <= _GEN_5332;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h53 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_83_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_83_flits_fired <= _GEN_13537;
      end
    end else begin
      rob_payload_83_flits_fired <= _GEN_13537;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h54 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_84_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_84_tsc <= _GEN_5205;
      end
    end else begin
      rob_payload_84_tsc <= _GEN_5205;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h54 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_84_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_84_rob_idx <= _GEN_5333;
      end
    end else begin
      rob_payload_84_rob_idx <= _GEN_5333;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h54 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_84_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_84_flits_fired <= _GEN_13538;
      end
    end else begin
      rob_payload_84_flits_fired <= _GEN_13538;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h55 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_85_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_85_tsc <= _GEN_5206;
      end
    end else begin
      rob_payload_85_tsc <= _GEN_5206;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h55 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_85_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_85_rob_idx <= _GEN_5334;
      end
    end else begin
      rob_payload_85_rob_idx <= _GEN_5334;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h55 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_85_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_85_flits_fired <= _GEN_13539;
      end
    end else begin
      rob_payload_85_flits_fired <= _GEN_13539;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h56 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_86_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_86_tsc <= _GEN_5207;
      end
    end else begin
      rob_payload_86_tsc <= _GEN_5207;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h56 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_86_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_86_rob_idx <= _GEN_5335;
      end
    end else begin
      rob_payload_86_rob_idx <= _GEN_5335;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h56 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_86_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_86_flits_fired <= _GEN_13540;
      end
    end else begin
      rob_payload_86_flits_fired <= _GEN_13540;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h57 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_87_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_87_tsc <= _GEN_5208;
      end
    end else begin
      rob_payload_87_tsc <= _GEN_5208;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h57 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_87_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_87_rob_idx <= _GEN_5336;
      end
    end else begin
      rob_payload_87_rob_idx <= _GEN_5336;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h57 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_87_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_87_flits_fired <= _GEN_13541;
      end
    end else begin
      rob_payload_87_flits_fired <= _GEN_13541;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h58 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_88_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_88_tsc <= _GEN_5209;
      end
    end else begin
      rob_payload_88_tsc <= _GEN_5209;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h58 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_88_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_88_rob_idx <= _GEN_5337;
      end
    end else begin
      rob_payload_88_rob_idx <= _GEN_5337;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h58 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_88_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_88_flits_fired <= _GEN_13542;
      end
    end else begin
      rob_payload_88_flits_fired <= _GEN_13542;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h59 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_89_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_89_tsc <= _GEN_5210;
      end
    end else begin
      rob_payload_89_tsc <= _GEN_5210;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h59 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_89_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_89_rob_idx <= _GEN_5338;
      end
    end else begin
      rob_payload_89_rob_idx <= _GEN_5338;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h59 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_89_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_89_flits_fired <= _GEN_13543;
      end
    end else begin
      rob_payload_89_flits_fired <= _GEN_13543;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5a == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_90_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_90_tsc <= _GEN_5211;
      end
    end else begin
      rob_payload_90_tsc <= _GEN_5211;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5a == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_90_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_90_rob_idx <= _GEN_5339;
      end
    end else begin
      rob_payload_90_rob_idx <= _GEN_5339;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h5a == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_90_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_90_flits_fired <= _GEN_13544;
      end
    end else begin
      rob_payload_90_flits_fired <= _GEN_13544;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5b == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_91_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_91_tsc <= _GEN_5212;
      end
    end else begin
      rob_payload_91_tsc <= _GEN_5212;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5b == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_91_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_91_rob_idx <= _GEN_5340;
      end
    end else begin
      rob_payload_91_rob_idx <= _GEN_5340;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h5b == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_91_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_91_flits_fired <= _GEN_13545;
      end
    end else begin
      rob_payload_91_flits_fired <= _GEN_13545;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5c == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_92_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_92_tsc <= _GEN_5213;
      end
    end else begin
      rob_payload_92_tsc <= _GEN_5213;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5c == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_92_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_92_rob_idx <= _GEN_5341;
      end
    end else begin
      rob_payload_92_rob_idx <= _GEN_5341;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h5c == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_92_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_92_flits_fired <= _GEN_13546;
      end
    end else begin
      rob_payload_92_flits_fired <= _GEN_13546;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5d == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_93_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_93_tsc <= _GEN_5214;
      end
    end else begin
      rob_payload_93_tsc <= _GEN_5214;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5d == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_93_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_93_rob_idx <= _GEN_5342;
      end
    end else begin
      rob_payload_93_rob_idx <= _GEN_5342;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h5d == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_93_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_93_flits_fired <= _GEN_13547;
      end
    end else begin
      rob_payload_93_flits_fired <= _GEN_13547;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5e == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_94_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_94_tsc <= _GEN_5215;
      end
    end else begin
      rob_payload_94_tsc <= _GEN_5215;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5e == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_94_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_94_rob_idx <= _GEN_5343;
      end
    end else begin
      rob_payload_94_rob_idx <= _GEN_5343;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h5e == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_94_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_94_flits_fired <= _GEN_13548;
      end
    end else begin
      rob_payload_94_flits_fired <= _GEN_13548;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5f == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_95_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_95_tsc <= _GEN_5216;
      end
    end else begin
      rob_payload_95_tsc <= _GEN_5216;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5f == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_95_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_95_rob_idx <= _GEN_5344;
      end
    end else begin
      rob_payload_95_rob_idx <= _GEN_5344;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h5f == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_95_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_95_flits_fired <= _GEN_13549;
      end
    end else begin
      rob_payload_95_flits_fired <= _GEN_13549;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h60 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_96_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_96_tsc <= _GEN_5217;
      end
    end else begin
      rob_payload_96_tsc <= _GEN_5217;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h60 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_96_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_96_rob_idx <= _GEN_5345;
      end
    end else begin
      rob_payload_96_rob_idx <= _GEN_5345;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h60 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_96_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_96_flits_fired <= _GEN_13550;
      end
    end else begin
      rob_payload_96_flits_fired <= _GEN_13550;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h61 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_97_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_97_tsc <= _GEN_5218;
      end
    end else begin
      rob_payload_97_tsc <= _GEN_5218;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h61 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_97_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_97_rob_idx <= _GEN_5346;
      end
    end else begin
      rob_payload_97_rob_idx <= _GEN_5346;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h61 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_97_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_97_flits_fired <= _GEN_13551;
      end
    end else begin
      rob_payload_97_flits_fired <= _GEN_13551;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h62 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_98_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_98_tsc <= _GEN_5219;
      end
    end else begin
      rob_payload_98_tsc <= _GEN_5219;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h62 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_98_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_98_rob_idx <= _GEN_5347;
      end
    end else begin
      rob_payload_98_rob_idx <= _GEN_5347;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h62 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_98_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_98_flits_fired <= _GEN_13552;
      end
    end else begin
      rob_payload_98_flits_fired <= _GEN_13552;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h63 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_99_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_99_tsc <= _GEN_5220;
      end
    end else begin
      rob_payload_99_tsc <= _GEN_5220;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h63 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_99_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_99_rob_idx <= _GEN_5348;
      end
    end else begin
      rob_payload_99_rob_idx <= _GEN_5348;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h63 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_99_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_99_flits_fired <= _GEN_13553;
      end
    end else begin
      rob_payload_99_flits_fired <= _GEN_13553;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h64 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_100_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_100_tsc <= _GEN_5221;
      end
    end else begin
      rob_payload_100_tsc <= _GEN_5221;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h64 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_100_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_100_rob_idx <= _GEN_5349;
      end
    end else begin
      rob_payload_100_rob_idx <= _GEN_5349;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h64 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_100_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_100_flits_fired <= _GEN_13554;
      end
    end else begin
      rob_payload_100_flits_fired <= _GEN_13554;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h65 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_101_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_101_tsc <= _GEN_5222;
      end
    end else begin
      rob_payload_101_tsc <= _GEN_5222;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h65 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_101_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_101_rob_idx <= _GEN_5350;
      end
    end else begin
      rob_payload_101_rob_idx <= _GEN_5350;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h65 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_101_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_101_flits_fired <= _GEN_13555;
      end
    end else begin
      rob_payload_101_flits_fired <= _GEN_13555;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h66 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_102_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_102_tsc <= _GEN_5223;
      end
    end else begin
      rob_payload_102_tsc <= _GEN_5223;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h66 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_102_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_102_rob_idx <= _GEN_5351;
      end
    end else begin
      rob_payload_102_rob_idx <= _GEN_5351;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h66 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_102_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_102_flits_fired <= _GEN_13556;
      end
    end else begin
      rob_payload_102_flits_fired <= _GEN_13556;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h67 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_103_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_103_tsc <= _GEN_5224;
      end
    end else begin
      rob_payload_103_tsc <= _GEN_5224;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h67 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_103_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_103_rob_idx <= _GEN_5352;
      end
    end else begin
      rob_payload_103_rob_idx <= _GEN_5352;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h67 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_103_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_103_flits_fired <= _GEN_13557;
      end
    end else begin
      rob_payload_103_flits_fired <= _GEN_13557;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h68 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_104_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_104_tsc <= _GEN_5225;
      end
    end else begin
      rob_payload_104_tsc <= _GEN_5225;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h68 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_104_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_104_rob_idx <= _GEN_5353;
      end
    end else begin
      rob_payload_104_rob_idx <= _GEN_5353;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h68 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_104_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_104_flits_fired <= _GEN_13558;
      end
    end else begin
      rob_payload_104_flits_fired <= _GEN_13558;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h69 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_105_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_105_tsc <= _GEN_5226;
      end
    end else begin
      rob_payload_105_tsc <= _GEN_5226;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h69 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_105_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_105_rob_idx <= _GEN_5354;
      end
    end else begin
      rob_payload_105_rob_idx <= _GEN_5354;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h69 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_105_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_105_flits_fired <= _GEN_13559;
      end
    end else begin
      rob_payload_105_flits_fired <= _GEN_13559;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6a == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_106_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_106_tsc <= _GEN_5227;
      end
    end else begin
      rob_payload_106_tsc <= _GEN_5227;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6a == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_106_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_106_rob_idx <= _GEN_5355;
      end
    end else begin
      rob_payload_106_rob_idx <= _GEN_5355;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h6a == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_106_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_106_flits_fired <= _GEN_13560;
      end
    end else begin
      rob_payload_106_flits_fired <= _GEN_13560;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6b == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_107_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_107_tsc <= _GEN_5228;
      end
    end else begin
      rob_payload_107_tsc <= _GEN_5228;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6b == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_107_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_107_rob_idx <= _GEN_5356;
      end
    end else begin
      rob_payload_107_rob_idx <= _GEN_5356;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h6b == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_107_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_107_flits_fired <= _GEN_13561;
      end
    end else begin
      rob_payload_107_flits_fired <= _GEN_13561;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6c == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_108_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_108_tsc <= _GEN_5229;
      end
    end else begin
      rob_payload_108_tsc <= _GEN_5229;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6c == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_108_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_108_rob_idx <= _GEN_5357;
      end
    end else begin
      rob_payload_108_rob_idx <= _GEN_5357;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h6c == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_108_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_108_flits_fired <= _GEN_13562;
      end
    end else begin
      rob_payload_108_flits_fired <= _GEN_13562;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6d == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_109_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_109_tsc <= _GEN_5230;
      end
    end else begin
      rob_payload_109_tsc <= _GEN_5230;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6d == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_109_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_109_rob_idx <= _GEN_5358;
      end
    end else begin
      rob_payload_109_rob_idx <= _GEN_5358;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h6d == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_109_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_109_flits_fired <= _GEN_13563;
      end
    end else begin
      rob_payload_109_flits_fired <= _GEN_13563;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6e == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_110_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_110_tsc <= _GEN_5231;
      end
    end else begin
      rob_payload_110_tsc <= _GEN_5231;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6e == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_110_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_110_rob_idx <= _GEN_5359;
      end
    end else begin
      rob_payload_110_rob_idx <= _GEN_5359;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h6e == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_110_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_110_flits_fired <= _GEN_13564;
      end
    end else begin
      rob_payload_110_flits_fired <= _GEN_13564;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6f == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_111_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_111_tsc <= _GEN_5232;
      end
    end else begin
      rob_payload_111_tsc <= _GEN_5232;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6f == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_111_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_111_rob_idx <= _GEN_5360;
      end
    end else begin
      rob_payload_111_rob_idx <= _GEN_5360;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h6f == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_111_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_111_flits_fired <= _GEN_13565;
      end
    end else begin
      rob_payload_111_flits_fired <= _GEN_13565;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h70 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_112_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_112_tsc <= _GEN_5233;
      end
    end else begin
      rob_payload_112_tsc <= _GEN_5233;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h70 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_112_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_112_rob_idx <= _GEN_5361;
      end
    end else begin
      rob_payload_112_rob_idx <= _GEN_5361;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h70 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_112_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_112_flits_fired <= _GEN_13566;
      end
    end else begin
      rob_payload_112_flits_fired <= _GEN_13566;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h71 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_113_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_113_tsc <= _GEN_5234;
      end
    end else begin
      rob_payload_113_tsc <= _GEN_5234;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h71 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_113_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_113_rob_idx <= _GEN_5362;
      end
    end else begin
      rob_payload_113_rob_idx <= _GEN_5362;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h71 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_113_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_113_flits_fired <= _GEN_13567;
      end
    end else begin
      rob_payload_113_flits_fired <= _GEN_13567;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h72 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_114_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_114_tsc <= _GEN_5235;
      end
    end else begin
      rob_payload_114_tsc <= _GEN_5235;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h72 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_114_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_114_rob_idx <= _GEN_5363;
      end
    end else begin
      rob_payload_114_rob_idx <= _GEN_5363;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h72 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_114_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_114_flits_fired <= _GEN_13568;
      end
    end else begin
      rob_payload_114_flits_fired <= _GEN_13568;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h73 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_115_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_115_tsc <= _GEN_5236;
      end
    end else begin
      rob_payload_115_tsc <= _GEN_5236;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h73 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_115_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_115_rob_idx <= _GEN_5364;
      end
    end else begin
      rob_payload_115_rob_idx <= _GEN_5364;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h73 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_115_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_115_flits_fired <= _GEN_13569;
      end
    end else begin
      rob_payload_115_flits_fired <= _GEN_13569;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h74 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_116_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_116_tsc <= _GEN_5237;
      end
    end else begin
      rob_payload_116_tsc <= _GEN_5237;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h74 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_116_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_116_rob_idx <= _GEN_5365;
      end
    end else begin
      rob_payload_116_rob_idx <= _GEN_5365;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h74 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_116_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_116_flits_fired <= _GEN_13570;
      end
    end else begin
      rob_payload_116_flits_fired <= _GEN_13570;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h75 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_117_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_117_tsc <= _GEN_5238;
      end
    end else begin
      rob_payload_117_tsc <= _GEN_5238;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h75 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_117_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_117_rob_idx <= _GEN_5366;
      end
    end else begin
      rob_payload_117_rob_idx <= _GEN_5366;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h75 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_117_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_117_flits_fired <= _GEN_13571;
      end
    end else begin
      rob_payload_117_flits_fired <= _GEN_13571;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h76 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_118_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_118_tsc <= _GEN_5239;
      end
    end else begin
      rob_payload_118_tsc <= _GEN_5239;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h76 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_118_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_118_rob_idx <= _GEN_5367;
      end
    end else begin
      rob_payload_118_rob_idx <= _GEN_5367;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h76 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_118_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_118_flits_fired <= _GEN_13572;
      end
    end else begin
      rob_payload_118_flits_fired <= _GEN_13572;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h77 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_119_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_119_tsc <= _GEN_5240;
      end
    end else begin
      rob_payload_119_tsc <= _GEN_5240;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h77 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_119_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_119_rob_idx <= _GEN_5368;
      end
    end else begin
      rob_payload_119_rob_idx <= _GEN_5368;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h77 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_119_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_119_flits_fired <= _GEN_13573;
      end
    end else begin
      rob_payload_119_flits_fired <= _GEN_13573;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h78 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_120_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_120_tsc <= _GEN_5241;
      end
    end else begin
      rob_payload_120_tsc <= _GEN_5241;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h78 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_120_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_120_rob_idx <= _GEN_5369;
      end
    end else begin
      rob_payload_120_rob_idx <= _GEN_5369;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h78 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_120_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_120_flits_fired <= _GEN_13574;
      end
    end else begin
      rob_payload_120_flits_fired <= _GEN_13574;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h79 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_121_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_121_tsc <= _GEN_5242;
      end
    end else begin
      rob_payload_121_tsc <= _GEN_5242;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h79 == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_121_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_121_rob_idx <= _GEN_5370;
      end
    end else begin
      rob_payload_121_rob_idx <= _GEN_5370;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h79 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_121_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_121_flits_fired <= _GEN_13575;
      end
    end else begin
      rob_payload_121_flits_fired <= _GEN_13575;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7a == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_122_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_122_tsc <= _GEN_5243;
      end
    end else begin
      rob_payload_122_tsc <= _GEN_5243;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7a == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_122_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_122_rob_idx <= _GEN_5371;
      end
    end else begin
      rob_payload_122_rob_idx <= _GEN_5371;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h7a == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_122_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_122_flits_fired <= _GEN_13576;
      end
    end else begin
      rob_payload_122_flits_fired <= _GEN_13576;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7b == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_123_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_123_tsc <= _GEN_5244;
      end
    end else begin
      rob_payload_123_tsc <= _GEN_5244;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7b == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_123_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_123_rob_idx <= _GEN_5372;
      end
    end else begin
      rob_payload_123_rob_idx <= _GEN_5372;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h7b == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_123_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_123_flits_fired <= _GEN_13577;
      end
    end else begin
      rob_payload_123_flits_fired <= _GEN_13577;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7c == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_124_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_124_tsc <= _GEN_5245;
      end
    end else begin
      rob_payload_124_tsc <= _GEN_5245;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7c == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_124_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_124_rob_idx <= _GEN_5373;
      end
    end else begin
      rob_payload_124_rob_idx <= _GEN_5373;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h7c == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_124_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_124_flits_fired <= _GEN_13578;
      end
    end else begin
      rob_payload_124_flits_fired <= _GEN_13578;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7d == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_125_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_125_tsc <= _GEN_5246;
      end
    end else begin
      rob_payload_125_tsc <= _GEN_5246;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7d == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_125_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_125_rob_idx <= _GEN_5374;
      end
    end else begin
      rob_payload_125_rob_idx <= _GEN_5374;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h7d == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_125_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_125_flits_fired <= _GEN_13579;
      end
    end else begin
      rob_payload_125_flits_fired <= _GEN_13579;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7e == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_126_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_126_tsc <= _GEN_5247;
      end
    end else begin
      rob_payload_126_tsc <= _GEN_5247;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7e == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_126_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_126_rob_idx <= _GEN_5375;
      end
    end else begin
      rob_payload_126_rob_idx <= _GEN_5375;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h7e == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_126_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_126_flits_fired <= _GEN_13580;
      end
    end else begin
      rob_payload_126_flits_fired <= _GEN_13580;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7f == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_127_tsc <= _rob_payload_WIRE_7[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_127_tsc <= _GEN_5248;
      end
    end else begin
      rob_payload_127_tsc <= _GEN_5248;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7f == rob_alloc_ids_3) begin // @[TestHarness.scala 179:36]
        rob_payload_127_rob_idx <= _rob_payload_WIRE_7[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_127_rob_idx <= _GEN_5376;
      end
    end else begin
      rob_payload_127_rob_idx <= _GEN_5376;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h7f == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_127_flits_fired <= _rob_payload_flits_fired_T_11; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_127_flits_fired <= _GEN_13581;
      end
    end else begin
      rob_payload_127_flits_fired <= _GEN_13581;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h0 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_0 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_0 <= _GEN_5505;
      end
    end else begin
      rob_egress_id_0 <= _GEN_5505;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_1 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_1 <= _GEN_5506;
      end
    end else begin
      rob_egress_id_1 <= _GEN_5506;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_2 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_2 <= _GEN_5507;
      end
    end else begin
      rob_egress_id_2 <= _GEN_5507;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_3 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_3 <= _GEN_5508;
      end
    end else begin
      rob_egress_id_3 <= _GEN_5508;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_4 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_4 <= _GEN_5509;
      end
    end else begin
      rob_egress_id_4 <= _GEN_5509;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_5 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_5 <= _GEN_5510;
      end
    end else begin
      rob_egress_id_5 <= _GEN_5510;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_6 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_6 <= _GEN_5511;
      end
    end else begin
      rob_egress_id_6 <= _GEN_5511;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_7 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_7 <= _GEN_5512;
      end
    end else begin
      rob_egress_id_7 <= _GEN_5512;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h8 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_8 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_8 <= _GEN_5513;
      end
    end else begin
      rob_egress_id_8 <= _GEN_5513;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h9 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_9 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_9 <= _GEN_5514;
      end
    end else begin
      rob_egress_id_9 <= _GEN_5514;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'ha == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_10 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_10 <= _GEN_5515;
      end
    end else begin
      rob_egress_id_10 <= _GEN_5515;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hb == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_11 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_11 <= _GEN_5516;
      end
    end else begin
      rob_egress_id_11 <= _GEN_5516;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hc == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_12 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_12 <= _GEN_5517;
      end
    end else begin
      rob_egress_id_12 <= _GEN_5517;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hd == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_13 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_13 <= _GEN_5518;
      end
    end else begin
      rob_egress_id_13 <= _GEN_5518;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'he == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_14 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_14 <= _GEN_5519;
      end
    end else begin
      rob_egress_id_14 <= _GEN_5519;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hf == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_15 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_15 <= _GEN_5520;
      end
    end else begin
      rob_egress_id_15 <= _GEN_5520;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h10 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_16 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_16 <= _GEN_5521;
      end
    end else begin
      rob_egress_id_16 <= _GEN_5521;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h11 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_17 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_17 <= _GEN_5522;
      end
    end else begin
      rob_egress_id_17 <= _GEN_5522;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h12 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_18 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_18 <= _GEN_5523;
      end
    end else begin
      rob_egress_id_18 <= _GEN_5523;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h13 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_19 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_19 <= _GEN_5524;
      end
    end else begin
      rob_egress_id_19 <= _GEN_5524;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h14 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_20 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_20 <= _GEN_5525;
      end
    end else begin
      rob_egress_id_20 <= _GEN_5525;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h15 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_21 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_21 <= _GEN_5526;
      end
    end else begin
      rob_egress_id_21 <= _GEN_5526;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h16 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_22 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_22 <= _GEN_5527;
      end
    end else begin
      rob_egress_id_22 <= _GEN_5527;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h17 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_23 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_23 <= _GEN_5528;
      end
    end else begin
      rob_egress_id_23 <= _GEN_5528;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h18 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_24 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_24 <= _GEN_5529;
      end
    end else begin
      rob_egress_id_24 <= _GEN_5529;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h19 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_25 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_25 <= _GEN_5530;
      end
    end else begin
      rob_egress_id_25 <= _GEN_5530;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1a == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_26 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_26 <= _GEN_5531;
      end
    end else begin
      rob_egress_id_26 <= _GEN_5531;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1b == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_27 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_27 <= _GEN_5532;
      end
    end else begin
      rob_egress_id_27 <= _GEN_5532;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1c == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_28 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_28 <= _GEN_5533;
      end
    end else begin
      rob_egress_id_28 <= _GEN_5533;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1d == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_29 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_29 <= _GEN_5534;
      end
    end else begin
      rob_egress_id_29 <= _GEN_5534;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1e == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_30 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_30 <= _GEN_5535;
      end
    end else begin
      rob_egress_id_30 <= _GEN_5535;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1f == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_31 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_31 <= _GEN_5536;
      end
    end else begin
      rob_egress_id_31 <= _GEN_5536;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h20 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_32 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_32 <= _GEN_5537;
      end
    end else begin
      rob_egress_id_32 <= _GEN_5537;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h21 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_33 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_33 <= _GEN_5538;
      end
    end else begin
      rob_egress_id_33 <= _GEN_5538;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h22 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_34 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_34 <= _GEN_5539;
      end
    end else begin
      rob_egress_id_34 <= _GEN_5539;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h23 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_35 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_35 <= _GEN_5540;
      end
    end else begin
      rob_egress_id_35 <= _GEN_5540;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h24 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_36 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_36 <= _GEN_5541;
      end
    end else begin
      rob_egress_id_36 <= _GEN_5541;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h25 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_37 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_37 <= _GEN_5542;
      end
    end else begin
      rob_egress_id_37 <= _GEN_5542;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h26 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_38 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_38 <= _GEN_5543;
      end
    end else begin
      rob_egress_id_38 <= _GEN_5543;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h27 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_39 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_39 <= _GEN_5544;
      end
    end else begin
      rob_egress_id_39 <= _GEN_5544;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h28 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_40 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_40 <= _GEN_5545;
      end
    end else begin
      rob_egress_id_40 <= _GEN_5545;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h29 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_41 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_41 <= _GEN_5546;
      end
    end else begin
      rob_egress_id_41 <= _GEN_5546;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2a == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_42 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_42 <= _GEN_5547;
      end
    end else begin
      rob_egress_id_42 <= _GEN_5547;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2b == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_43 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_43 <= _GEN_5548;
      end
    end else begin
      rob_egress_id_43 <= _GEN_5548;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2c == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_44 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_44 <= _GEN_5549;
      end
    end else begin
      rob_egress_id_44 <= _GEN_5549;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2d == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_45 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_45 <= _GEN_5550;
      end
    end else begin
      rob_egress_id_45 <= _GEN_5550;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2e == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_46 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_46 <= _GEN_5551;
      end
    end else begin
      rob_egress_id_46 <= _GEN_5551;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2f == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_47 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_47 <= _GEN_5552;
      end
    end else begin
      rob_egress_id_47 <= _GEN_5552;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h30 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_48 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_48 <= _GEN_5553;
      end
    end else begin
      rob_egress_id_48 <= _GEN_5553;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h31 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_49 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_49 <= _GEN_5554;
      end
    end else begin
      rob_egress_id_49 <= _GEN_5554;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h32 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_50 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_50 <= _GEN_5555;
      end
    end else begin
      rob_egress_id_50 <= _GEN_5555;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h33 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_51 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_51 <= _GEN_5556;
      end
    end else begin
      rob_egress_id_51 <= _GEN_5556;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h34 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_52 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_52 <= _GEN_5557;
      end
    end else begin
      rob_egress_id_52 <= _GEN_5557;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h35 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_53 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_53 <= _GEN_5558;
      end
    end else begin
      rob_egress_id_53 <= _GEN_5558;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h36 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_54 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_54 <= _GEN_5559;
      end
    end else begin
      rob_egress_id_54 <= _GEN_5559;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h37 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_55 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_55 <= _GEN_5560;
      end
    end else begin
      rob_egress_id_55 <= _GEN_5560;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h38 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_56 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_56 <= _GEN_5561;
      end
    end else begin
      rob_egress_id_56 <= _GEN_5561;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h39 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_57 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_57 <= _GEN_5562;
      end
    end else begin
      rob_egress_id_57 <= _GEN_5562;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3a == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_58 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_58 <= _GEN_5563;
      end
    end else begin
      rob_egress_id_58 <= _GEN_5563;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3b == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_59 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_59 <= _GEN_5564;
      end
    end else begin
      rob_egress_id_59 <= _GEN_5564;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3c == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_60 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_60 <= _GEN_5565;
      end
    end else begin
      rob_egress_id_60 <= _GEN_5565;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3d == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_61 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_61 <= _GEN_5566;
      end
    end else begin
      rob_egress_id_61 <= _GEN_5566;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3e == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_62 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_62 <= _GEN_5567;
      end
    end else begin
      rob_egress_id_62 <= _GEN_5567;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3f == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_63 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_63 <= _GEN_5568;
      end
    end else begin
      rob_egress_id_63 <= _GEN_5568;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h40 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_64 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_64 <= _GEN_5569;
      end
    end else begin
      rob_egress_id_64 <= _GEN_5569;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h41 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_65 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_65 <= _GEN_5570;
      end
    end else begin
      rob_egress_id_65 <= _GEN_5570;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h42 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_66 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_66 <= _GEN_5571;
      end
    end else begin
      rob_egress_id_66 <= _GEN_5571;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h43 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_67 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_67 <= _GEN_5572;
      end
    end else begin
      rob_egress_id_67 <= _GEN_5572;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h44 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_68 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_68 <= _GEN_5573;
      end
    end else begin
      rob_egress_id_68 <= _GEN_5573;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h45 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_69 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_69 <= _GEN_5574;
      end
    end else begin
      rob_egress_id_69 <= _GEN_5574;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h46 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_70 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_70 <= _GEN_5575;
      end
    end else begin
      rob_egress_id_70 <= _GEN_5575;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h47 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_71 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_71 <= _GEN_5576;
      end
    end else begin
      rob_egress_id_71 <= _GEN_5576;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h48 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_72 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_72 <= _GEN_5577;
      end
    end else begin
      rob_egress_id_72 <= _GEN_5577;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h49 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_73 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_73 <= _GEN_5578;
      end
    end else begin
      rob_egress_id_73 <= _GEN_5578;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4a == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_74 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_74 <= _GEN_5579;
      end
    end else begin
      rob_egress_id_74 <= _GEN_5579;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4b == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_75 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_75 <= _GEN_5580;
      end
    end else begin
      rob_egress_id_75 <= _GEN_5580;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4c == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_76 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_76 <= _GEN_5581;
      end
    end else begin
      rob_egress_id_76 <= _GEN_5581;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4d == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_77 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_77 <= _GEN_5582;
      end
    end else begin
      rob_egress_id_77 <= _GEN_5582;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4e == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_78 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_78 <= _GEN_5583;
      end
    end else begin
      rob_egress_id_78 <= _GEN_5583;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4f == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_79 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_79 <= _GEN_5584;
      end
    end else begin
      rob_egress_id_79 <= _GEN_5584;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h50 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_80 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_80 <= _GEN_5585;
      end
    end else begin
      rob_egress_id_80 <= _GEN_5585;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h51 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_81 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_81 <= _GEN_5586;
      end
    end else begin
      rob_egress_id_81 <= _GEN_5586;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h52 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_82 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_82 <= _GEN_5587;
      end
    end else begin
      rob_egress_id_82 <= _GEN_5587;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h53 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_83 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_83 <= _GEN_5588;
      end
    end else begin
      rob_egress_id_83 <= _GEN_5588;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h54 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_84 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_84 <= _GEN_5589;
      end
    end else begin
      rob_egress_id_84 <= _GEN_5589;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h55 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_85 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_85 <= _GEN_5590;
      end
    end else begin
      rob_egress_id_85 <= _GEN_5590;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h56 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_86 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_86 <= _GEN_5591;
      end
    end else begin
      rob_egress_id_86 <= _GEN_5591;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h57 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_87 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_87 <= _GEN_5592;
      end
    end else begin
      rob_egress_id_87 <= _GEN_5592;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h58 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_88 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_88 <= _GEN_5593;
      end
    end else begin
      rob_egress_id_88 <= _GEN_5593;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h59 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_89 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_89 <= _GEN_5594;
      end
    end else begin
      rob_egress_id_89 <= _GEN_5594;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5a == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_90 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_90 <= _GEN_5595;
      end
    end else begin
      rob_egress_id_90 <= _GEN_5595;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5b == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_91 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_91 <= _GEN_5596;
      end
    end else begin
      rob_egress_id_91 <= _GEN_5596;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5c == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_92 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_92 <= _GEN_5597;
      end
    end else begin
      rob_egress_id_92 <= _GEN_5597;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5d == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_93 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_93 <= _GEN_5598;
      end
    end else begin
      rob_egress_id_93 <= _GEN_5598;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5e == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_94 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_94 <= _GEN_5599;
      end
    end else begin
      rob_egress_id_94 <= _GEN_5599;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5f == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_95 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_95 <= _GEN_5600;
      end
    end else begin
      rob_egress_id_95 <= _GEN_5600;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h60 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_96 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_96 <= _GEN_5601;
      end
    end else begin
      rob_egress_id_96 <= _GEN_5601;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h61 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_97 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_97 <= _GEN_5602;
      end
    end else begin
      rob_egress_id_97 <= _GEN_5602;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h62 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_98 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_98 <= _GEN_5603;
      end
    end else begin
      rob_egress_id_98 <= _GEN_5603;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h63 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_99 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_99 <= _GEN_5604;
      end
    end else begin
      rob_egress_id_99 <= _GEN_5604;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h64 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_100 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_100 <= _GEN_5605;
      end
    end else begin
      rob_egress_id_100 <= _GEN_5605;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h65 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_101 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_101 <= _GEN_5606;
      end
    end else begin
      rob_egress_id_101 <= _GEN_5606;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h66 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_102 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_102 <= _GEN_5607;
      end
    end else begin
      rob_egress_id_102 <= _GEN_5607;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h67 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_103 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_103 <= _GEN_5608;
      end
    end else begin
      rob_egress_id_103 <= _GEN_5608;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h68 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_104 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_104 <= _GEN_5609;
      end
    end else begin
      rob_egress_id_104 <= _GEN_5609;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h69 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_105 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_105 <= _GEN_5610;
      end
    end else begin
      rob_egress_id_105 <= _GEN_5610;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6a == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_106 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_106 <= _GEN_5611;
      end
    end else begin
      rob_egress_id_106 <= _GEN_5611;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6b == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_107 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_107 <= _GEN_5612;
      end
    end else begin
      rob_egress_id_107 <= _GEN_5612;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6c == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_108 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_108 <= _GEN_5613;
      end
    end else begin
      rob_egress_id_108 <= _GEN_5613;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6d == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_109 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_109 <= _GEN_5614;
      end
    end else begin
      rob_egress_id_109 <= _GEN_5614;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6e == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_110 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_110 <= _GEN_5615;
      end
    end else begin
      rob_egress_id_110 <= _GEN_5615;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6f == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_111 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_111 <= _GEN_5616;
      end
    end else begin
      rob_egress_id_111 <= _GEN_5616;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h70 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_112 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_112 <= _GEN_5617;
      end
    end else begin
      rob_egress_id_112 <= _GEN_5617;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h71 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_113 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_113 <= _GEN_5618;
      end
    end else begin
      rob_egress_id_113 <= _GEN_5618;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h72 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_114 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_114 <= _GEN_5619;
      end
    end else begin
      rob_egress_id_114 <= _GEN_5619;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h73 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_115 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_115 <= _GEN_5620;
      end
    end else begin
      rob_egress_id_115 <= _GEN_5620;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h74 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_116 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_116 <= _GEN_5621;
      end
    end else begin
      rob_egress_id_116 <= _GEN_5621;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h75 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_117 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_117 <= _GEN_5622;
      end
    end else begin
      rob_egress_id_117 <= _GEN_5622;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h76 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_118 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_118 <= _GEN_5623;
      end
    end else begin
      rob_egress_id_118 <= _GEN_5623;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h77 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_119 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_119 <= _GEN_5624;
      end
    end else begin
      rob_egress_id_119 <= _GEN_5624;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h78 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_120 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_120 <= _GEN_5625;
      end
    end else begin
      rob_egress_id_120 <= _GEN_5625;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h79 == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_121 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_121 <= _GEN_5626;
      end
    end else begin
      rob_egress_id_121 <= _GEN_5626;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7a == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_122 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_122 <= _GEN_5627;
      end
    end else begin
      rob_egress_id_122 <= _GEN_5627;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7b == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_123 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_123 <= _GEN_5628;
      end
    end else begin
      rob_egress_id_123 <= _GEN_5628;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7c == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_124 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_124 <= _GEN_5629;
      end
    end else begin
      rob_egress_id_124 <= _GEN_5629;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7d == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_125 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_125 <= _GEN_5630;
      end
    end else begin
      rob_egress_id_125 <= _GEN_5630;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7e == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_126 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_126 <= _GEN_5631;
      end
    end else begin
      rob_egress_id_126 <= _GEN_5631;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7f == rob_alloc_ids_3) begin // @[TestHarness.scala 180:36]
        rob_egress_id_127 <= _rob_egress_id_T_65; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_127 <= _GEN_5632;
      end
    end else begin
      rob_egress_id_127 <= _GEN_5632;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h0 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_0 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_0 <= _GEN_5633;
      end
    end else begin
      rob_ingress_id_0 <= _GEN_5633;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_1 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_1 <= _GEN_5634;
      end
    end else begin
      rob_ingress_id_1 <= _GEN_5634;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_2 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_2 <= _GEN_5635;
      end
    end else begin
      rob_ingress_id_2 <= _GEN_5635;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_3 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_3 <= _GEN_5636;
      end
    end else begin
      rob_ingress_id_3 <= _GEN_5636;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_4 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_4 <= _GEN_5637;
      end
    end else begin
      rob_ingress_id_4 <= _GEN_5637;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_5 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_5 <= _GEN_5638;
      end
    end else begin
      rob_ingress_id_5 <= _GEN_5638;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_6 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_6 <= _GEN_5639;
      end
    end else begin
      rob_ingress_id_6 <= _GEN_5639;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_7 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_7 <= _GEN_5640;
      end
    end else begin
      rob_ingress_id_7 <= _GEN_5640;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h8 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_8 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_8 <= _GEN_5641;
      end
    end else begin
      rob_ingress_id_8 <= _GEN_5641;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h9 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_9 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_9 <= _GEN_5642;
      end
    end else begin
      rob_ingress_id_9 <= _GEN_5642;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'ha == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_10 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_10 <= _GEN_5643;
      end
    end else begin
      rob_ingress_id_10 <= _GEN_5643;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hb == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_11 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_11 <= _GEN_5644;
      end
    end else begin
      rob_ingress_id_11 <= _GEN_5644;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hc == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_12 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_12 <= _GEN_5645;
      end
    end else begin
      rob_ingress_id_12 <= _GEN_5645;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hd == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_13 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_13 <= _GEN_5646;
      end
    end else begin
      rob_ingress_id_13 <= _GEN_5646;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'he == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_14 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_14 <= _GEN_5647;
      end
    end else begin
      rob_ingress_id_14 <= _GEN_5647;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hf == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_15 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_15 <= _GEN_5648;
      end
    end else begin
      rob_ingress_id_15 <= _GEN_5648;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h10 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_16 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_16 <= _GEN_5649;
      end
    end else begin
      rob_ingress_id_16 <= _GEN_5649;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h11 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_17 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_17 <= _GEN_5650;
      end
    end else begin
      rob_ingress_id_17 <= _GEN_5650;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h12 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_18 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_18 <= _GEN_5651;
      end
    end else begin
      rob_ingress_id_18 <= _GEN_5651;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h13 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_19 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_19 <= _GEN_5652;
      end
    end else begin
      rob_ingress_id_19 <= _GEN_5652;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h14 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_20 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_20 <= _GEN_5653;
      end
    end else begin
      rob_ingress_id_20 <= _GEN_5653;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h15 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_21 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_21 <= _GEN_5654;
      end
    end else begin
      rob_ingress_id_21 <= _GEN_5654;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h16 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_22 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_22 <= _GEN_5655;
      end
    end else begin
      rob_ingress_id_22 <= _GEN_5655;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h17 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_23 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_23 <= _GEN_5656;
      end
    end else begin
      rob_ingress_id_23 <= _GEN_5656;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h18 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_24 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_24 <= _GEN_5657;
      end
    end else begin
      rob_ingress_id_24 <= _GEN_5657;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h19 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_25 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_25 <= _GEN_5658;
      end
    end else begin
      rob_ingress_id_25 <= _GEN_5658;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1a == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_26 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_26 <= _GEN_5659;
      end
    end else begin
      rob_ingress_id_26 <= _GEN_5659;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1b == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_27 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_27 <= _GEN_5660;
      end
    end else begin
      rob_ingress_id_27 <= _GEN_5660;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1c == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_28 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_28 <= _GEN_5661;
      end
    end else begin
      rob_ingress_id_28 <= _GEN_5661;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1d == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_29 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_29 <= _GEN_5662;
      end
    end else begin
      rob_ingress_id_29 <= _GEN_5662;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1e == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_30 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_30 <= _GEN_5663;
      end
    end else begin
      rob_ingress_id_30 <= _GEN_5663;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1f == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_31 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_31 <= _GEN_5664;
      end
    end else begin
      rob_ingress_id_31 <= _GEN_5664;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h20 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_32 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_32 <= _GEN_5665;
      end
    end else begin
      rob_ingress_id_32 <= _GEN_5665;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h21 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_33 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_33 <= _GEN_5666;
      end
    end else begin
      rob_ingress_id_33 <= _GEN_5666;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h22 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_34 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_34 <= _GEN_5667;
      end
    end else begin
      rob_ingress_id_34 <= _GEN_5667;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h23 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_35 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_35 <= _GEN_5668;
      end
    end else begin
      rob_ingress_id_35 <= _GEN_5668;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h24 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_36 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_36 <= _GEN_5669;
      end
    end else begin
      rob_ingress_id_36 <= _GEN_5669;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h25 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_37 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_37 <= _GEN_5670;
      end
    end else begin
      rob_ingress_id_37 <= _GEN_5670;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h26 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_38 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_38 <= _GEN_5671;
      end
    end else begin
      rob_ingress_id_38 <= _GEN_5671;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h27 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_39 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_39 <= _GEN_5672;
      end
    end else begin
      rob_ingress_id_39 <= _GEN_5672;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h28 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_40 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_40 <= _GEN_5673;
      end
    end else begin
      rob_ingress_id_40 <= _GEN_5673;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h29 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_41 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_41 <= _GEN_5674;
      end
    end else begin
      rob_ingress_id_41 <= _GEN_5674;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2a == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_42 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_42 <= _GEN_5675;
      end
    end else begin
      rob_ingress_id_42 <= _GEN_5675;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2b == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_43 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_43 <= _GEN_5676;
      end
    end else begin
      rob_ingress_id_43 <= _GEN_5676;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2c == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_44 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_44 <= _GEN_5677;
      end
    end else begin
      rob_ingress_id_44 <= _GEN_5677;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2d == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_45 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_45 <= _GEN_5678;
      end
    end else begin
      rob_ingress_id_45 <= _GEN_5678;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2e == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_46 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_46 <= _GEN_5679;
      end
    end else begin
      rob_ingress_id_46 <= _GEN_5679;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2f == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_47 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_47 <= _GEN_5680;
      end
    end else begin
      rob_ingress_id_47 <= _GEN_5680;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h30 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_48 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_48 <= _GEN_5681;
      end
    end else begin
      rob_ingress_id_48 <= _GEN_5681;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h31 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_49 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_49 <= _GEN_5682;
      end
    end else begin
      rob_ingress_id_49 <= _GEN_5682;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h32 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_50 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_50 <= _GEN_5683;
      end
    end else begin
      rob_ingress_id_50 <= _GEN_5683;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h33 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_51 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_51 <= _GEN_5684;
      end
    end else begin
      rob_ingress_id_51 <= _GEN_5684;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h34 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_52 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_52 <= _GEN_5685;
      end
    end else begin
      rob_ingress_id_52 <= _GEN_5685;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h35 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_53 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_53 <= _GEN_5686;
      end
    end else begin
      rob_ingress_id_53 <= _GEN_5686;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h36 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_54 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_54 <= _GEN_5687;
      end
    end else begin
      rob_ingress_id_54 <= _GEN_5687;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h37 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_55 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_55 <= _GEN_5688;
      end
    end else begin
      rob_ingress_id_55 <= _GEN_5688;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h38 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_56 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_56 <= _GEN_5689;
      end
    end else begin
      rob_ingress_id_56 <= _GEN_5689;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h39 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_57 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_57 <= _GEN_5690;
      end
    end else begin
      rob_ingress_id_57 <= _GEN_5690;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3a == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_58 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_58 <= _GEN_5691;
      end
    end else begin
      rob_ingress_id_58 <= _GEN_5691;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3b == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_59 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_59 <= _GEN_5692;
      end
    end else begin
      rob_ingress_id_59 <= _GEN_5692;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3c == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_60 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_60 <= _GEN_5693;
      end
    end else begin
      rob_ingress_id_60 <= _GEN_5693;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3d == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_61 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_61 <= _GEN_5694;
      end
    end else begin
      rob_ingress_id_61 <= _GEN_5694;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3e == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_62 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_62 <= _GEN_5695;
      end
    end else begin
      rob_ingress_id_62 <= _GEN_5695;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3f == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_63 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_63 <= _GEN_5696;
      end
    end else begin
      rob_ingress_id_63 <= _GEN_5696;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h40 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_64 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_64 <= _GEN_5697;
      end
    end else begin
      rob_ingress_id_64 <= _GEN_5697;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h41 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_65 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_65 <= _GEN_5698;
      end
    end else begin
      rob_ingress_id_65 <= _GEN_5698;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h42 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_66 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_66 <= _GEN_5699;
      end
    end else begin
      rob_ingress_id_66 <= _GEN_5699;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h43 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_67 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_67 <= _GEN_5700;
      end
    end else begin
      rob_ingress_id_67 <= _GEN_5700;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h44 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_68 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_68 <= _GEN_5701;
      end
    end else begin
      rob_ingress_id_68 <= _GEN_5701;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h45 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_69 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_69 <= _GEN_5702;
      end
    end else begin
      rob_ingress_id_69 <= _GEN_5702;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h46 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_70 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_70 <= _GEN_5703;
      end
    end else begin
      rob_ingress_id_70 <= _GEN_5703;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h47 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_71 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_71 <= _GEN_5704;
      end
    end else begin
      rob_ingress_id_71 <= _GEN_5704;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h48 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_72 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_72 <= _GEN_5705;
      end
    end else begin
      rob_ingress_id_72 <= _GEN_5705;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h49 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_73 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_73 <= _GEN_5706;
      end
    end else begin
      rob_ingress_id_73 <= _GEN_5706;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4a == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_74 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_74 <= _GEN_5707;
      end
    end else begin
      rob_ingress_id_74 <= _GEN_5707;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4b == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_75 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_75 <= _GEN_5708;
      end
    end else begin
      rob_ingress_id_75 <= _GEN_5708;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4c == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_76 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_76 <= _GEN_5709;
      end
    end else begin
      rob_ingress_id_76 <= _GEN_5709;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4d == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_77 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_77 <= _GEN_5710;
      end
    end else begin
      rob_ingress_id_77 <= _GEN_5710;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4e == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_78 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_78 <= _GEN_5711;
      end
    end else begin
      rob_ingress_id_78 <= _GEN_5711;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4f == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_79 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_79 <= _GEN_5712;
      end
    end else begin
      rob_ingress_id_79 <= _GEN_5712;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h50 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_80 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_80 <= _GEN_5713;
      end
    end else begin
      rob_ingress_id_80 <= _GEN_5713;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h51 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_81 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_81 <= _GEN_5714;
      end
    end else begin
      rob_ingress_id_81 <= _GEN_5714;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h52 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_82 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_82 <= _GEN_5715;
      end
    end else begin
      rob_ingress_id_82 <= _GEN_5715;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h53 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_83 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_83 <= _GEN_5716;
      end
    end else begin
      rob_ingress_id_83 <= _GEN_5716;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h54 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_84 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_84 <= _GEN_5717;
      end
    end else begin
      rob_ingress_id_84 <= _GEN_5717;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h55 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_85 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_85 <= _GEN_5718;
      end
    end else begin
      rob_ingress_id_85 <= _GEN_5718;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h56 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_86 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_86 <= _GEN_5719;
      end
    end else begin
      rob_ingress_id_86 <= _GEN_5719;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h57 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_87 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_87 <= _GEN_5720;
      end
    end else begin
      rob_ingress_id_87 <= _GEN_5720;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h58 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_88 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_88 <= _GEN_5721;
      end
    end else begin
      rob_ingress_id_88 <= _GEN_5721;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h59 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_89 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_89 <= _GEN_5722;
      end
    end else begin
      rob_ingress_id_89 <= _GEN_5722;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5a == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_90 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_90 <= _GEN_5723;
      end
    end else begin
      rob_ingress_id_90 <= _GEN_5723;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5b == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_91 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_91 <= _GEN_5724;
      end
    end else begin
      rob_ingress_id_91 <= _GEN_5724;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5c == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_92 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_92 <= _GEN_5725;
      end
    end else begin
      rob_ingress_id_92 <= _GEN_5725;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5d == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_93 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_93 <= _GEN_5726;
      end
    end else begin
      rob_ingress_id_93 <= _GEN_5726;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5e == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_94 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_94 <= _GEN_5727;
      end
    end else begin
      rob_ingress_id_94 <= _GEN_5727;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5f == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_95 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_95 <= _GEN_5728;
      end
    end else begin
      rob_ingress_id_95 <= _GEN_5728;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h60 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_96 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_96 <= _GEN_5729;
      end
    end else begin
      rob_ingress_id_96 <= _GEN_5729;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h61 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_97 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_97 <= _GEN_5730;
      end
    end else begin
      rob_ingress_id_97 <= _GEN_5730;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h62 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_98 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_98 <= _GEN_5731;
      end
    end else begin
      rob_ingress_id_98 <= _GEN_5731;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h63 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_99 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_99 <= _GEN_5732;
      end
    end else begin
      rob_ingress_id_99 <= _GEN_5732;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h64 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_100 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_100 <= _GEN_5733;
      end
    end else begin
      rob_ingress_id_100 <= _GEN_5733;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h65 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_101 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_101 <= _GEN_5734;
      end
    end else begin
      rob_ingress_id_101 <= _GEN_5734;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h66 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_102 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_102 <= _GEN_5735;
      end
    end else begin
      rob_ingress_id_102 <= _GEN_5735;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h67 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_103 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_103 <= _GEN_5736;
      end
    end else begin
      rob_ingress_id_103 <= _GEN_5736;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h68 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_104 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_104 <= _GEN_5737;
      end
    end else begin
      rob_ingress_id_104 <= _GEN_5737;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h69 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_105 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_105 <= _GEN_5738;
      end
    end else begin
      rob_ingress_id_105 <= _GEN_5738;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6a == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_106 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_106 <= _GEN_5739;
      end
    end else begin
      rob_ingress_id_106 <= _GEN_5739;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6b == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_107 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_107 <= _GEN_5740;
      end
    end else begin
      rob_ingress_id_107 <= _GEN_5740;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6c == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_108 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_108 <= _GEN_5741;
      end
    end else begin
      rob_ingress_id_108 <= _GEN_5741;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6d == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_109 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_109 <= _GEN_5742;
      end
    end else begin
      rob_ingress_id_109 <= _GEN_5742;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6e == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_110 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_110 <= _GEN_5743;
      end
    end else begin
      rob_ingress_id_110 <= _GEN_5743;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6f == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_111 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_111 <= _GEN_5744;
      end
    end else begin
      rob_ingress_id_111 <= _GEN_5744;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h70 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_112 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_112 <= _GEN_5745;
      end
    end else begin
      rob_ingress_id_112 <= _GEN_5745;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h71 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_113 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_113 <= _GEN_5746;
      end
    end else begin
      rob_ingress_id_113 <= _GEN_5746;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h72 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_114 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_114 <= _GEN_5747;
      end
    end else begin
      rob_ingress_id_114 <= _GEN_5747;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h73 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_115 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_115 <= _GEN_5748;
      end
    end else begin
      rob_ingress_id_115 <= _GEN_5748;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h74 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_116 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_116 <= _GEN_5749;
      end
    end else begin
      rob_ingress_id_116 <= _GEN_5749;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h75 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_117 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_117 <= _GEN_5750;
      end
    end else begin
      rob_ingress_id_117 <= _GEN_5750;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h76 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_118 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_118 <= _GEN_5751;
      end
    end else begin
      rob_ingress_id_118 <= _GEN_5751;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h77 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_119 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_119 <= _GEN_5752;
      end
    end else begin
      rob_ingress_id_119 <= _GEN_5752;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h78 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_120 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_120 <= _GEN_5753;
      end
    end else begin
      rob_ingress_id_120 <= _GEN_5753;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h79 == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_121 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_121 <= _GEN_5754;
      end
    end else begin
      rob_ingress_id_121 <= _GEN_5754;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7a == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_122 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_122 <= _GEN_5755;
      end
    end else begin
      rob_ingress_id_122 <= _GEN_5755;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7b == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_123 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_123 <= _GEN_5756;
      end
    end else begin
      rob_ingress_id_123 <= _GEN_5756;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7c == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_124 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_124 <= _GEN_5757;
      end
    end else begin
      rob_ingress_id_124 <= _GEN_5757;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7d == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_125 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_125 <= _GEN_5758;
      end
    end else begin
      rob_ingress_id_125 <= _GEN_5758;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7e == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_126 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_126 <= _GEN_5759;
      end
    end else begin
      rob_ingress_id_126 <= _GEN_5759;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7f == rob_alloc_ids_3) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_127 <= 2'h3; // @[TestHarness.scala 181:36]
      end else begin
        rob_ingress_id_127 <= _GEN_5760;
      end
    end else begin
      rob_ingress_id_127 <= _GEN_5760;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h0 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_0 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_0 <= _GEN_5761;
      end
    end else begin
      rob_n_flits_0 <= _GEN_5761;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_1 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_1 <= _GEN_5762;
      end
    end else begin
      rob_n_flits_1 <= _GEN_5762;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_2 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_2 <= _GEN_5763;
      end
    end else begin
      rob_n_flits_2 <= _GEN_5763;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_3 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_3 <= _GEN_5764;
      end
    end else begin
      rob_n_flits_3 <= _GEN_5764;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_4 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_4 <= _GEN_5765;
      end
    end else begin
      rob_n_flits_4 <= _GEN_5765;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_5 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_5 <= _GEN_5766;
      end
    end else begin
      rob_n_flits_5 <= _GEN_5766;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_6 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_6 <= _GEN_5767;
      end
    end else begin
      rob_n_flits_6 <= _GEN_5767;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_7 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_7 <= _GEN_5768;
      end
    end else begin
      rob_n_flits_7 <= _GEN_5768;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h8 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_8 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_8 <= _GEN_5769;
      end
    end else begin
      rob_n_flits_8 <= _GEN_5769;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h9 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_9 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_9 <= _GEN_5770;
      end
    end else begin
      rob_n_flits_9 <= _GEN_5770;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'ha == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_10 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_10 <= _GEN_5771;
      end
    end else begin
      rob_n_flits_10 <= _GEN_5771;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hb == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_11 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_11 <= _GEN_5772;
      end
    end else begin
      rob_n_flits_11 <= _GEN_5772;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hc == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_12 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_12 <= _GEN_5773;
      end
    end else begin
      rob_n_flits_12 <= _GEN_5773;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hd == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_13 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_13 <= _GEN_5774;
      end
    end else begin
      rob_n_flits_13 <= _GEN_5774;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'he == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_14 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_14 <= _GEN_5775;
      end
    end else begin
      rob_n_flits_14 <= _GEN_5775;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hf == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_15 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_15 <= _GEN_5776;
      end
    end else begin
      rob_n_flits_15 <= _GEN_5776;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h10 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_16 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_16 <= _GEN_5777;
      end
    end else begin
      rob_n_flits_16 <= _GEN_5777;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h11 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_17 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_17 <= _GEN_5778;
      end
    end else begin
      rob_n_flits_17 <= _GEN_5778;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h12 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_18 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_18 <= _GEN_5779;
      end
    end else begin
      rob_n_flits_18 <= _GEN_5779;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h13 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_19 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_19 <= _GEN_5780;
      end
    end else begin
      rob_n_flits_19 <= _GEN_5780;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h14 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_20 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_20 <= _GEN_5781;
      end
    end else begin
      rob_n_flits_20 <= _GEN_5781;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h15 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_21 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_21 <= _GEN_5782;
      end
    end else begin
      rob_n_flits_21 <= _GEN_5782;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h16 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_22 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_22 <= _GEN_5783;
      end
    end else begin
      rob_n_flits_22 <= _GEN_5783;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h17 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_23 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_23 <= _GEN_5784;
      end
    end else begin
      rob_n_flits_23 <= _GEN_5784;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h18 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_24 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_24 <= _GEN_5785;
      end
    end else begin
      rob_n_flits_24 <= _GEN_5785;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h19 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_25 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_25 <= _GEN_5786;
      end
    end else begin
      rob_n_flits_25 <= _GEN_5786;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1a == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_26 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_26 <= _GEN_5787;
      end
    end else begin
      rob_n_flits_26 <= _GEN_5787;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1b == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_27 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_27 <= _GEN_5788;
      end
    end else begin
      rob_n_flits_27 <= _GEN_5788;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1c == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_28 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_28 <= _GEN_5789;
      end
    end else begin
      rob_n_flits_28 <= _GEN_5789;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1d == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_29 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_29 <= _GEN_5790;
      end
    end else begin
      rob_n_flits_29 <= _GEN_5790;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1e == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_30 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_30 <= _GEN_5791;
      end
    end else begin
      rob_n_flits_30 <= _GEN_5791;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1f == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_31 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_31 <= _GEN_5792;
      end
    end else begin
      rob_n_flits_31 <= _GEN_5792;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h20 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_32 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_32 <= _GEN_5793;
      end
    end else begin
      rob_n_flits_32 <= _GEN_5793;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h21 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_33 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_33 <= _GEN_5794;
      end
    end else begin
      rob_n_flits_33 <= _GEN_5794;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h22 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_34 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_34 <= _GEN_5795;
      end
    end else begin
      rob_n_flits_34 <= _GEN_5795;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h23 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_35 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_35 <= _GEN_5796;
      end
    end else begin
      rob_n_flits_35 <= _GEN_5796;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h24 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_36 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_36 <= _GEN_5797;
      end
    end else begin
      rob_n_flits_36 <= _GEN_5797;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h25 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_37 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_37 <= _GEN_5798;
      end
    end else begin
      rob_n_flits_37 <= _GEN_5798;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h26 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_38 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_38 <= _GEN_5799;
      end
    end else begin
      rob_n_flits_38 <= _GEN_5799;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h27 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_39 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_39 <= _GEN_5800;
      end
    end else begin
      rob_n_flits_39 <= _GEN_5800;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h28 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_40 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_40 <= _GEN_5801;
      end
    end else begin
      rob_n_flits_40 <= _GEN_5801;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h29 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_41 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_41 <= _GEN_5802;
      end
    end else begin
      rob_n_flits_41 <= _GEN_5802;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2a == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_42 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_42 <= _GEN_5803;
      end
    end else begin
      rob_n_flits_42 <= _GEN_5803;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2b == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_43 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_43 <= _GEN_5804;
      end
    end else begin
      rob_n_flits_43 <= _GEN_5804;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2c == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_44 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_44 <= _GEN_5805;
      end
    end else begin
      rob_n_flits_44 <= _GEN_5805;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2d == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_45 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_45 <= _GEN_5806;
      end
    end else begin
      rob_n_flits_45 <= _GEN_5806;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2e == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_46 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_46 <= _GEN_5807;
      end
    end else begin
      rob_n_flits_46 <= _GEN_5807;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2f == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_47 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_47 <= _GEN_5808;
      end
    end else begin
      rob_n_flits_47 <= _GEN_5808;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h30 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_48 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_48 <= _GEN_5809;
      end
    end else begin
      rob_n_flits_48 <= _GEN_5809;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h31 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_49 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_49 <= _GEN_5810;
      end
    end else begin
      rob_n_flits_49 <= _GEN_5810;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h32 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_50 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_50 <= _GEN_5811;
      end
    end else begin
      rob_n_flits_50 <= _GEN_5811;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h33 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_51 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_51 <= _GEN_5812;
      end
    end else begin
      rob_n_flits_51 <= _GEN_5812;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h34 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_52 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_52 <= _GEN_5813;
      end
    end else begin
      rob_n_flits_52 <= _GEN_5813;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h35 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_53 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_53 <= _GEN_5814;
      end
    end else begin
      rob_n_flits_53 <= _GEN_5814;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h36 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_54 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_54 <= _GEN_5815;
      end
    end else begin
      rob_n_flits_54 <= _GEN_5815;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h37 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_55 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_55 <= _GEN_5816;
      end
    end else begin
      rob_n_flits_55 <= _GEN_5816;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h38 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_56 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_56 <= _GEN_5817;
      end
    end else begin
      rob_n_flits_56 <= _GEN_5817;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h39 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_57 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_57 <= _GEN_5818;
      end
    end else begin
      rob_n_flits_57 <= _GEN_5818;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3a == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_58 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_58 <= _GEN_5819;
      end
    end else begin
      rob_n_flits_58 <= _GEN_5819;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3b == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_59 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_59 <= _GEN_5820;
      end
    end else begin
      rob_n_flits_59 <= _GEN_5820;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3c == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_60 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_60 <= _GEN_5821;
      end
    end else begin
      rob_n_flits_60 <= _GEN_5821;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3d == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_61 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_61 <= _GEN_5822;
      end
    end else begin
      rob_n_flits_61 <= _GEN_5822;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3e == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_62 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_62 <= _GEN_5823;
      end
    end else begin
      rob_n_flits_62 <= _GEN_5823;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3f == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_63 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_63 <= _GEN_5824;
      end
    end else begin
      rob_n_flits_63 <= _GEN_5824;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h40 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_64 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_64 <= _GEN_5825;
      end
    end else begin
      rob_n_flits_64 <= _GEN_5825;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h41 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_65 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_65 <= _GEN_5826;
      end
    end else begin
      rob_n_flits_65 <= _GEN_5826;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h42 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_66 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_66 <= _GEN_5827;
      end
    end else begin
      rob_n_flits_66 <= _GEN_5827;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h43 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_67 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_67 <= _GEN_5828;
      end
    end else begin
      rob_n_flits_67 <= _GEN_5828;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h44 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_68 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_68 <= _GEN_5829;
      end
    end else begin
      rob_n_flits_68 <= _GEN_5829;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h45 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_69 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_69 <= _GEN_5830;
      end
    end else begin
      rob_n_flits_69 <= _GEN_5830;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h46 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_70 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_70 <= _GEN_5831;
      end
    end else begin
      rob_n_flits_70 <= _GEN_5831;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h47 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_71 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_71 <= _GEN_5832;
      end
    end else begin
      rob_n_flits_71 <= _GEN_5832;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h48 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_72 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_72 <= _GEN_5833;
      end
    end else begin
      rob_n_flits_72 <= _GEN_5833;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h49 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_73 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_73 <= _GEN_5834;
      end
    end else begin
      rob_n_flits_73 <= _GEN_5834;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4a == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_74 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_74 <= _GEN_5835;
      end
    end else begin
      rob_n_flits_74 <= _GEN_5835;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4b == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_75 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_75 <= _GEN_5836;
      end
    end else begin
      rob_n_flits_75 <= _GEN_5836;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4c == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_76 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_76 <= _GEN_5837;
      end
    end else begin
      rob_n_flits_76 <= _GEN_5837;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4d == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_77 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_77 <= _GEN_5838;
      end
    end else begin
      rob_n_flits_77 <= _GEN_5838;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4e == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_78 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_78 <= _GEN_5839;
      end
    end else begin
      rob_n_flits_78 <= _GEN_5839;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4f == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_79 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_79 <= _GEN_5840;
      end
    end else begin
      rob_n_flits_79 <= _GEN_5840;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h50 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_80 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_80 <= _GEN_5841;
      end
    end else begin
      rob_n_flits_80 <= _GEN_5841;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h51 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_81 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_81 <= _GEN_5842;
      end
    end else begin
      rob_n_flits_81 <= _GEN_5842;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h52 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_82 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_82 <= _GEN_5843;
      end
    end else begin
      rob_n_flits_82 <= _GEN_5843;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h53 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_83 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_83 <= _GEN_5844;
      end
    end else begin
      rob_n_flits_83 <= _GEN_5844;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h54 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_84 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_84 <= _GEN_5845;
      end
    end else begin
      rob_n_flits_84 <= _GEN_5845;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h55 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_85 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_85 <= _GEN_5846;
      end
    end else begin
      rob_n_flits_85 <= _GEN_5846;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h56 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_86 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_86 <= _GEN_5847;
      end
    end else begin
      rob_n_flits_86 <= _GEN_5847;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h57 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_87 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_87 <= _GEN_5848;
      end
    end else begin
      rob_n_flits_87 <= _GEN_5848;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h58 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_88 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_88 <= _GEN_5849;
      end
    end else begin
      rob_n_flits_88 <= _GEN_5849;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h59 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_89 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_89 <= _GEN_5850;
      end
    end else begin
      rob_n_flits_89 <= _GEN_5850;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5a == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_90 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_90 <= _GEN_5851;
      end
    end else begin
      rob_n_flits_90 <= _GEN_5851;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5b == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_91 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_91 <= _GEN_5852;
      end
    end else begin
      rob_n_flits_91 <= _GEN_5852;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5c == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_92 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_92 <= _GEN_5853;
      end
    end else begin
      rob_n_flits_92 <= _GEN_5853;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5d == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_93 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_93 <= _GEN_5854;
      end
    end else begin
      rob_n_flits_93 <= _GEN_5854;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5e == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_94 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_94 <= _GEN_5855;
      end
    end else begin
      rob_n_flits_94 <= _GEN_5855;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5f == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_95 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_95 <= _GEN_5856;
      end
    end else begin
      rob_n_flits_95 <= _GEN_5856;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h60 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_96 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_96 <= _GEN_5857;
      end
    end else begin
      rob_n_flits_96 <= _GEN_5857;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h61 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_97 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_97 <= _GEN_5858;
      end
    end else begin
      rob_n_flits_97 <= _GEN_5858;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h62 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_98 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_98 <= _GEN_5859;
      end
    end else begin
      rob_n_flits_98 <= _GEN_5859;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h63 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_99 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_99 <= _GEN_5860;
      end
    end else begin
      rob_n_flits_99 <= _GEN_5860;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h64 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_100 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_100 <= _GEN_5861;
      end
    end else begin
      rob_n_flits_100 <= _GEN_5861;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h65 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_101 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_101 <= _GEN_5862;
      end
    end else begin
      rob_n_flits_101 <= _GEN_5862;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h66 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_102 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_102 <= _GEN_5863;
      end
    end else begin
      rob_n_flits_102 <= _GEN_5863;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h67 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_103 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_103 <= _GEN_5864;
      end
    end else begin
      rob_n_flits_103 <= _GEN_5864;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h68 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_104 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_104 <= _GEN_5865;
      end
    end else begin
      rob_n_flits_104 <= _GEN_5865;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h69 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_105 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_105 <= _GEN_5866;
      end
    end else begin
      rob_n_flits_105 <= _GEN_5866;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6a == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_106 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_106 <= _GEN_5867;
      end
    end else begin
      rob_n_flits_106 <= _GEN_5867;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6b == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_107 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_107 <= _GEN_5868;
      end
    end else begin
      rob_n_flits_107 <= _GEN_5868;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6c == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_108 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_108 <= _GEN_5869;
      end
    end else begin
      rob_n_flits_108 <= _GEN_5869;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6d == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_109 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_109 <= _GEN_5870;
      end
    end else begin
      rob_n_flits_109 <= _GEN_5870;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6e == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_110 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_110 <= _GEN_5871;
      end
    end else begin
      rob_n_flits_110 <= _GEN_5871;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6f == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_111 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_111 <= _GEN_5872;
      end
    end else begin
      rob_n_flits_111 <= _GEN_5872;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h70 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_112 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_112 <= _GEN_5873;
      end
    end else begin
      rob_n_flits_112 <= _GEN_5873;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h71 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_113 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_113 <= _GEN_5874;
      end
    end else begin
      rob_n_flits_113 <= _GEN_5874;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h72 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_114 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_114 <= _GEN_5875;
      end
    end else begin
      rob_n_flits_114 <= _GEN_5875;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h73 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_115 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_115 <= _GEN_5876;
      end
    end else begin
      rob_n_flits_115 <= _GEN_5876;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h74 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_116 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_116 <= _GEN_5877;
      end
    end else begin
      rob_n_flits_116 <= _GEN_5877;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h75 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_117 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_117 <= _GEN_5878;
      end
    end else begin
      rob_n_flits_117 <= _GEN_5878;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h76 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_118 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_118 <= _GEN_5879;
      end
    end else begin
      rob_n_flits_118 <= _GEN_5879;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h77 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_119 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_119 <= _GEN_5880;
      end
    end else begin
      rob_n_flits_119 <= _GEN_5880;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h78 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_120 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_120 <= _GEN_5881;
      end
    end else begin
      rob_n_flits_120 <= _GEN_5881;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h79 == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_121 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_121 <= _GEN_5882;
      end
    end else begin
      rob_n_flits_121 <= _GEN_5882;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7a == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_122 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_122 <= _GEN_5883;
      end
    end else begin
      rob_n_flits_122 <= _GEN_5883;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7b == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_123 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_123 <= _GEN_5884;
      end
    end else begin
      rob_n_flits_123 <= _GEN_5884;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7c == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_124 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_124 <= _GEN_5885;
      end
    end else begin
      rob_n_flits_124 <= _GEN_5885;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7d == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_125 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_125 <= _GEN_5886;
      end
    end else begin
      rob_n_flits_125 <= _GEN_5886;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7e == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_126 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_126 <= _GEN_5887;
      end
    end else begin
      rob_n_flits_126 <= _GEN_5887;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7f == rob_alloc_ids_3) begin // @[TestHarness.scala 182:36]
        rob_n_flits_127 <= _rob_n_flits_T_69; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_127 <= _GEN_5888;
      end
    end else begin
      rob_n_flits_127 <= _GEN_5888;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h0 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_0 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_0 <= _GEN_13326;
      end
    end else begin
      rob_flits_returned_0 <= _GEN_13326;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h1 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_1 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_1 <= _GEN_13327;
      end
    end else begin
      rob_flits_returned_1 <= _GEN_13327;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h2 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_2 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_2 <= _GEN_13328;
      end
    end else begin
      rob_flits_returned_2 <= _GEN_13328;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h3 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_3 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_3 <= _GEN_13329;
      end
    end else begin
      rob_flits_returned_3 <= _GEN_13329;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h4 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_4 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_4 <= _GEN_13330;
      end
    end else begin
      rob_flits_returned_4 <= _GEN_13330;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h5 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_5 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_5 <= _GEN_13331;
      end
    end else begin
      rob_flits_returned_5 <= _GEN_13331;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h6 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_6 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_6 <= _GEN_13332;
      end
    end else begin
      rob_flits_returned_6 <= _GEN_13332;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h7 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_7 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_7 <= _GEN_13333;
      end
    end else begin
      rob_flits_returned_7 <= _GEN_13333;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h8 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_8 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_8 <= _GEN_13334;
      end
    end else begin
      rob_flits_returned_8 <= _GEN_13334;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h9 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_9 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_9 <= _GEN_13335;
      end
    end else begin
      rob_flits_returned_9 <= _GEN_13335;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'ha == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_10 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_10 <= _GEN_13336;
      end
    end else begin
      rob_flits_returned_10 <= _GEN_13336;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'hb == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_11 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_11 <= _GEN_13337;
      end
    end else begin
      rob_flits_returned_11 <= _GEN_13337;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'hc == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_12 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_12 <= _GEN_13338;
      end
    end else begin
      rob_flits_returned_12 <= _GEN_13338;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'hd == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_13 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_13 <= _GEN_13339;
      end
    end else begin
      rob_flits_returned_13 <= _GEN_13339;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'he == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_14 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_14 <= _GEN_13340;
      end
    end else begin
      rob_flits_returned_14 <= _GEN_13340;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'hf == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_15 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_15 <= _GEN_13341;
      end
    end else begin
      rob_flits_returned_15 <= _GEN_13341;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h10 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_16 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_16 <= _GEN_13342;
      end
    end else begin
      rob_flits_returned_16 <= _GEN_13342;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h11 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_17 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_17 <= _GEN_13343;
      end
    end else begin
      rob_flits_returned_17 <= _GEN_13343;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h12 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_18 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_18 <= _GEN_13344;
      end
    end else begin
      rob_flits_returned_18 <= _GEN_13344;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h13 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_19 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_19 <= _GEN_13345;
      end
    end else begin
      rob_flits_returned_19 <= _GEN_13345;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h14 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_20 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_20 <= _GEN_13346;
      end
    end else begin
      rob_flits_returned_20 <= _GEN_13346;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h15 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_21 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_21 <= _GEN_13347;
      end
    end else begin
      rob_flits_returned_21 <= _GEN_13347;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h16 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_22 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_22 <= _GEN_13348;
      end
    end else begin
      rob_flits_returned_22 <= _GEN_13348;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h17 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_23 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_23 <= _GEN_13349;
      end
    end else begin
      rob_flits_returned_23 <= _GEN_13349;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h18 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_24 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_24 <= _GEN_13350;
      end
    end else begin
      rob_flits_returned_24 <= _GEN_13350;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h19 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_25 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_25 <= _GEN_13351;
      end
    end else begin
      rob_flits_returned_25 <= _GEN_13351;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h1a == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_26 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_26 <= _GEN_13352;
      end
    end else begin
      rob_flits_returned_26 <= _GEN_13352;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h1b == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_27 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_27 <= _GEN_13353;
      end
    end else begin
      rob_flits_returned_27 <= _GEN_13353;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h1c == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_28 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_28 <= _GEN_13354;
      end
    end else begin
      rob_flits_returned_28 <= _GEN_13354;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h1d == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_29 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_29 <= _GEN_13355;
      end
    end else begin
      rob_flits_returned_29 <= _GEN_13355;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h1e == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_30 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_30 <= _GEN_13356;
      end
    end else begin
      rob_flits_returned_30 <= _GEN_13356;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h1f == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_31 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_31 <= _GEN_13357;
      end
    end else begin
      rob_flits_returned_31 <= _GEN_13357;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h20 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_32 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_32 <= _GEN_13358;
      end
    end else begin
      rob_flits_returned_32 <= _GEN_13358;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h21 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_33 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_33 <= _GEN_13359;
      end
    end else begin
      rob_flits_returned_33 <= _GEN_13359;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h22 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_34 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_34 <= _GEN_13360;
      end
    end else begin
      rob_flits_returned_34 <= _GEN_13360;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h23 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_35 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_35 <= _GEN_13361;
      end
    end else begin
      rob_flits_returned_35 <= _GEN_13361;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h24 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_36 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_36 <= _GEN_13362;
      end
    end else begin
      rob_flits_returned_36 <= _GEN_13362;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h25 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_37 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_37 <= _GEN_13363;
      end
    end else begin
      rob_flits_returned_37 <= _GEN_13363;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h26 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_38 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_38 <= _GEN_13364;
      end
    end else begin
      rob_flits_returned_38 <= _GEN_13364;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h27 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_39 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_39 <= _GEN_13365;
      end
    end else begin
      rob_flits_returned_39 <= _GEN_13365;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h28 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_40 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_40 <= _GEN_13366;
      end
    end else begin
      rob_flits_returned_40 <= _GEN_13366;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h29 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_41 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_41 <= _GEN_13367;
      end
    end else begin
      rob_flits_returned_41 <= _GEN_13367;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h2a == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_42 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_42 <= _GEN_13368;
      end
    end else begin
      rob_flits_returned_42 <= _GEN_13368;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h2b == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_43 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_43 <= _GEN_13369;
      end
    end else begin
      rob_flits_returned_43 <= _GEN_13369;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h2c == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_44 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_44 <= _GEN_13370;
      end
    end else begin
      rob_flits_returned_44 <= _GEN_13370;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h2d == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_45 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_45 <= _GEN_13371;
      end
    end else begin
      rob_flits_returned_45 <= _GEN_13371;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h2e == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_46 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_46 <= _GEN_13372;
      end
    end else begin
      rob_flits_returned_46 <= _GEN_13372;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h2f == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_47 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_47 <= _GEN_13373;
      end
    end else begin
      rob_flits_returned_47 <= _GEN_13373;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h30 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_48 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_48 <= _GEN_13374;
      end
    end else begin
      rob_flits_returned_48 <= _GEN_13374;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h31 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_49 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_49 <= _GEN_13375;
      end
    end else begin
      rob_flits_returned_49 <= _GEN_13375;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h32 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_50 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_50 <= _GEN_13376;
      end
    end else begin
      rob_flits_returned_50 <= _GEN_13376;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h33 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_51 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_51 <= _GEN_13377;
      end
    end else begin
      rob_flits_returned_51 <= _GEN_13377;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h34 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_52 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_52 <= _GEN_13378;
      end
    end else begin
      rob_flits_returned_52 <= _GEN_13378;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h35 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_53 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_53 <= _GEN_13379;
      end
    end else begin
      rob_flits_returned_53 <= _GEN_13379;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h36 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_54 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_54 <= _GEN_13380;
      end
    end else begin
      rob_flits_returned_54 <= _GEN_13380;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h37 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_55 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_55 <= _GEN_13381;
      end
    end else begin
      rob_flits_returned_55 <= _GEN_13381;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h38 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_56 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_56 <= _GEN_13382;
      end
    end else begin
      rob_flits_returned_56 <= _GEN_13382;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h39 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_57 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_57 <= _GEN_13383;
      end
    end else begin
      rob_flits_returned_57 <= _GEN_13383;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h3a == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_58 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_58 <= _GEN_13384;
      end
    end else begin
      rob_flits_returned_58 <= _GEN_13384;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h3b == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_59 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_59 <= _GEN_13385;
      end
    end else begin
      rob_flits_returned_59 <= _GEN_13385;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h3c == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_60 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_60 <= _GEN_13386;
      end
    end else begin
      rob_flits_returned_60 <= _GEN_13386;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h3d == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_61 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_61 <= _GEN_13387;
      end
    end else begin
      rob_flits_returned_61 <= _GEN_13387;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h3e == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_62 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_62 <= _GEN_13388;
      end
    end else begin
      rob_flits_returned_62 <= _GEN_13388;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h3f == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_63 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_63 <= _GEN_13389;
      end
    end else begin
      rob_flits_returned_63 <= _GEN_13389;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h40 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_64 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_64 <= _GEN_13390;
      end
    end else begin
      rob_flits_returned_64 <= _GEN_13390;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h41 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_65 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_65 <= _GEN_13391;
      end
    end else begin
      rob_flits_returned_65 <= _GEN_13391;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h42 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_66 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_66 <= _GEN_13392;
      end
    end else begin
      rob_flits_returned_66 <= _GEN_13392;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h43 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_67 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_67 <= _GEN_13393;
      end
    end else begin
      rob_flits_returned_67 <= _GEN_13393;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h44 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_68 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_68 <= _GEN_13394;
      end
    end else begin
      rob_flits_returned_68 <= _GEN_13394;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h45 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_69 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_69 <= _GEN_13395;
      end
    end else begin
      rob_flits_returned_69 <= _GEN_13395;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h46 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_70 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_70 <= _GEN_13396;
      end
    end else begin
      rob_flits_returned_70 <= _GEN_13396;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h47 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_71 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_71 <= _GEN_13397;
      end
    end else begin
      rob_flits_returned_71 <= _GEN_13397;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h48 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_72 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_72 <= _GEN_13398;
      end
    end else begin
      rob_flits_returned_72 <= _GEN_13398;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h49 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_73 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_73 <= _GEN_13399;
      end
    end else begin
      rob_flits_returned_73 <= _GEN_13399;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h4a == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_74 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_74 <= _GEN_13400;
      end
    end else begin
      rob_flits_returned_74 <= _GEN_13400;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h4b == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_75 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_75 <= _GEN_13401;
      end
    end else begin
      rob_flits_returned_75 <= _GEN_13401;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h4c == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_76 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_76 <= _GEN_13402;
      end
    end else begin
      rob_flits_returned_76 <= _GEN_13402;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h4d == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_77 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_77 <= _GEN_13403;
      end
    end else begin
      rob_flits_returned_77 <= _GEN_13403;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h4e == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_78 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_78 <= _GEN_13404;
      end
    end else begin
      rob_flits_returned_78 <= _GEN_13404;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h4f == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_79 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_79 <= _GEN_13405;
      end
    end else begin
      rob_flits_returned_79 <= _GEN_13405;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h50 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_80 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_80 <= _GEN_13406;
      end
    end else begin
      rob_flits_returned_80 <= _GEN_13406;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h51 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_81 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_81 <= _GEN_13407;
      end
    end else begin
      rob_flits_returned_81 <= _GEN_13407;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h52 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_82 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_82 <= _GEN_13408;
      end
    end else begin
      rob_flits_returned_82 <= _GEN_13408;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h53 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_83 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_83 <= _GEN_13409;
      end
    end else begin
      rob_flits_returned_83 <= _GEN_13409;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h54 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_84 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_84 <= _GEN_13410;
      end
    end else begin
      rob_flits_returned_84 <= _GEN_13410;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h55 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_85 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_85 <= _GEN_13411;
      end
    end else begin
      rob_flits_returned_85 <= _GEN_13411;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h56 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_86 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_86 <= _GEN_13412;
      end
    end else begin
      rob_flits_returned_86 <= _GEN_13412;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h57 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_87 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_87 <= _GEN_13413;
      end
    end else begin
      rob_flits_returned_87 <= _GEN_13413;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h58 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_88 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_88 <= _GEN_13414;
      end
    end else begin
      rob_flits_returned_88 <= _GEN_13414;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h59 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_89 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_89 <= _GEN_13415;
      end
    end else begin
      rob_flits_returned_89 <= _GEN_13415;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h5a == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_90 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_90 <= _GEN_13416;
      end
    end else begin
      rob_flits_returned_90 <= _GEN_13416;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h5b == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_91 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_91 <= _GEN_13417;
      end
    end else begin
      rob_flits_returned_91 <= _GEN_13417;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h5c == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_92 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_92 <= _GEN_13418;
      end
    end else begin
      rob_flits_returned_92 <= _GEN_13418;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h5d == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_93 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_93 <= _GEN_13419;
      end
    end else begin
      rob_flits_returned_93 <= _GEN_13419;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h5e == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_94 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_94 <= _GEN_13420;
      end
    end else begin
      rob_flits_returned_94 <= _GEN_13420;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h5f == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_95 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_95 <= _GEN_13421;
      end
    end else begin
      rob_flits_returned_95 <= _GEN_13421;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h60 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_96 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_96 <= _GEN_13422;
      end
    end else begin
      rob_flits_returned_96 <= _GEN_13422;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h61 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_97 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_97 <= _GEN_13423;
      end
    end else begin
      rob_flits_returned_97 <= _GEN_13423;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h62 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_98 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_98 <= _GEN_13424;
      end
    end else begin
      rob_flits_returned_98 <= _GEN_13424;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h63 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_99 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_99 <= _GEN_13425;
      end
    end else begin
      rob_flits_returned_99 <= _GEN_13425;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h64 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_100 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_100 <= _GEN_13426;
      end
    end else begin
      rob_flits_returned_100 <= _GEN_13426;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h65 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_101 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_101 <= _GEN_13427;
      end
    end else begin
      rob_flits_returned_101 <= _GEN_13427;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h66 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_102 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_102 <= _GEN_13428;
      end
    end else begin
      rob_flits_returned_102 <= _GEN_13428;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h67 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_103 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_103 <= _GEN_13429;
      end
    end else begin
      rob_flits_returned_103 <= _GEN_13429;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h68 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_104 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_104 <= _GEN_13430;
      end
    end else begin
      rob_flits_returned_104 <= _GEN_13430;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h69 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_105 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_105 <= _GEN_13431;
      end
    end else begin
      rob_flits_returned_105 <= _GEN_13431;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h6a == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_106 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_106 <= _GEN_13432;
      end
    end else begin
      rob_flits_returned_106 <= _GEN_13432;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h6b == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_107 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_107 <= _GEN_13433;
      end
    end else begin
      rob_flits_returned_107 <= _GEN_13433;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h6c == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_108 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_108 <= _GEN_13434;
      end
    end else begin
      rob_flits_returned_108 <= _GEN_13434;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h6d == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_109 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_109 <= _GEN_13435;
      end
    end else begin
      rob_flits_returned_109 <= _GEN_13435;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h6e == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_110 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_110 <= _GEN_13436;
      end
    end else begin
      rob_flits_returned_110 <= _GEN_13436;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h6f == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_111 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_111 <= _GEN_13437;
      end
    end else begin
      rob_flits_returned_111 <= _GEN_13437;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h70 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_112 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_112 <= _GEN_13438;
      end
    end else begin
      rob_flits_returned_112 <= _GEN_13438;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h71 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_113 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_113 <= _GEN_13439;
      end
    end else begin
      rob_flits_returned_113 <= _GEN_13439;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h72 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_114 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_114 <= _GEN_13440;
      end
    end else begin
      rob_flits_returned_114 <= _GEN_13440;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h73 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_115 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_115 <= _GEN_13441;
      end
    end else begin
      rob_flits_returned_115 <= _GEN_13441;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h74 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_116 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_116 <= _GEN_13442;
      end
    end else begin
      rob_flits_returned_116 <= _GEN_13442;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h75 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_117 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_117 <= _GEN_13443;
      end
    end else begin
      rob_flits_returned_117 <= _GEN_13443;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h76 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_118 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_118 <= _GEN_13444;
      end
    end else begin
      rob_flits_returned_118 <= _GEN_13444;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h77 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_119 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_119 <= _GEN_13445;
      end
    end else begin
      rob_flits_returned_119 <= _GEN_13445;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h78 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_120 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_120 <= _GEN_13446;
      end
    end else begin
      rob_flits_returned_120 <= _GEN_13446;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h79 == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_121 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_121 <= _GEN_13447;
      end
    end else begin
      rob_flits_returned_121 <= _GEN_13447;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h7a == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_122 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_122 <= _GEN_13448;
      end
    end else begin
      rob_flits_returned_122 <= _GEN_13448;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h7b == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_123 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_123 <= _GEN_13449;
      end
    end else begin
      rob_flits_returned_123 <= _GEN_13449;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h7c == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_124 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_124 <= _GEN_13450;
      end
    end else begin
      rob_flits_returned_124 <= _GEN_13450;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h7d == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_125 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_125 <= _GEN_13451;
      end
    end else begin
      rob_flits_returned_125 <= _GEN_13451;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h7e == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_126 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_126 <= _GEN_13452;
      end
    end else begin
      rob_flits_returned_126 <= _GEN_13452;
    end
    if (_T_259) begin // @[TestHarness.scala 199:26]
      if (7'h7f == out_payload_3_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_127 <= _rob_flits_returned_T_11; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_127 <= _GEN_13453;
      end
    end else begin
      rob_flits_returned_127 <= _GEN_13453;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h0 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_0 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_0 <= _GEN_6017;
      end
    end else begin
      rob_tscs_0 <= _GEN_6017;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_1 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_1 <= _GEN_6018;
      end
    end else begin
      rob_tscs_1 <= _GEN_6018;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_2 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_2 <= _GEN_6019;
      end
    end else begin
      rob_tscs_2 <= _GEN_6019;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_3 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_3 <= _GEN_6020;
      end
    end else begin
      rob_tscs_3 <= _GEN_6020;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_4 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_4 <= _GEN_6021;
      end
    end else begin
      rob_tscs_4 <= _GEN_6021;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_5 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_5 <= _GEN_6022;
      end
    end else begin
      rob_tscs_5 <= _GEN_6022;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_6 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_6 <= _GEN_6023;
      end
    end else begin
      rob_tscs_6 <= _GEN_6023;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_7 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_7 <= _GEN_6024;
      end
    end else begin
      rob_tscs_7 <= _GEN_6024;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h8 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_8 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_8 <= _GEN_6025;
      end
    end else begin
      rob_tscs_8 <= _GEN_6025;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h9 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_9 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_9 <= _GEN_6026;
      end
    end else begin
      rob_tscs_9 <= _GEN_6026;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'ha == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_10 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_10 <= _GEN_6027;
      end
    end else begin
      rob_tscs_10 <= _GEN_6027;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hb == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_11 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_11 <= _GEN_6028;
      end
    end else begin
      rob_tscs_11 <= _GEN_6028;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hc == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_12 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_12 <= _GEN_6029;
      end
    end else begin
      rob_tscs_12 <= _GEN_6029;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hd == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_13 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_13 <= _GEN_6030;
      end
    end else begin
      rob_tscs_13 <= _GEN_6030;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'he == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_14 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_14 <= _GEN_6031;
      end
    end else begin
      rob_tscs_14 <= _GEN_6031;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hf == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_15 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_15 <= _GEN_6032;
      end
    end else begin
      rob_tscs_15 <= _GEN_6032;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h10 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_16 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_16 <= _GEN_6033;
      end
    end else begin
      rob_tscs_16 <= _GEN_6033;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h11 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_17 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_17 <= _GEN_6034;
      end
    end else begin
      rob_tscs_17 <= _GEN_6034;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h12 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_18 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_18 <= _GEN_6035;
      end
    end else begin
      rob_tscs_18 <= _GEN_6035;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h13 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_19 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_19 <= _GEN_6036;
      end
    end else begin
      rob_tscs_19 <= _GEN_6036;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h14 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_20 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_20 <= _GEN_6037;
      end
    end else begin
      rob_tscs_20 <= _GEN_6037;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h15 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_21 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_21 <= _GEN_6038;
      end
    end else begin
      rob_tscs_21 <= _GEN_6038;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h16 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_22 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_22 <= _GEN_6039;
      end
    end else begin
      rob_tscs_22 <= _GEN_6039;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h17 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_23 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_23 <= _GEN_6040;
      end
    end else begin
      rob_tscs_23 <= _GEN_6040;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h18 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_24 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_24 <= _GEN_6041;
      end
    end else begin
      rob_tscs_24 <= _GEN_6041;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h19 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_25 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_25 <= _GEN_6042;
      end
    end else begin
      rob_tscs_25 <= _GEN_6042;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1a == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_26 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_26 <= _GEN_6043;
      end
    end else begin
      rob_tscs_26 <= _GEN_6043;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1b == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_27 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_27 <= _GEN_6044;
      end
    end else begin
      rob_tscs_27 <= _GEN_6044;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1c == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_28 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_28 <= _GEN_6045;
      end
    end else begin
      rob_tscs_28 <= _GEN_6045;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1d == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_29 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_29 <= _GEN_6046;
      end
    end else begin
      rob_tscs_29 <= _GEN_6046;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1e == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_30 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_30 <= _GEN_6047;
      end
    end else begin
      rob_tscs_30 <= _GEN_6047;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1f == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_31 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_31 <= _GEN_6048;
      end
    end else begin
      rob_tscs_31 <= _GEN_6048;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h20 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_32 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_32 <= _GEN_6049;
      end
    end else begin
      rob_tscs_32 <= _GEN_6049;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h21 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_33 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_33 <= _GEN_6050;
      end
    end else begin
      rob_tscs_33 <= _GEN_6050;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h22 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_34 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_34 <= _GEN_6051;
      end
    end else begin
      rob_tscs_34 <= _GEN_6051;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h23 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_35 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_35 <= _GEN_6052;
      end
    end else begin
      rob_tscs_35 <= _GEN_6052;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h24 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_36 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_36 <= _GEN_6053;
      end
    end else begin
      rob_tscs_36 <= _GEN_6053;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h25 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_37 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_37 <= _GEN_6054;
      end
    end else begin
      rob_tscs_37 <= _GEN_6054;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h26 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_38 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_38 <= _GEN_6055;
      end
    end else begin
      rob_tscs_38 <= _GEN_6055;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h27 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_39 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_39 <= _GEN_6056;
      end
    end else begin
      rob_tscs_39 <= _GEN_6056;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h28 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_40 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_40 <= _GEN_6057;
      end
    end else begin
      rob_tscs_40 <= _GEN_6057;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h29 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_41 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_41 <= _GEN_6058;
      end
    end else begin
      rob_tscs_41 <= _GEN_6058;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2a == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_42 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_42 <= _GEN_6059;
      end
    end else begin
      rob_tscs_42 <= _GEN_6059;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2b == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_43 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_43 <= _GEN_6060;
      end
    end else begin
      rob_tscs_43 <= _GEN_6060;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2c == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_44 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_44 <= _GEN_6061;
      end
    end else begin
      rob_tscs_44 <= _GEN_6061;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2d == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_45 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_45 <= _GEN_6062;
      end
    end else begin
      rob_tscs_45 <= _GEN_6062;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2e == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_46 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_46 <= _GEN_6063;
      end
    end else begin
      rob_tscs_46 <= _GEN_6063;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2f == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_47 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_47 <= _GEN_6064;
      end
    end else begin
      rob_tscs_47 <= _GEN_6064;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h30 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_48 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_48 <= _GEN_6065;
      end
    end else begin
      rob_tscs_48 <= _GEN_6065;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h31 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_49 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_49 <= _GEN_6066;
      end
    end else begin
      rob_tscs_49 <= _GEN_6066;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h32 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_50 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_50 <= _GEN_6067;
      end
    end else begin
      rob_tscs_50 <= _GEN_6067;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h33 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_51 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_51 <= _GEN_6068;
      end
    end else begin
      rob_tscs_51 <= _GEN_6068;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h34 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_52 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_52 <= _GEN_6069;
      end
    end else begin
      rob_tscs_52 <= _GEN_6069;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h35 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_53 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_53 <= _GEN_6070;
      end
    end else begin
      rob_tscs_53 <= _GEN_6070;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h36 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_54 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_54 <= _GEN_6071;
      end
    end else begin
      rob_tscs_54 <= _GEN_6071;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h37 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_55 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_55 <= _GEN_6072;
      end
    end else begin
      rob_tscs_55 <= _GEN_6072;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h38 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_56 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_56 <= _GEN_6073;
      end
    end else begin
      rob_tscs_56 <= _GEN_6073;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h39 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_57 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_57 <= _GEN_6074;
      end
    end else begin
      rob_tscs_57 <= _GEN_6074;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3a == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_58 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_58 <= _GEN_6075;
      end
    end else begin
      rob_tscs_58 <= _GEN_6075;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3b == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_59 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_59 <= _GEN_6076;
      end
    end else begin
      rob_tscs_59 <= _GEN_6076;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3c == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_60 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_60 <= _GEN_6077;
      end
    end else begin
      rob_tscs_60 <= _GEN_6077;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3d == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_61 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_61 <= _GEN_6078;
      end
    end else begin
      rob_tscs_61 <= _GEN_6078;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3e == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_62 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_62 <= _GEN_6079;
      end
    end else begin
      rob_tscs_62 <= _GEN_6079;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3f == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_63 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_63 <= _GEN_6080;
      end
    end else begin
      rob_tscs_63 <= _GEN_6080;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h40 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_64 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_64 <= _GEN_6081;
      end
    end else begin
      rob_tscs_64 <= _GEN_6081;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h41 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_65 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_65 <= _GEN_6082;
      end
    end else begin
      rob_tscs_65 <= _GEN_6082;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h42 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_66 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_66 <= _GEN_6083;
      end
    end else begin
      rob_tscs_66 <= _GEN_6083;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h43 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_67 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_67 <= _GEN_6084;
      end
    end else begin
      rob_tscs_67 <= _GEN_6084;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h44 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_68 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_68 <= _GEN_6085;
      end
    end else begin
      rob_tscs_68 <= _GEN_6085;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h45 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_69 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_69 <= _GEN_6086;
      end
    end else begin
      rob_tscs_69 <= _GEN_6086;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h46 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_70 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_70 <= _GEN_6087;
      end
    end else begin
      rob_tscs_70 <= _GEN_6087;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h47 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_71 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_71 <= _GEN_6088;
      end
    end else begin
      rob_tscs_71 <= _GEN_6088;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h48 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_72 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_72 <= _GEN_6089;
      end
    end else begin
      rob_tscs_72 <= _GEN_6089;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h49 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_73 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_73 <= _GEN_6090;
      end
    end else begin
      rob_tscs_73 <= _GEN_6090;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4a == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_74 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_74 <= _GEN_6091;
      end
    end else begin
      rob_tscs_74 <= _GEN_6091;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4b == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_75 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_75 <= _GEN_6092;
      end
    end else begin
      rob_tscs_75 <= _GEN_6092;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4c == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_76 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_76 <= _GEN_6093;
      end
    end else begin
      rob_tscs_76 <= _GEN_6093;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4d == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_77 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_77 <= _GEN_6094;
      end
    end else begin
      rob_tscs_77 <= _GEN_6094;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4e == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_78 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_78 <= _GEN_6095;
      end
    end else begin
      rob_tscs_78 <= _GEN_6095;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4f == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_79 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_79 <= _GEN_6096;
      end
    end else begin
      rob_tscs_79 <= _GEN_6096;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h50 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_80 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_80 <= _GEN_6097;
      end
    end else begin
      rob_tscs_80 <= _GEN_6097;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h51 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_81 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_81 <= _GEN_6098;
      end
    end else begin
      rob_tscs_81 <= _GEN_6098;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h52 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_82 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_82 <= _GEN_6099;
      end
    end else begin
      rob_tscs_82 <= _GEN_6099;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h53 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_83 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_83 <= _GEN_6100;
      end
    end else begin
      rob_tscs_83 <= _GEN_6100;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h54 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_84 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_84 <= _GEN_6101;
      end
    end else begin
      rob_tscs_84 <= _GEN_6101;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h55 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_85 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_85 <= _GEN_6102;
      end
    end else begin
      rob_tscs_85 <= _GEN_6102;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h56 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_86 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_86 <= _GEN_6103;
      end
    end else begin
      rob_tscs_86 <= _GEN_6103;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h57 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_87 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_87 <= _GEN_6104;
      end
    end else begin
      rob_tscs_87 <= _GEN_6104;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h58 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_88 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_88 <= _GEN_6105;
      end
    end else begin
      rob_tscs_88 <= _GEN_6105;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h59 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_89 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_89 <= _GEN_6106;
      end
    end else begin
      rob_tscs_89 <= _GEN_6106;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5a == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_90 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_90 <= _GEN_6107;
      end
    end else begin
      rob_tscs_90 <= _GEN_6107;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5b == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_91 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_91 <= _GEN_6108;
      end
    end else begin
      rob_tscs_91 <= _GEN_6108;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5c == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_92 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_92 <= _GEN_6109;
      end
    end else begin
      rob_tscs_92 <= _GEN_6109;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5d == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_93 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_93 <= _GEN_6110;
      end
    end else begin
      rob_tscs_93 <= _GEN_6110;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5e == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_94 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_94 <= _GEN_6111;
      end
    end else begin
      rob_tscs_94 <= _GEN_6111;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5f == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_95 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_95 <= _GEN_6112;
      end
    end else begin
      rob_tscs_95 <= _GEN_6112;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h60 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_96 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_96 <= _GEN_6113;
      end
    end else begin
      rob_tscs_96 <= _GEN_6113;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h61 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_97 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_97 <= _GEN_6114;
      end
    end else begin
      rob_tscs_97 <= _GEN_6114;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h62 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_98 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_98 <= _GEN_6115;
      end
    end else begin
      rob_tscs_98 <= _GEN_6115;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h63 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_99 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_99 <= _GEN_6116;
      end
    end else begin
      rob_tscs_99 <= _GEN_6116;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h64 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_100 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_100 <= _GEN_6117;
      end
    end else begin
      rob_tscs_100 <= _GEN_6117;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h65 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_101 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_101 <= _GEN_6118;
      end
    end else begin
      rob_tscs_101 <= _GEN_6118;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h66 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_102 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_102 <= _GEN_6119;
      end
    end else begin
      rob_tscs_102 <= _GEN_6119;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h67 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_103 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_103 <= _GEN_6120;
      end
    end else begin
      rob_tscs_103 <= _GEN_6120;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h68 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_104 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_104 <= _GEN_6121;
      end
    end else begin
      rob_tscs_104 <= _GEN_6121;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h69 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_105 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_105 <= _GEN_6122;
      end
    end else begin
      rob_tscs_105 <= _GEN_6122;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6a == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_106 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_106 <= _GEN_6123;
      end
    end else begin
      rob_tscs_106 <= _GEN_6123;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6b == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_107 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_107 <= _GEN_6124;
      end
    end else begin
      rob_tscs_107 <= _GEN_6124;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6c == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_108 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_108 <= _GEN_6125;
      end
    end else begin
      rob_tscs_108 <= _GEN_6125;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6d == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_109 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_109 <= _GEN_6126;
      end
    end else begin
      rob_tscs_109 <= _GEN_6126;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6e == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_110 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_110 <= _GEN_6127;
      end
    end else begin
      rob_tscs_110 <= _GEN_6127;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6f == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_111 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_111 <= _GEN_6128;
      end
    end else begin
      rob_tscs_111 <= _GEN_6128;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h70 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_112 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_112 <= _GEN_6129;
      end
    end else begin
      rob_tscs_112 <= _GEN_6129;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h71 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_113 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_113 <= _GEN_6130;
      end
    end else begin
      rob_tscs_113 <= _GEN_6130;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h72 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_114 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_114 <= _GEN_6131;
      end
    end else begin
      rob_tscs_114 <= _GEN_6131;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h73 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_115 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_115 <= _GEN_6132;
      end
    end else begin
      rob_tscs_115 <= _GEN_6132;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h74 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_116 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_116 <= _GEN_6133;
      end
    end else begin
      rob_tscs_116 <= _GEN_6133;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h75 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_117 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_117 <= _GEN_6134;
      end
    end else begin
      rob_tscs_117 <= _GEN_6134;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h76 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_118 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_118 <= _GEN_6135;
      end
    end else begin
      rob_tscs_118 <= _GEN_6135;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h77 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_119 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_119 <= _GEN_6136;
      end
    end else begin
      rob_tscs_119 <= _GEN_6136;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h78 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_120 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_120 <= _GEN_6137;
      end
    end else begin
      rob_tscs_120 <= _GEN_6137;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h79 == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_121 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_121 <= _GEN_6138;
      end
    end else begin
      rob_tscs_121 <= _GEN_6138;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7a == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_122 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_122 <= _GEN_6139;
      end
    end else begin
      rob_tscs_122 <= _GEN_6139;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7b == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_123 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_123 <= _GEN_6140;
      end
    end else begin
      rob_tscs_123 <= _GEN_6140;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7c == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_124 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_124 <= _GEN_6141;
      end
    end else begin
      rob_tscs_124 <= _GEN_6141;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7d == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_125 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_125 <= _GEN_6142;
      end
    end else begin
      rob_tscs_125 <= _GEN_6142;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7e == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_126 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_126 <= _GEN_6143;
      end
    end else begin
      rob_tscs_126 <= _GEN_6143;
    end
    if (igen_3_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7f == rob_alloc_ids_3) begin // @[TestHarness.scala 184:36]
        rob_tscs_127 <= _rob_tscs_T_31; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_127 <= _GEN_6144;
      end
    end else begin
      rob_tscs_127 <= _GEN_6144;
    end
    if (reset) begin // @[TestHarness.scala 164:24]
      io_success_REG <= 1'h0; // @[TestHarness.scala 164:24]
    end else begin
      io_success_REG <= success; // @[TestHarness.scala 164:24]
    end
    if (reset) begin // @[TestHarness.scala 196:31]
      packet_valid <= 1'h0; // @[TestHarness.scala 196:31]
    end else if (_T_118) begin // @[TestHarness.scala 199:26]
      if (io_from_noc_0_flit_bits_tail) begin // @[TestHarness.scala 216:31]
        packet_valid <= 1'h0; // @[TestHarness.scala 216:46]
      end else begin
        packet_valid <= _GEN_9729;
      end
    end
    packet_rob_idx <= _GEN_9989[6:0];
    if (reset) begin // @[TestHarness.scala 196:31]
      packet_valid_1 <= 1'h0; // @[TestHarness.scala 196:31]
    end else if (_T_165) begin // @[TestHarness.scala 199:26]
      if (io_from_noc_1_flit_bits_tail) begin // @[TestHarness.scala 216:31]
        packet_valid_1 <= 1'h0; // @[TestHarness.scala 216:46]
      end else begin
        packet_valid_1 <= _GEN_11526;
      end
    end
    packet_rob_idx_1 <= _GEN_11786[6:0];
    if (reset) begin // @[TestHarness.scala 196:31]
      packet_valid_2 <= 1'h0; // @[TestHarness.scala 196:31]
    end else if (_T_212) begin // @[TestHarness.scala 199:26]
      if (io_from_noc_2_flit_bits_tail) begin // @[TestHarness.scala 216:31]
        packet_valid_2 <= 1'h0; // @[TestHarness.scala 216:46]
      end else begin
        packet_valid_2 <= _GEN_13323;
      end
    end
    packet_rob_idx_2 <= _GEN_13583[6:0];
    if (reset) begin // @[TestHarness.scala 196:31]
      packet_valid_3 <= 1'h0; // @[TestHarness.scala 196:31]
    end else if (_T_259) begin // @[TestHarness.scala 199:26]
      if (io_from_noc_3_flit_bits_tail) begin // @[TestHarness.scala 216:31]
        packet_valid_3 <= 1'h0; // @[TestHarness.scala 216:46]
      end else begin
        packet_valid_3 <= _GEN_15120;
      end
    end
    packet_rob_idx_3 <= _GEN_15380[6:0];
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~idle_counter[10])) begin
          $fwrite(32'h80000002,"Assertion failed\n    at TestHarness.scala:148 assert(!idle_counter(10))\n"); // @[TestHarness.scala 148:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (success & _T_3) begin
          $fwrite(32'h80000002,"%d flits, %d cycles\n",flits,tsc); // @[TestHarness.scala 166:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_118 & _T_3 & ~_T_76[0]) begin
          $fwrite(32'h80000002,
            "Assertion failed: out[0] unexpected response\n    at TestHarness.scala:201 assert(rob_valids(rob_idx), cf\"out[${i.toString}] unexpected response\")\n"
            ); // @[TestHarness.scala 201:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_15519 & ~(_T_82 == io_from_noc_0_flit_bits_payload)) begin
          $fwrite(32'h80000002,
            "Assertion failed: out[0] incorrect payload\n    at TestHarness.scala:202 assert(rob_payload(rob_idx).asUInt === o.flit.bits.payload.asUInt, cf\"out[${i.toString}] incorrect payload\");\n"
            ); // @[TestHarness.scala 202:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_15519 & ~(io_from_noc_0_flit_bits_ingress_id == _GEN_8704)) begin
          $fwrite(32'h80000002,
            "Assertion failed: out[0] incorrect source\n    at TestHarness.scala:203 assert(o.flit.bits.ingress_id === rob_ingress_id(rob_idx), cf\"out[${i.toString}] incorrect source\")\n"
            ); // @[TestHarness.scala 203:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_15519 & ~(2'h0 == _GEN_8832)) begin
          $fwrite(32'h80000002,
            "Assertion failed: out[0] incorrect destination\n    at TestHarness.scala:204 assert(i.U === rob_egress_id(rob_idx), cf\"out[${i.toString}] incorrect destination\")\n"
            ); // @[TestHarness.scala 204:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_15519 & ~(_GEN_8960 < _GEN_9088)) begin
          $fwrite(32'h80000002,
            "Assertion failed: out[0] too many flits returned\n    at TestHarness.scala:205 assert(rob_flits_returned(rob_idx) < rob_n_flits(rob_idx), cf\"out[${i.toString}] too many flits returned\")\n"
            ); // @[TestHarness.scala 205:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_15519 & ~(~packet_valid & io_from_noc_0_flit_bits_head | out_payload_rob_idx == _GEN_15381)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at TestHarness.scala:206 assert((!packet_valid && o.flit.bits.head) || rob_idx === packet_rob_idx)\n"
            ); // @[TestHarness.scala 206:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_118 & _T_110 & _T_3) begin
          $fwrite(32'h80000002,"%d, 0, %d\n",_GEN_8704,tsc - out_payload_tsc); // @[TestHarness.scala 210:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_165 & _T_3 & ~_T_123[0]) begin
          $fwrite(32'h80000002,
            "Assertion failed: out[1] unexpected response\n    at TestHarness.scala:201 assert(rob_valids(rob_idx), cf\"out[${i.toString}] unexpected response\")\n"
            ); // @[TestHarness.scala 201:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_15526 & ~(_T_129 == io_from_noc_1_flit_bits_payload)) begin
          $fwrite(32'h80000002,
            "Assertion failed: out[1] incorrect payload\n    at TestHarness.scala:202 assert(rob_payload(rob_idx).asUInt === o.flit.bits.payload.asUInt, cf\"out[${i.toString}] incorrect payload\");\n"
            ); // @[TestHarness.scala 202:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_15526 & ~(io_from_noc_1_flit_bits_ingress_id == _GEN_10501)) begin
          $fwrite(32'h80000002,
            "Assertion failed: out[1] incorrect source\n    at TestHarness.scala:203 assert(o.flit.bits.ingress_id === rob_ingress_id(rob_idx), cf\"out[${i.toString}] incorrect source\")\n"
            ); // @[TestHarness.scala 203:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_15526 & ~(2'h1 == _GEN_10629)) begin
          $fwrite(32'h80000002,
            "Assertion failed: out[1] incorrect destination\n    at TestHarness.scala:204 assert(i.U === rob_egress_id(rob_idx), cf\"out[${i.toString}] incorrect destination\")\n"
            ); // @[TestHarness.scala 204:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_15526 & ~(_GEN_10757 < _GEN_10885)) begin
          $fwrite(32'h80000002,
            "Assertion failed: out[1] too many flits returned\n    at TestHarness.scala:205 assert(rob_flits_returned(rob_idx) < rob_n_flits(rob_idx), cf\"out[${i.toString}] too many flits returned\")\n"
            ); // @[TestHarness.scala 205:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_15526 & ~(~packet_valid_1 & io_from_noc_1_flit_bits_head | out_payload_1_rob_idx == _GEN_15382)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at TestHarness.scala:206 assert((!packet_valid && o.flit.bits.head) || rob_idx === packet_rob_idx)\n"
            ); // @[TestHarness.scala 206:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_165 & _T_157 & _T_3) begin
          $fwrite(32'h80000002,"%d, 1, %d\n",_GEN_10501,tsc - out_payload_1_tsc); // @[TestHarness.scala 210:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_212 & _T_3 & ~_T_170[0]) begin
          $fwrite(32'h80000002,
            "Assertion failed: out[2] unexpected response\n    at TestHarness.scala:201 assert(rob_valids(rob_idx), cf\"out[${i.toString}] unexpected response\")\n"
            ); // @[TestHarness.scala 201:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_15533 & ~(_T_176 == io_from_noc_2_flit_bits_payload)) begin
          $fwrite(32'h80000002,
            "Assertion failed: out[2] incorrect payload\n    at TestHarness.scala:202 assert(rob_payload(rob_idx).asUInt === o.flit.bits.payload.asUInt, cf\"out[${i.toString}] incorrect payload\");\n"
            ); // @[TestHarness.scala 202:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_15533 & ~(io_from_noc_2_flit_bits_ingress_id == _GEN_12298)) begin
          $fwrite(32'h80000002,
            "Assertion failed: out[2] incorrect source\n    at TestHarness.scala:203 assert(o.flit.bits.ingress_id === rob_ingress_id(rob_idx), cf\"out[${i.toString}] incorrect source\")\n"
            ); // @[TestHarness.scala 203:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_15533 & ~(2'h2 == _GEN_12426)) begin
          $fwrite(32'h80000002,
            "Assertion failed: out[2] incorrect destination\n    at TestHarness.scala:204 assert(i.U === rob_egress_id(rob_idx), cf\"out[${i.toString}] incorrect destination\")\n"
            ); // @[TestHarness.scala 204:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_15533 & ~(_GEN_12554 < _GEN_12682)) begin
          $fwrite(32'h80000002,
            "Assertion failed: out[2] too many flits returned\n    at TestHarness.scala:205 assert(rob_flits_returned(rob_idx) < rob_n_flits(rob_idx), cf\"out[${i.toString}] too many flits returned\")\n"
            ); // @[TestHarness.scala 205:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_15533 & ~(~packet_valid_2 & io_from_noc_2_flit_bits_head | out_payload_2_rob_idx == _GEN_15383)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at TestHarness.scala:206 assert((!packet_valid && o.flit.bits.head) || rob_idx === packet_rob_idx)\n"
            ); // @[TestHarness.scala 206:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_212 & _T_204 & _T_3) begin
          $fwrite(32'h80000002,"%d, 2, %d\n",_GEN_12298,tsc - out_payload_2_tsc); // @[TestHarness.scala 210:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_259 & _T_3 & ~_T_217[0]) begin
          $fwrite(32'h80000002,
            "Assertion failed: out[3] unexpected response\n    at TestHarness.scala:201 assert(rob_valids(rob_idx), cf\"out[${i.toString}] unexpected response\")\n"
            ); // @[TestHarness.scala 201:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_15540 & ~(_T_223 == io_from_noc_3_flit_bits_payload)) begin
          $fwrite(32'h80000002,
            "Assertion failed: out[3] incorrect payload\n    at TestHarness.scala:202 assert(rob_payload(rob_idx).asUInt === o.flit.bits.payload.asUInt, cf\"out[${i.toString}] incorrect payload\");\n"
            ); // @[TestHarness.scala 202:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_15540 & ~(io_from_noc_3_flit_bits_ingress_id == _GEN_14095)) begin
          $fwrite(32'h80000002,
            "Assertion failed: out[3] incorrect source\n    at TestHarness.scala:203 assert(o.flit.bits.ingress_id === rob_ingress_id(rob_idx), cf\"out[${i.toString}] incorrect source\")\n"
            ); // @[TestHarness.scala 203:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_15540 & ~(2'h3 == _GEN_14223)) begin
          $fwrite(32'h80000002,
            "Assertion failed: out[3] incorrect destination\n    at TestHarness.scala:204 assert(i.U === rob_egress_id(rob_idx), cf\"out[${i.toString}] incorrect destination\")\n"
            ); // @[TestHarness.scala 204:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_15540 & ~(_GEN_14351 < _GEN_14479)) begin
          $fwrite(32'h80000002,
            "Assertion failed: out[3] too many flits returned\n    at TestHarness.scala:205 assert(rob_flits_returned(rob_idx) < rob_n_flits(rob_idx), cf\"out[${i.toString}] too many flits returned\")\n"
            ); // @[TestHarness.scala 205:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_15540 & ~(~packet_valid_3 & io_from_noc_3_flit_bits_head | out_payload_3_rob_idx == _GEN_15384)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at TestHarness.scala:206 assert((!packet_valid && o.flit.bits.head) || rob_idx === packet_rob_idx)\n"
            ); // @[TestHarness.scala 206:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_259 & _T_251 & _T_3) begin
          $fwrite(32'h80000002,"%d, 3, %d\n",_GEN_14095,tsc - out_payload_3_tsc); // @[TestHarness.scala 210:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[0] & _T_3 & ~(_T_264 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 0 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[1] & _T_3 & ~(_T_271 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 1 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[2] & _T_3 & ~(_T_278 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 2 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[3] & _T_3 & ~(_T_285 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 3 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[4] & _T_3 & ~(_T_292 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 4 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[5] & _T_3 & ~(_T_299 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 5 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[6] & _T_3 & ~(_T_306 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 6 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[7] & _T_3 & ~(_T_313 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 7 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[8] & _T_3 & ~(_T_320 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 8 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[9] & _T_3 & ~(_T_327 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 9 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[10] & _T_3 & ~(_T_334 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 10 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[11] & _T_3 & ~(_T_341 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 11 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[12] & _T_3 & ~(_T_348 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 12 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[13] & _T_3 & ~(_T_355 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 13 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[14] & _T_3 & ~(_T_362 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 14 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[15] & _T_3 & ~(_T_369 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 15 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[16] & _T_3 & ~(_T_376 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 16 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[17] & _T_3 & ~(_T_383 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 17 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[18] & _T_3 & ~(_T_390 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 18 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[19] & _T_3 & ~(_T_397 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 19 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[20] & _T_3 & ~(_T_404 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 20 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[21] & _T_3 & ~(_T_411 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 21 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[22] & _T_3 & ~(_T_418 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 22 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[23] & _T_3 & ~(_T_425 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 23 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[24] & _T_3 & ~(_T_432 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 24 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[25] & _T_3 & ~(_T_439 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 25 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[26] & _T_3 & ~(_T_446 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 26 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[27] & _T_3 & ~(_T_453 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 27 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[28] & _T_3 & ~(_T_460 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 28 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[29] & _T_3 & ~(_T_467 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 29 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[30] & _T_3 & ~(_T_474 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 30 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[31] & _T_3 & ~(_T_481 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 31 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[32] & _T_3 & ~(_T_488 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 32 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[33] & _T_3 & ~(_T_495 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 33 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[34] & _T_3 & ~(_T_502 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 34 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[35] & _T_3 & ~(_T_509 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 35 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[36] & _T_3 & ~(_T_516 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 36 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[37] & _T_3 & ~(_T_523 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 37 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[38] & _T_3 & ~(_T_530 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 38 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[39] & _T_3 & ~(_T_537 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 39 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[40] & _T_3 & ~(_T_544 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 40 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[41] & _T_3 & ~(_T_551 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 41 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[42] & _T_3 & ~(_T_558 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 42 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[43] & _T_3 & ~(_T_565 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 43 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[44] & _T_3 & ~(_T_572 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 44 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[45] & _T_3 & ~(_T_579 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 45 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[46] & _T_3 & ~(_T_586 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 46 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[47] & _T_3 & ~(_T_593 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 47 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[48] & _T_3 & ~(_T_600 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 48 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[49] & _T_3 & ~(_T_607 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 49 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[50] & _T_3 & ~(_T_614 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 50 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[51] & _T_3 & ~(_T_621 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 51 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[52] & _T_3 & ~(_T_628 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 52 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[53] & _T_3 & ~(_T_635 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 53 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[54] & _T_3 & ~(_T_642 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 54 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[55] & _T_3 & ~(_T_649 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 55 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[56] & _T_3 & ~(_T_656 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 56 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[57] & _T_3 & ~(_T_663 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 57 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[58] & _T_3 & ~(_T_670 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 58 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[59] & _T_3 & ~(_T_677 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 59 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[60] & _T_3 & ~(_T_684 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 60 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[61] & _T_3 & ~(_T_691 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 61 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[62] & _T_3 & ~(_T_698 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 62 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[63] & _T_3 & ~(_T_705 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 63 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[64] & _T_3 & ~(_T_712 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 64 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[65] & _T_3 & ~(_T_719 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 65 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[66] & _T_3 & ~(_T_726 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 66 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[67] & _T_3 & ~(_T_733 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 67 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[68] & _T_3 & ~(_T_740 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 68 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[69] & _T_3 & ~(_T_747 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 69 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[70] & _T_3 & ~(_T_754 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 70 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[71] & _T_3 & ~(_T_761 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 71 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[72] & _T_3 & ~(_T_768 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 72 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[73] & _T_3 & ~(_T_775 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 73 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[74] & _T_3 & ~(_T_782 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 74 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[75] & _T_3 & ~(_T_789 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 75 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[76] & _T_3 & ~(_T_796 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 76 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[77] & _T_3 & ~(_T_803 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 77 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[78] & _T_3 & ~(_T_810 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 78 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[79] & _T_3 & ~(_T_817 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 79 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[80] & _T_3 & ~(_T_824 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 80 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[81] & _T_3 & ~(_T_831 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 81 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[82] & _T_3 & ~(_T_838 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 82 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[83] & _T_3 & ~(_T_845 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 83 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[84] & _T_3 & ~(_T_852 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 84 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[85] & _T_3 & ~(_T_859 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 85 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[86] & _T_3 & ~(_T_866 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 86 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[87] & _T_3 & ~(_T_873 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 87 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[88] & _T_3 & ~(_T_880 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 88 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[89] & _T_3 & ~(_T_887 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 89 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[90] & _T_3 & ~(_T_894 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 90 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[91] & _T_3 & ~(_T_901 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 91 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[92] & _T_3 & ~(_T_908 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 92 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[93] & _T_3 & ~(_T_915 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 93 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[94] & _T_3 & ~(_T_922 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 94 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[95] & _T_3 & ~(_T_929 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 95 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[96] & _T_3 & ~(_T_936 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 96 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[97] & _T_3 & ~(_T_943 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 97 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[98] & _T_3 & ~(_T_950 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 98 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[99] & _T_3 & ~(_T_957 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 99 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[100] & _T_3 & ~(_T_964 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 100 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[101] & _T_3 & ~(_T_971 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 101 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[102] & _T_3 & ~(_T_978 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 102 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[103] & _T_3 & ~(_T_985 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 103 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[104] & _T_3 & ~(_T_992 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 104 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[105] & _T_3 & ~(_T_999 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 105 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[106] & _T_3 & ~(_T_1006 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 106 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[107] & _T_3 & ~(_T_1013 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 107 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[108] & _T_3 & ~(_T_1020 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 108 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[109] & _T_3 & ~(_T_1027 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 109 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[110] & _T_3 & ~(_T_1034 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 110 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[111] & _T_3 & ~(_T_1041 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 111 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[112] & _T_3 & ~(_T_1048 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 112 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[113] & _T_3 & ~(_T_1055 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 113 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[114] & _T_3 & ~(_T_1062 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 114 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[115] & _T_3 & ~(_T_1069 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 115 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[116] & _T_3 & ~(_T_1076 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 116 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[117] & _T_3 & ~(_T_1083 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 117 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[118] & _T_3 & ~(_T_1090 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 118 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[119] & _T_3 & ~(_T_1097 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 119 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[120] & _T_3 & ~(_T_1104 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 120 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[121] & _T_3 & ~(_T_1111 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 121 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[122] & _T_3 & ~(_T_1118 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 122 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[123] & _T_3 & ~(_T_1125 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 123 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[124] & _T_3 & ~(_T_1132 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 124 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[125] & _T_3 & ~(_T_1139 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 125 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[126] & _T_3 & ~(_T_1146 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 126 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[127] & _T_3 & ~(_T_1153 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 127 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  txs = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  flits = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  tsc = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  idle_counter = _RAND_3[10:0];
  _RAND_4 = {4{`RANDOM}};
  rob_valids = _RAND_4[127:0];
  _RAND_5 = {1{`RANDOM}};
  rob_payload_0_tsc = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  rob_payload_0_rob_idx = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  rob_payload_0_flits_fired = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  rob_payload_1_tsc = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  rob_payload_1_rob_idx = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  rob_payload_1_flits_fired = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  rob_payload_2_tsc = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  rob_payload_2_rob_idx = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  rob_payload_2_flits_fired = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  rob_payload_3_tsc = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  rob_payload_3_rob_idx = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  rob_payload_3_flits_fired = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  rob_payload_4_tsc = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  rob_payload_4_rob_idx = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  rob_payload_4_flits_fired = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  rob_payload_5_tsc = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  rob_payload_5_rob_idx = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  rob_payload_5_flits_fired = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  rob_payload_6_tsc = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  rob_payload_6_rob_idx = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  rob_payload_6_flits_fired = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  rob_payload_7_tsc = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  rob_payload_7_rob_idx = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  rob_payload_7_flits_fired = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  rob_payload_8_tsc = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  rob_payload_8_rob_idx = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  rob_payload_8_flits_fired = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  rob_payload_9_tsc = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  rob_payload_9_rob_idx = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  rob_payload_9_flits_fired = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  rob_payload_10_tsc = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  rob_payload_10_rob_idx = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  rob_payload_10_flits_fired = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  rob_payload_11_tsc = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  rob_payload_11_rob_idx = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  rob_payload_11_flits_fired = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  rob_payload_12_tsc = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  rob_payload_12_rob_idx = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  rob_payload_12_flits_fired = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  rob_payload_13_tsc = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  rob_payload_13_rob_idx = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  rob_payload_13_flits_fired = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  rob_payload_14_tsc = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  rob_payload_14_rob_idx = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  rob_payload_14_flits_fired = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  rob_payload_15_tsc = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  rob_payload_15_rob_idx = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  rob_payload_15_flits_fired = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  rob_payload_16_tsc = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  rob_payload_16_rob_idx = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  rob_payload_16_flits_fired = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  rob_payload_17_tsc = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  rob_payload_17_rob_idx = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  rob_payload_17_flits_fired = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  rob_payload_18_tsc = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  rob_payload_18_rob_idx = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  rob_payload_18_flits_fired = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  rob_payload_19_tsc = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  rob_payload_19_rob_idx = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  rob_payload_19_flits_fired = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  rob_payload_20_tsc = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  rob_payload_20_rob_idx = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  rob_payload_20_flits_fired = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  rob_payload_21_tsc = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  rob_payload_21_rob_idx = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  rob_payload_21_flits_fired = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  rob_payload_22_tsc = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  rob_payload_22_rob_idx = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  rob_payload_22_flits_fired = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  rob_payload_23_tsc = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  rob_payload_23_rob_idx = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  rob_payload_23_flits_fired = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  rob_payload_24_tsc = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  rob_payload_24_rob_idx = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  rob_payload_24_flits_fired = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  rob_payload_25_tsc = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  rob_payload_25_rob_idx = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  rob_payload_25_flits_fired = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  rob_payload_26_tsc = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  rob_payload_26_rob_idx = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  rob_payload_26_flits_fired = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  rob_payload_27_tsc = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  rob_payload_27_rob_idx = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  rob_payload_27_flits_fired = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  rob_payload_28_tsc = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  rob_payload_28_rob_idx = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  rob_payload_28_flits_fired = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  rob_payload_29_tsc = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  rob_payload_29_rob_idx = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  rob_payload_29_flits_fired = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  rob_payload_30_tsc = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  rob_payload_30_rob_idx = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  rob_payload_30_flits_fired = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  rob_payload_31_tsc = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  rob_payload_31_rob_idx = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  rob_payload_31_flits_fired = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  rob_payload_32_tsc = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  rob_payload_32_rob_idx = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  rob_payload_32_flits_fired = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  rob_payload_33_tsc = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  rob_payload_33_rob_idx = _RAND_105[15:0];
  _RAND_106 = {1{`RANDOM}};
  rob_payload_33_flits_fired = _RAND_106[15:0];
  _RAND_107 = {1{`RANDOM}};
  rob_payload_34_tsc = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  rob_payload_34_rob_idx = _RAND_108[15:0];
  _RAND_109 = {1{`RANDOM}};
  rob_payload_34_flits_fired = _RAND_109[15:0];
  _RAND_110 = {1{`RANDOM}};
  rob_payload_35_tsc = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  rob_payload_35_rob_idx = _RAND_111[15:0];
  _RAND_112 = {1{`RANDOM}};
  rob_payload_35_flits_fired = _RAND_112[15:0];
  _RAND_113 = {1{`RANDOM}};
  rob_payload_36_tsc = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  rob_payload_36_rob_idx = _RAND_114[15:0];
  _RAND_115 = {1{`RANDOM}};
  rob_payload_36_flits_fired = _RAND_115[15:0];
  _RAND_116 = {1{`RANDOM}};
  rob_payload_37_tsc = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  rob_payload_37_rob_idx = _RAND_117[15:0];
  _RAND_118 = {1{`RANDOM}};
  rob_payload_37_flits_fired = _RAND_118[15:0];
  _RAND_119 = {1{`RANDOM}};
  rob_payload_38_tsc = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  rob_payload_38_rob_idx = _RAND_120[15:0];
  _RAND_121 = {1{`RANDOM}};
  rob_payload_38_flits_fired = _RAND_121[15:0];
  _RAND_122 = {1{`RANDOM}};
  rob_payload_39_tsc = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  rob_payload_39_rob_idx = _RAND_123[15:0];
  _RAND_124 = {1{`RANDOM}};
  rob_payload_39_flits_fired = _RAND_124[15:0];
  _RAND_125 = {1{`RANDOM}};
  rob_payload_40_tsc = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  rob_payload_40_rob_idx = _RAND_126[15:0];
  _RAND_127 = {1{`RANDOM}};
  rob_payload_40_flits_fired = _RAND_127[15:0];
  _RAND_128 = {1{`RANDOM}};
  rob_payload_41_tsc = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  rob_payload_41_rob_idx = _RAND_129[15:0];
  _RAND_130 = {1{`RANDOM}};
  rob_payload_41_flits_fired = _RAND_130[15:0];
  _RAND_131 = {1{`RANDOM}};
  rob_payload_42_tsc = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  rob_payload_42_rob_idx = _RAND_132[15:0];
  _RAND_133 = {1{`RANDOM}};
  rob_payload_42_flits_fired = _RAND_133[15:0];
  _RAND_134 = {1{`RANDOM}};
  rob_payload_43_tsc = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  rob_payload_43_rob_idx = _RAND_135[15:0];
  _RAND_136 = {1{`RANDOM}};
  rob_payload_43_flits_fired = _RAND_136[15:0];
  _RAND_137 = {1{`RANDOM}};
  rob_payload_44_tsc = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  rob_payload_44_rob_idx = _RAND_138[15:0];
  _RAND_139 = {1{`RANDOM}};
  rob_payload_44_flits_fired = _RAND_139[15:0];
  _RAND_140 = {1{`RANDOM}};
  rob_payload_45_tsc = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  rob_payload_45_rob_idx = _RAND_141[15:0];
  _RAND_142 = {1{`RANDOM}};
  rob_payload_45_flits_fired = _RAND_142[15:0];
  _RAND_143 = {1{`RANDOM}};
  rob_payload_46_tsc = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  rob_payload_46_rob_idx = _RAND_144[15:0];
  _RAND_145 = {1{`RANDOM}};
  rob_payload_46_flits_fired = _RAND_145[15:0];
  _RAND_146 = {1{`RANDOM}};
  rob_payload_47_tsc = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  rob_payload_47_rob_idx = _RAND_147[15:0];
  _RAND_148 = {1{`RANDOM}};
  rob_payload_47_flits_fired = _RAND_148[15:0];
  _RAND_149 = {1{`RANDOM}};
  rob_payload_48_tsc = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  rob_payload_48_rob_idx = _RAND_150[15:0];
  _RAND_151 = {1{`RANDOM}};
  rob_payload_48_flits_fired = _RAND_151[15:0];
  _RAND_152 = {1{`RANDOM}};
  rob_payload_49_tsc = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  rob_payload_49_rob_idx = _RAND_153[15:0];
  _RAND_154 = {1{`RANDOM}};
  rob_payload_49_flits_fired = _RAND_154[15:0];
  _RAND_155 = {1{`RANDOM}};
  rob_payload_50_tsc = _RAND_155[31:0];
  _RAND_156 = {1{`RANDOM}};
  rob_payload_50_rob_idx = _RAND_156[15:0];
  _RAND_157 = {1{`RANDOM}};
  rob_payload_50_flits_fired = _RAND_157[15:0];
  _RAND_158 = {1{`RANDOM}};
  rob_payload_51_tsc = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  rob_payload_51_rob_idx = _RAND_159[15:0];
  _RAND_160 = {1{`RANDOM}};
  rob_payload_51_flits_fired = _RAND_160[15:0];
  _RAND_161 = {1{`RANDOM}};
  rob_payload_52_tsc = _RAND_161[31:0];
  _RAND_162 = {1{`RANDOM}};
  rob_payload_52_rob_idx = _RAND_162[15:0];
  _RAND_163 = {1{`RANDOM}};
  rob_payload_52_flits_fired = _RAND_163[15:0];
  _RAND_164 = {1{`RANDOM}};
  rob_payload_53_tsc = _RAND_164[31:0];
  _RAND_165 = {1{`RANDOM}};
  rob_payload_53_rob_idx = _RAND_165[15:0];
  _RAND_166 = {1{`RANDOM}};
  rob_payload_53_flits_fired = _RAND_166[15:0];
  _RAND_167 = {1{`RANDOM}};
  rob_payload_54_tsc = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  rob_payload_54_rob_idx = _RAND_168[15:0];
  _RAND_169 = {1{`RANDOM}};
  rob_payload_54_flits_fired = _RAND_169[15:0];
  _RAND_170 = {1{`RANDOM}};
  rob_payload_55_tsc = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  rob_payload_55_rob_idx = _RAND_171[15:0];
  _RAND_172 = {1{`RANDOM}};
  rob_payload_55_flits_fired = _RAND_172[15:0];
  _RAND_173 = {1{`RANDOM}};
  rob_payload_56_tsc = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  rob_payload_56_rob_idx = _RAND_174[15:0];
  _RAND_175 = {1{`RANDOM}};
  rob_payload_56_flits_fired = _RAND_175[15:0];
  _RAND_176 = {1{`RANDOM}};
  rob_payload_57_tsc = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  rob_payload_57_rob_idx = _RAND_177[15:0];
  _RAND_178 = {1{`RANDOM}};
  rob_payload_57_flits_fired = _RAND_178[15:0];
  _RAND_179 = {1{`RANDOM}};
  rob_payload_58_tsc = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  rob_payload_58_rob_idx = _RAND_180[15:0];
  _RAND_181 = {1{`RANDOM}};
  rob_payload_58_flits_fired = _RAND_181[15:0];
  _RAND_182 = {1{`RANDOM}};
  rob_payload_59_tsc = _RAND_182[31:0];
  _RAND_183 = {1{`RANDOM}};
  rob_payload_59_rob_idx = _RAND_183[15:0];
  _RAND_184 = {1{`RANDOM}};
  rob_payload_59_flits_fired = _RAND_184[15:0];
  _RAND_185 = {1{`RANDOM}};
  rob_payload_60_tsc = _RAND_185[31:0];
  _RAND_186 = {1{`RANDOM}};
  rob_payload_60_rob_idx = _RAND_186[15:0];
  _RAND_187 = {1{`RANDOM}};
  rob_payload_60_flits_fired = _RAND_187[15:0];
  _RAND_188 = {1{`RANDOM}};
  rob_payload_61_tsc = _RAND_188[31:0];
  _RAND_189 = {1{`RANDOM}};
  rob_payload_61_rob_idx = _RAND_189[15:0];
  _RAND_190 = {1{`RANDOM}};
  rob_payload_61_flits_fired = _RAND_190[15:0];
  _RAND_191 = {1{`RANDOM}};
  rob_payload_62_tsc = _RAND_191[31:0];
  _RAND_192 = {1{`RANDOM}};
  rob_payload_62_rob_idx = _RAND_192[15:0];
  _RAND_193 = {1{`RANDOM}};
  rob_payload_62_flits_fired = _RAND_193[15:0];
  _RAND_194 = {1{`RANDOM}};
  rob_payload_63_tsc = _RAND_194[31:0];
  _RAND_195 = {1{`RANDOM}};
  rob_payload_63_rob_idx = _RAND_195[15:0];
  _RAND_196 = {1{`RANDOM}};
  rob_payload_63_flits_fired = _RAND_196[15:0];
  _RAND_197 = {1{`RANDOM}};
  rob_payload_64_tsc = _RAND_197[31:0];
  _RAND_198 = {1{`RANDOM}};
  rob_payload_64_rob_idx = _RAND_198[15:0];
  _RAND_199 = {1{`RANDOM}};
  rob_payload_64_flits_fired = _RAND_199[15:0];
  _RAND_200 = {1{`RANDOM}};
  rob_payload_65_tsc = _RAND_200[31:0];
  _RAND_201 = {1{`RANDOM}};
  rob_payload_65_rob_idx = _RAND_201[15:0];
  _RAND_202 = {1{`RANDOM}};
  rob_payload_65_flits_fired = _RAND_202[15:0];
  _RAND_203 = {1{`RANDOM}};
  rob_payload_66_tsc = _RAND_203[31:0];
  _RAND_204 = {1{`RANDOM}};
  rob_payload_66_rob_idx = _RAND_204[15:0];
  _RAND_205 = {1{`RANDOM}};
  rob_payload_66_flits_fired = _RAND_205[15:0];
  _RAND_206 = {1{`RANDOM}};
  rob_payload_67_tsc = _RAND_206[31:0];
  _RAND_207 = {1{`RANDOM}};
  rob_payload_67_rob_idx = _RAND_207[15:0];
  _RAND_208 = {1{`RANDOM}};
  rob_payload_67_flits_fired = _RAND_208[15:0];
  _RAND_209 = {1{`RANDOM}};
  rob_payload_68_tsc = _RAND_209[31:0];
  _RAND_210 = {1{`RANDOM}};
  rob_payload_68_rob_idx = _RAND_210[15:0];
  _RAND_211 = {1{`RANDOM}};
  rob_payload_68_flits_fired = _RAND_211[15:0];
  _RAND_212 = {1{`RANDOM}};
  rob_payload_69_tsc = _RAND_212[31:0];
  _RAND_213 = {1{`RANDOM}};
  rob_payload_69_rob_idx = _RAND_213[15:0];
  _RAND_214 = {1{`RANDOM}};
  rob_payload_69_flits_fired = _RAND_214[15:0];
  _RAND_215 = {1{`RANDOM}};
  rob_payload_70_tsc = _RAND_215[31:0];
  _RAND_216 = {1{`RANDOM}};
  rob_payload_70_rob_idx = _RAND_216[15:0];
  _RAND_217 = {1{`RANDOM}};
  rob_payload_70_flits_fired = _RAND_217[15:0];
  _RAND_218 = {1{`RANDOM}};
  rob_payload_71_tsc = _RAND_218[31:0];
  _RAND_219 = {1{`RANDOM}};
  rob_payload_71_rob_idx = _RAND_219[15:0];
  _RAND_220 = {1{`RANDOM}};
  rob_payload_71_flits_fired = _RAND_220[15:0];
  _RAND_221 = {1{`RANDOM}};
  rob_payload_72_tsc = _RAND_221[31:0];
  _RAND_222 = {1{`RANDOM}};
  rob_payload_72_rob_idx = _RAND_222[15:0];
  _RAND_223 = {1{`RANDOM}};
  rob_payload_72_flits_fired = _RAND_223[15:0];
  _RAND_224 = {1{`RANDOM}};
  rob_payload_73_tsc = _RAND_224[31:0];
  _RAND_225 = {1{`RANDOM}};
  rob_payload_73_rob_idx = _RAND_225[15:0];
  _RAND_226 = {1{`RANDOM}};
  rob_payload_73_flits_fired = _RAND_226[15:0];
  _RAND_227 = {1{`RANDOM}};
  rob_payload_74_tsc = _RAND_227[31:0];
  _RAND_228 = {1{`RANDOM}};
  rob_payload_74_rob_idx = _RAND_228[15:0];
  _RAND_229 = {1{`RANDOM}};
  rob_payload_74_flits_fired = _RAND_229[15:0];
  _RAND_230 = {1{`RANDOM}};
  rob_payload_75_tsc = _RAND_230[31:0];
  _RAND_231 = {1{`RANDOM}};
  rob_payload_75_rob_idx = _RAND_231[15:0];
  _RAND_232 = {1{`RANDOM}};
  rob_payload_75_flits_fired = _RAND_232[15:0];
  _RAND_233 = {1{`RANDOM}};
  rob_payload_76_tsc = _RAND_233[31:0];
  _RAND_234 = {1{`RANDOM}};
  rob_payload_76_rob_idx = _RAND_234[15:0];
  _RAND_235 = {1{`RANDOM}};
  rob_payload_76_flits_fired = _RAND_235[15:0];
  _RAND_236 = {1{`RANDOM}};
  rob_payload_77_tsc = _RAND_236[31:0];
  _RAND_237 = {1{`RANDOM}};
  rob_payload_77_rob_idx = _RAND_237[15:0];
  _RAND_238 = {1{`RANDOM}};
  rob_payload_77_flits_fired = _RAND_238[15:0];
  _RAND_239 = {1{`RANDOM}};
  rob_payload_78_tsc = _RAND_239[31:0];
  _RAND_240 = {1{`RANDOM}};
  rob_payload_78_rob_idx = _RAND_240[15:0];
  _RAND_241 = {1{`RANDOM}};
  rob_payload_78_flits_fired = _RAND_241[15:0];
  _RAND_242 = {1{`RANDOM}};
  rob_payload_79_tsc = _RAND_242[31:0];
  _RAND_243 = {1{`RANDOM}};
  rob_payload_79_rob_idx = _RAND_243[15:0];
  _RAND_244 = {1{`RANDOM}};
  rob_payload_79_flits_fired = _RAND_244[15:0];
  _RAND_245 = {1{`RANDOM}};
  rob_payload_80_tsc = _RAND_245[31:0];
  _RAND_246 = {1{`RANDOM}};
  rob_payload_80_rob_idx = _RAND_246[15:0];
  _RAND_247 = {1{`RANDOM}};
  rob_payload_80_flits_fired = _RAND_247[15:0];
  _RAND_248 = {1{`RANDOM}};
  rob_payload_81_tsc = _RAND_248[31:0];
  _RAND_249 = {1{`RANDOM}};
  rob_payload_81_rob_idx = _RAND_249[15:0];
  _RAND_250 = {1{`RANDOM}};
  rob_payload_81_flits_fired = _RAND_250[15:0];
  _RAND_251 = {1{`RANDOM}};
  rob_payload_82_tsc = _RAND_251[31:0];
  _RAND_252 = {1{`RANDOM}};
  rob_payload_82_rob_idx = _RAND_252[15:0];
  _RAND_253 = {1{`RANDOM}};
  rob_payload_82_flits_fired = _RAND_253[15:0];
  _RAND_254 = {1{`RANDOM}};
  rob_payload_83_tsc = _RAND_254[31:0];
  _RAND_255 = {1{`RANDOM}};
  rob_payload_83_rob_idx = _RAND_255[15:0];
  _RAND_256 = {1{`RANDOM}};
  rob_payload_83_flits_fired = _RAND_256[15:0];
  _RAND_257 = {1{`RANDOM}};
  rob_payload_84_tsc = _RAND_257[31:0];
  _RAND_258 = {1{`RANDOM}};
  rob_payload_84_rob_idx = _RAND_258[15:0];
  _RAND_259 = {1{`RANDOM}};
  rob_payload_84_flits_fired = _RAND_259[15:0];
  _RAND_260 = {1{`RANDOM}};
  rob_payload_85_tsc = _RAND_260[31:0];
  _RAND_261 = {1{`RANDOM}};
  rob_payload_85_rob_idx = _RAND_261[15:0];
  _RAND_262 = {1{`RANDOM}};
  rob_payload_85_flits_fired = _RAND_262[15:0];
  _RAND_263 = {1{`RANDOM}};
  rob_payload_86_tsc = _RAND_263[31:0];
  _RAND_264 = {1{`RANDOM}};
  rob_payload_86_rob_idx = _RAND_264[15:0];
  _RAND_265 = {1{`RANDOM}};
  rob_payload_86_flits_fired = _RAND_265[15:0];
  _RAND_266 = {1{`RANDOM}};
  rob_payload_87_tsc = _RAND_266[31:0];
  _RAND_267 = {1{`RANDOM}};
  rob_payload_87_rob_idx = _RAND_267[15:0];
  _RAND_268 = {1{`RANDOM}};
  rob_payload_87_flits_fired = _RAND_268[15:0];
  _RAND_269 = {1{`RANDOM}};
  rob_payload_88_tsc = _RAND_269[31:0];
  _RAND_270 = {1{`RANDOM}};
  rob_payload_88_rob_idx = _RAND_270[15:0];
  _RAND_271 = {1{`RANDOM}};
  rob_payload_88_flits_fired = _RAND_271[15:0];
  _RAND_272 = {1{`RANDOM}};
  rob_payload_89_tsc = _RAND_272[31:0];
  _RAND_273 = {1{`RANDOM}};
  rob_payload_89_rob_idx = _RAND_273[15:0];
  _RAND_274 = {1{`RANDOM}};
  rob_payload_89_flits_fired = _RAND_274[15:0];
  _RAND_275 = {1{`RANDOM}};
  rob_payload_90_tsc = _RAND_275[31:0];
  _RAND_276 = {1{`RANDOM}};
  rob_payload_90_rob_idx = _RAND_276[15:0];
  _RAND_277 = {1{`RANDOM}};
  rob_payload_90_flits_fired = _RAND_277[15:0];
  _RAND_278 = {1{`RANDOM}};
  rob_payload_91_tsc = _RAND_278[31:0];
  _RAND_279 = {1{`RANDOM}};
  rob_payload_91_rob_idx = _RAND_279[15:0];
  _RAND_280 = {1{`RANDOM}};
  rob_payload_91_flits_fired = _RAND_280[15:0];
  _RAND_281 = {1{`RANDOM}};
  rob_payload_92_tsc = _RAND_281[31:0];
  _RAND_282 = {1{`RANDOM}};
  rob_payload_92_rob_idx = _RAND_282[15:0];
  _RAND_283 = {1{`RANDOM}};
  rob_payload_92_flits_fired = _RAND_283[15:0];
  _RAND_284 = {1{`RANDOM}};
  rob_payload_93_tsc = _RAND_284[31:0];
  _RAND_285 = {1{`RANDOM}};
  rob_payload_93_rob_idx = _RAND_285[15:0];
  _RAND_286 = {1{`RANDOM}};
  rob_payload_93_flits_fired = _RAND_286[15:0];
  _RAND_287 = {1{`RANDOM}};
  rob_payload_94_tsc = _RAND_287[31:0];
  _RAND_288 = {1{`RANDOM}};
  rob_payload_94_rob_idx = _RAND_288[15:0];
  _RAND_289 = {1{`RANDOM}};
  rob_payload_94_flits_fired = _RAND_289[15:0];
  _RAND_290 = {1{`RANDOM}};
  rob_payload_95_tsc = _RAND_290[31:0];
  _RAND_291 = {1{`RANDOM}};
  rob_payload_95_rob_idx = _RAND_291[15:0];
  _RAND_292 = {1{`RANDOM}};
  rob_payload_95_flits_fired = _RAND_292[15:0];
  _RAND_293 = {1{`RANDOM}};
  rob_payload_96_tsc = _RAND_293[31:0];
  _RAND_294 = {1{`RANDOM}};
  rob_payload_96_rob_idx = _RAND_294[15:0];
  _RAND_295 = {1{`RANDOM}};
  rob_payload_96_flits_fired = _RAND_295[15:0];
  _RAND_296 = {1{`RANDOM}};
  rob_payload_97_tsc = _RAND_296[31:0];
  _RAND_297 = {1{`RANDOM}};
  rob_payload_97_rob_idx = _RAND_297[15:0];
  _RAND_298 = {1{`RANDOM}};
  rob_payload_97_flits_fired = _RAND_298[15:0];
  _RAND_299 = {1{`RANDOM}};
  rob_payload_98_tsc = _RAND_299[31:0];
  _RAND_300 = {1{`RANDOM}};
  rob_payload_98_rob_idx = _RAND_300[15:0];
  _RAND_301 = {1{`RANDOM}};
  rob_payload_98_flits_fired = _RAND_301[15:0];
  _RAND_302 = {1{`RANDOM}};
  rob_payload_99_tsc = _RAND_302[31:0];
  _RAND_303 = {1{`RANDOM}};
  rob_payload_99_rob_idx = _RAND_303[15:0];
  _RAND_304 = {1{`RANDOM}};
  rob_payload_99_flits_fired = _RAND_304[15:0];
  _RAND_305 = {1{`RANDOM}};
  rob_payload_100_tsc = _RAND_305[31:0];
  _RAND_306 = {1{`RANDOM}};
  rob_payload_100_rob_idx = _RAND_306[15:0];
  _RAND_307 = {1{`RANDOM}};
  rob_payload_100_flits_fired = _RAND_307[15:0];
  _RAND_308 = {1{`RANDOM}};
  rob_payload_101_tsc = _RAND_308[31:0];
  _RAND_309 = {1{`RANDOM}};
  rob_payload_101_rob_idx = _RAND_309[15:0];
  _RAND_310 = {1{`RANDOM}};
  rob_payload_101_flits_fired = _RAND_310[15:0];
  _RAND_311 = {1{`RANDOM}};
  rob_payload_102_tsc = _RAND_311[31:0];
  _RAND_312 = {1{`RANDOM}};
  rob_payload_102_rob_idx = _RAND_312[15:0];
  _RAND_313 = {1{`RANDOM}};
  rob_payload_102_flits_fired = _RAND_313[15:0];
  _RAND_314 = {1{`RANDOM}};
  rob_payload_103_tsc = _RAND_314[31:0];
  _RAND_315 = {1{`RANDOM}};
  rob_payload_103_rob_idx = _RAND_315[15:0];
  _RAND_316 = {1{`RANDOM}};
  rob_payload_103_flits_fired = _RAND_316[15:0];
  _RAND_317 = {1{`RANDOM}};
  rob_payload_104_tsc = _RAND_317[31:0];
  _RAND_318 = {1{`RANDOM}};
  rob_payload_104_rob_idx = _RAND_318[15:0];
  _RAND_319 = {1{`RANDOM}};
  rob_payload_104_flits_fired = _RAND_319[15:0];
  _RAND_320 = {1{`RANDOM}};
  rob_payload_105_tsc = _RAND_320[31:0];
  _RAND_321 = {1{`RANDOM}};
  rob_payload_105_rob_idx = _RAND_321[15:0];
  _RAND_322 = {1{`RANDOM}};
  rob_payload_105_flits_fired = _RAND_322[15:0];
  _RAND_323 = {1{`RANDOM}};
  rob_payload_106_tsc = _RAND_323[31:0];
  _RAND_324 = {1{`RANDOM}};
  rob_payload_106_rob_idx = _RAND_324[15:0];
  _RAND_325 = {1{`RANDOM}};
  rob_payload_106_flits_fired = _RAND_325[15:0];
  _RAND_326 = {1{`RANDOM}};
  rob_payload_107_tsc = _RAND_326[31:0];
  _RAND_327 = {1{`RANDOM}};
  rob_payload_107_rob_idx = _RAND_327[15:0];
  _RAND_328 = {1{`RANDOM}};
  rob_payload_107_flits_fired = _RAND_328[15:0];
  _RAND_329 = {1{`RANDOM}};
  rob_payload_108_tsc = _RAND_329[31:0];
  _RAND_330 = {1{`RANDOM}};
  rob_payload_108_rob_idx = _RAND_330[15:0];
  _RAND_331 = {1{`RANDOM}};
  rob_payload_108_flits_fired = _RAND_331[15:0];
  _RAND_332 = {1{`RANDOM}};
  rob_payload_109_tsc = _RAND_332[31:0];
  _RAND_333 = {1{`RANDOM}};
  rob_payload_109_rob_idx = _RAND_333[15:0];
  _RAND_334 = {1{`RANDOM}};
  rob_payload_109_flits_fired = _RAND_334[15:0];
  _RAND_335 = {1{`RANDOM}};
  rob_payload_110_tsc = _RAND_335[31:0];
  _RAND_336 = {1{`RANDOM}};
  rob_payload_110_rob_idx = _RAND_336[15:0];
  _RAND_337 = {1{`RANDOM}};
  rob_payload_110_flits_fired = _RAND_337[15:0];
  _RAND_338 = {1{`RANDOM}};
  rob_payload_111_tsc = _RAND_338[31:0];
  _RAND_339 = {1{`RANDOM}};
  rob_payload_111_rob_idx = _RAND_339[15:0];
  _RAND_340 = {1{`RANDOM}};
  rob_payload_111_flits_fired = _RAND_340[15:0];
  _RAND_341 = {1{`RANDOM}};
  rob_payload_112_tsc = _RAND_341[31:0];
  _RAND_342 = {1{`RANDOM}};
  rob_payload_112_rob_idx = _RAND_342[15:0];
  _RAND_343 = {1{`RANDOM}};
  rob_payload_112_flits_fired = _RAND_343[15:0];
  _RAND_344 = {1{`RANDOM}};
  rob_payload_113_tsc = _RAND_344[31:0];
  _RAND_345 = {1{`RANDOM}};
  rob_payload_113_rob_idx = _RAND_345[15:0];
  _RAND_346 = {1{`RANDOM}};
  rob_payload_113_flits_fired = _RAND_346[15:0];
  _RAND_347 = {1{`RANDOM}};
  rob_payload_114_tsc = _RAND_347[31:0];
  _RAND_348 = {1{`RANDOM}};
  rob_payload_114_rob_idx = _RAND_348[15:0];
  _RAND_349 = {1{`RANDOM}};
  rob_payload_114_flits_fired = _RAND_349[15:0];
  _RAND_350 = {1{`RANDOM}};
  rob_payload_115_tsc = _RAND_350[31:0];
  _RAND_351 = {1{`RANDOM}};
  rob_payload_115_rob_idx = _RAND_351[15:0];
  _RAND_352 = {1{`RANDOM}};
  rob_payload_115_flits_fired = _RAND_352[15:0];
  _RAND_353 = {1{`RANDOM}};
  rob_payload_116_tsc = _RAND_353[31:0];
  _RAND_354 = {1{`RANDOM}};
  rob_payload_116_rob_idx = _RAND_354[15:0];
  _RAND_355 = {1{`RANDOM}};
  rob_payload_116_flits_fired = _RAND_355[15:0];
  _RAND_356 = {1{`RANDOM}};
  rob_payload_117_tsc = _RAND_356[31:0];
  _RAND_357 = {1{`RANDOM}};
  rob_payload_117_rob_idx = _RAND_357[15:0];
  _RAND_358 = {1{`RANDOM}};
  rob_payload_117_flits_fired = _RAND_358[15:0];
  _RAND_359 = {1{`RANDOM}};
  rob_payload_118_tsc = _RAND_359[31:0];
  _RAND_360 = {1{`RANDOM}};
  rob_payload_118_rob_idx = _RAND_360[15:0];
  _RAND_361 = {1{`RANDOM}};
  rob_payload_118_flits_fired = _RAND_361[15:0];
  _RAND_362 = {1{`RANDOM}};
  rob_payload_119_tsc = _RAND_362[31:0];
  _RAND_363 = {1{`RANDOM}};
  rob_payload_119_rob_idx = _RAND_363[15:0];
  _RAND_364 = {1{`RANDOM}};
  rob_payload_119_flits_fired = _RAND_364[15:0];
  _RAND_365 = {1{`RANDOM}};
  rob_payload_120_tsc = _RAND_365[31:0];
  _RAND_366 = {1{`RANDOM}};
  rob_payload_120_rob_idx = _RAND_366[15:0];
  _RAND_367 = {1{`RANDOM}};
  rob_payload_120_flits_fired = _RAND_367[15:0];
  _RAND_368 = {1{`RANDOM}};
  rob_payload_121_tsc = _RAND_368[31:0];
  _RAND_369 = {1{`RANDOM}};
  rob_payload_121_rob_idx = _RAND_369[15:0];
  _RAND_370 = {1{`RANDOM}};
  rob_payload_121_flits_fired = _RAND_370[15:0];
  _RAND_371 = {1{`RANDOM}};
  rob_payload_122_tsc = _RAND_371[31:0];
  _RAND_372 = {1{`RANDOM}};
  rob_payload_122_rob_idx = _RAND_372[15:0];
  _RAND_373 = {1{`RANDOM}};
  rob_payload_122_flits_fired = _RAND_373[15:0];
  _RAND_374 = {1{`RANDOM}};
  rob_payload_123_tsc = _RAND_374[31:0];
  _RAND_375 = {1{`RANDOM}};
  rob_payload_123_rob_idx = _RAND_375[15:0];
  _RAND_376 = {1{`RANDOM}};
  rob_payload_123_flits_fired = _RAND_376[15:0];
  _RAND_377 = {1{`RANDOM}};
  rob_payload_124_tsc = _RAND_377[31:0];
  _RAND_378 = {1{`RANDOM}};
  rob_payload_124_rob_idx = _RAND_378[15:0];
  _RAND_379 = {1{`RANDOM}};
  rob_payload_124_flits_fired = _RAND_379[15:0];
  _RAND_380 = {1{`RANDOM}};
  rob_payload_125_tsc = _RAND_380[31:0];
  _RAND_381 = {1{`RANDOM}};
  rob_payload_125_rob_idx = _RAND_381[15:0];
  _RAND_382 = {1{`RANDOM}};
  rob_payload_125_flits_fired = _RAND_382[15:0];
  _RAND_383 = {1{`RANDOM}};
  rob_payload_126_tsc = _RAND_383[31:0];
  _RAND_384 = {1{`RANDOM}};
  rob_payload_126_rob_idx = _RAND_384[15:0];
  _RAND_385 = {1{`RANDOM}};
  rob_payload_126_flits_fired = _RAND_385[15:0];
  _RAND_386 = {1{`RANDOM}};
  rob_payload_127_tsc = _RAND_386[31:0];
  _RAND_387 = {1{`RANDOM}};
  rob_payload_127_rob_idx = _RAND_387[15:0];
  _RAND_388 = {1{`RANDOM}};
  rob_payload_127_flits_fired = _RAND_388[15:0];
  _RAND_389 = {1{`RANDOM}};
  rob_egress_id_0 = _RAND_389[1:0];
  _RAND_390 = {1{`RANDOM}};
  rob_egress_id_1 = _RAND_390[1:0];
  _RAND_391 = {1{`RANDOM}};
  rob_egress_id_2 = _RAND_391[1:0];
  _RAND_392 = {1{`RANDOM}};
  rob_egress_id_3 = _RAND_392[1:0];
  _RAND_393 = {1{`RANDOM}};
  rob_egress_id_4 = _RAND_393[1:0];
  _RAND_394 = {1{`RANDOM}};
  rob_egress_id_5 = _RAND_394[1:0];
  _RAND_395 = {1{`RANDOM}};
  rob_egress_id_6 = _RAND_395[1:0];
  _RAND_396 = {1{`RANDOM}};
  rob_egress_id_7 = _RAND_396[1:0];
  _RAND_397 = {1{`RANDOM}};
  rob_egress_id_8 = _RAND_397[1:0];
  _RAND_398 = {1{`RANDOM}};
  rob_egress_id_9 = _RAND_398[1:0];
  _RAND_399 = {1{`RANDOM}};
  rob_egress_id_10 = _RAND_399[1:0];
  _RAND_400 = {1{`RANDOM}};
  rob_egress_id_11 = _RAND_400[1:0];
  _RAND_401 = {1{`RANDOM}};
  rob_egress_id_12 = _RAND_401[1:0];
  _RAND_402 = {1{`RANDOM}};
  rob_egress_id_13 = _RAND_402[1:0];
  _RAND_403 = {1{`RANDOM}};
  rob_egress_id_14 = _RAND_403[1:0];
  _RAND_404 = {1{`RANDOM}};
  rob_egress_id_15 = _RAND_404[1:0];
  _RAND_405 = {1{`RANDOM}};
  rob_egress_id_16 = _RAND_405[1:0];
  _RAND_406 = {1{`RANDOM}};
  rob_egress_id_17 = _RAND_406[1:0];
  _RAND_407 = {1{`RANDOM}};
  rob_egress_id_18 = _RAND_407[1:0];
  _RAND_408 = {1{`RANDOM}};
  rob_egress_id_19 = _RAND_408[1:0];
  _RAND_409 = {1{`RANDOM}};
  rob_egress_id_20 = _RAND_409[1:0];
  _RAND_410 = {1{`RANDOM}};
  rob_egress_id_21 = _RAND_410[1:0];
  _RAND_411 = {1{`RANDOM}};
  rob_egress_id_22 = _RAND_411[1:0];
  _RAND_412 = {1{`RANDOM}};
  rob_egress_id_23 = _RAND_412[1:0];
  _RAND_413 = {1{`RANDOM}};
  rob_egress_id_24 = _RAND_413[1:0];
  _RAND_414 = {1{`RANDOM}};
  rob_egress_id_25 = _RAND_414[1:0];
  _RAND_415 = {1{`RANDOM}};
  rob_egress_id_26 = _RAND_415[1:0];
  _RAND_416 = {1{`RANDOM}};
  rob_egress_id_27 = _RAND_416[1:0];
  _RAND_417 = {1{`RANDOM}};
  rob_egress_id_28 = _RAND_417[1:0];
  _RAND_418 = {1{`RANDOM}};
  rob_egress_id_29 = _RAND_418[1:0];
  _RAND_419 = {1{`RANDOM}};
  rob_egress_id_30 = _RAND_419[1:0];
  _RAND_420 = {1{`RANDOM}};
  rob_egress_id_31 = _RAND_420[1:0];
  _RAND_421 = {1{`RANDOM}};
  rob_egress_id_32 = _RAND_421[1:0];
  _RAND_422 = {1{`RANDOM}};
  rob_egress_id_33 = _RAND_422[1:0];
  _RAND_423 = {1{`RANDOM}};
  rob_egress_id_34 = _RAND_423[1:0];
  _RAND_424 = {1{`RANDOM}};
  rob_egress_id_35 = _RAND_424[1:0];
  _RAND_425 = {1{`RANDOM}};
  rob_egress_id_36 = _RAND_425[1:0];
  _RAND_426 = {1{`RANDOM}};
  rob_egress_id_37 = _RAND_426[1:0];
  _RAND_427 = {1{`RANDOM}};
  rob_egress_id_38 = _RAND_427[1:0];
  _RAND_428 = {1{`RANDOM}};
  rob_egress_id_39 = _RAND_428[1:0];
  _RAND_429 = {1{`RANDOM}};
  rob_egress_id_40 = _RAND_429[1:0];
  _RAND_430 = {1{`RANDOM}};
  rob_egress_id_41 = _RAND_430[1:0];
  _RAND_431 = {1{`RANDOM}};
  rob_egress_id_42 = _RAND_431[1:0];
  _RAND_432 = {1{`RANDOM}};
  rob_egress_id_43 = _RAND_432[1:0];
  _RAND_433 = {1{`RANDOM}};
  rob_egress_id_44 = _RAND_433[1:0];
  _RAND_434 = {1{`RANDOM}};
  rob_egress_id_45 = _RAND_434[1:0];
  _RAND_435 = {1{`RANDOM}};
  rob_egress_id_46 = _RAND_435[1:0];
  _RAND_436 = {1{`RANDOM}};
  rob_egress_id_47 = _RAND_436[1:0];
  _RAND_437 = {1{`RANDOM}};
  rob_egress_id_48 = _RAND_437[1:0];
  _RAND_438 = {1{`RANDOM}};
  rob_egress_id_49 = _RAND_438[1:0];
  _RAND_439 = {1{`RANDOM}};
  rob_egress_id_50 = _RAND_439[1:0];
  _RAND_440 = {1{`RANDOM}};
  rob_egress_id_51 = _RAND_440[1:0];
  _RAND_441 = {1{`RANDOM}};
  rob_egress_id_52 = _RAND_441[1:0];
  _RAND_442 = {1{`RANDOM}};
  rob_egress_id_53 = _RAND_442[1:0];
  _RAND_443 = {1{`RANDOM}};
  rob_egress_id_54 = _RAND_443[1:0];
  _RAND_444 = {1{`RANDOM}};
  rob_egress_id_55 = _RAND_444[1:0];
  _RAND_445 = {1{`RANDOM}};
  rob_egress_id_56 = _RAND_445[1:0];
  _RAND_446 = {1{`RANDOM}};
  rob_egress_id_57 = _RAND_446[1:0];
  _RAND_447 = {1{`RANDOM}};
  rob_egress_id_58 = _RAND_447[1:0];
  _RAND_448 = {1{`RANDOM}};
  rob_egress_id_59 = _RAND_448[1:0];
  _RAND_449 = {1{`RANDOM}};
  rob_egress_id_60 = _RAND_449[1:0];
  _RAND_450 = {1{`RANDOM}};
  rob_egress_id_61 = _RAND_450[1:0];
  _RAND_451 = {1{`RANDOM}};
  rob_egress_id_62 = _RAND_451[1:0];
  _RAND_452 = {1{`RANDOM}};
  rob_egress_id_63 = _RAND_452[1:0];
  _RAND_453 = {1{`RANDOM}};
  rob_egress_id_64 = _RAND_453[1:0];
  _RAND_454 = {1{`RANDOM}};
  rob_egress_id_65 = _RAND_454[1:0];
  _RAND_455 = {1{`RANDOM}};
  rob_egress_id_66 = _RAND_455[1:0];
  _RAND_456 = {1{`RANDOM}};
  rob_egress_id_67 = _RAND_456[1:0];
  _RAND_457 = {1{`RANDOM}};
  rob_egress_id_68 = _RAND_457[1:0];
  _RAND_458 = {1{`RANDOM}};
  rob_egress_id_69 = _RAND_458[1:0];
  _RAND_459 = {1{`RANDOM}};
  rob_egress_id_70 = _RAND_459[1:0];
  _RAND_460 = {1{`RANDOM}};
  rob_egress_id_71 = _RAND_460[1:0];
  _RAND_461 = {1{`RANDOM}};
  rob_egress_id_72 = _RAND_461[1:0];
  _RAND_462 = {1{`RANDOM}};
  rob_egress_id_73 = _RAND_462[1:0];
  _RAND_463 = {1{`RANDOM}};
  rob_egress_id_74 = _RAND_463[1:0];
  _RAND_464 = {1{`RANDOM}};
  rob_egress_id_75 = _RAND_464[1:0];
  _RAND_465 = {1{`RANDOM}};
  rob_egress_id_76 = _RAND_465[1:0];
  _RAND_466 = {1{`RANDOM}};
  rob_egress_id_77 = _RAND_466[1:0];
  _RAND_467 = {1{`RANDOM}};
  rob_egress_id_78 = _RAND_467[1:0];
  _RAND_468 = {1{`RANDOM}};
  rob_egress_id_79 = _RAND_468[1:0];
  _RAND_469 = {1{`RANDOM}};
  rob_egress_id_80 = _RAND_469[1:0];
  _RAND_470 = {1{`RANDOM}};
  rob_egress_id_81 = _RAND_470[1:0];
  _RAND_471 = {1{`RANDOM}};
  rob_egress_id_82 = _RAND_471[1:0];
  _RAND_472 = {1{`RANDOM}};
  rob_egress_id_83 = _RAND_472[1:0];
  _RAND_473 = {1{`RANDOM}};
  rob_egress_id_84 = _RAND_473[1:0];
  _RAND_474 = {1{`RANDOM}};
  rob_egress_id_85 = _RAND_474[1:0];
  _RAND_475 = {1{`RANDOM}};
  rob_egress_id_86 = _RAND_475[1:0];
  _RAND_476 = {1{`RANDOM}};
  rob_egress_id_87 = _RAND_476[1:0];
  _RAND_477 = {1{`RANDOM}};
  rob_egress_id_88 = _RAND_477[1:0];
  _RAND_478 = {1{`RANDOM}};
  rob_egress_id_89 = _RAND_478[1:0];
  _RAND_479 = {1{`RANDOM}};
  rob_egress_id_90 = _RAND_479[1:0];
  _RAND_480 = {1{`RANDOM}};
  rob_egress_id_91 = _RAND_480[1:0];
  _RAND_481 = {1{`RANDOM}};
  rob_egress_id_92 = _RAND_481[1:0];
  _RAND_482 = {1{`RANDOM}};
  rob_egress_id_93 = _RAND_482[1:0];
  _RAND_483 = {1{`RANDOM}};
  rob_egress_id_94 = _RAND_483[1:0];
  _RAND_484 = {1{`RANDOM}};
  rob_egress_id_95 = _RAND_484[1:0];
  _RAND_485 = {1{`RANDOM}};
  rob_egress_id_96 = _RAND_485[1:0];
  _RAND_486 = {1{`RANDOM}};
  rob_egress_id_97 = _RAND_486[1:0];
  _RAND_487 = {1{`RANDOM}};
  rob_egress_id_98 = _RAND_487[1:0];
  _RAND_488 = {1{`RANDOM}};
  rob_egress_id_99 = _RAND_488[1:0];
  _RAND_489 = {1{`RANDOM}};
  rob_egress_id_100 = _RAND_489[1:0];
  _RAND_490 = {1{`RANDOM}};
  rob_egress_id_101 = _RAND_490[1:0];
  _RAND_491 = {1{`RANDOM}};
  rob_egress_id_102 = _RAND_491[1:0];
  _RAND_492 = {1{`RANDOM}};
  rob_egress_id_103 = _RAND_492[1:0];
  _RAND_493 = {1{`RANDOM}};
  rob_egress_id_104 = _RAND_493[1:0];
  _RAND_494 = {1{`RANDOM}};
  rob_egress_id_105 = _RAND_494[1:0];
  _RAND_495 = {1{`RANDOM}};
  rob_egress_id_106 = _RAND_495[1:0];
  _RAND_496 = {1{`RANDOM}};
  rob_egress_id_107 = _RAND_496[1:0];
  _RAND_497 = {1{`RANDOM}};
  rob_egress_id_108 = _RAND_497[1:0];
  _RAND_498 = {1{`RANDOM}};
  rob_egress_id_109 = _RAND_498[1:0];
  _RAND_499 = {1{`RANDOM}};
  rob_egress_id_110 = _RAND_499[1:0];
  _RAND_500 = {1{`RANDOM}};
  rob_egress_id_111 = _RAND_500[1:0];
  _RAND_501 = {1{`RANDOM}};
  rob_egress_id_112 = _RAND_501[1:0];
  _RAND_502 = {1{`RANDOM}};
  rob_egress_id_113 = _RAND_502[1:0];
  _RAND_503 = {1{`RANDOM}};
  rob_egress_id_114 = _RAND_503[1:0];
  _RAND_504 = {1{`RANDOM}};
  rob_egress_id_115 = _RAND_504[1:0];
  _RAND_505 = {1{`RANDOM}};
  rob_egress_id_116 = _RAND_505[1:0];
  _RAND_506 = {1{`RANDOM}};
  rob_egress_id_117 = _RAND_506[1:0];
  _RAND_507 = {1{`RANDOM}};
  rob_egress_id_118 = _RAND_507[1:0];
  _RAND_508 = {1{`RANDOM}};
  rob_egress_id_119 = _RAND_508[1:0];
  _RAND_509 = {1{`RANDOM}};
  rob_egress_id_120 = _RAND_509[1:0];
  _RAND_510 = {1{`RANDOM}};
  rob_egress_id_121 = _RAND_510[1:0];
  _RAND_511 = {1{`RANDOM}};
  rob_egress_id_122 = _RAND_511[1:0];
  _RAND_512 = {1{`RANDOM}};
  rob_egress_id_123 = _RAND_512[1:0];
  _RAND_513 = {1{`RANDOM}};
  rob_egress_id_124 = _RAND_513[1:0];
  _RAND_514 = {1{`RANDOM}};
  rob_egress_id_125 = _RAND_514[1:0];
  _RAND_515 = {1{`RANDOM}};
  rob_egress_id_126 = _RAND_515[1:0];
  _RAND_516 = {1{`RANDOM}};
  rob_egress_id_127 = _RAND_516[1:0];
  _RAND_517 = {1{`RANDOM}};
  rob_ingress_id_0 = _RAND_517[1:0];
  _RAND_518 = {1{`RANDOM}};
  rob_ingress_id_1 = _RAND_518[1:0];
  _RAND_519 = {1{`RANDOM}};
  rob_ingress_id_2 = _RAND_519[1:0];
  _RAND_520 = {1{`RANDOM}};
  rob_ingress_id_3 = _RAND_520[1:0];
  _RAND_521 = {1{`RANDOM}};
  rob_ingress_id_4 = _RAND_521[1:0];
  _RAND_522 = {1{`RANDOM}};
  rob_ingress_id_5 = _RAND_522[1:0];
  _RAND_523 = {1{`RANDOM}};
  rob_ingress_id_6 = _RAND_523[1:0];
  _RAND_524 = {1{`RANDOM}};
  rob_ingress_id_7 = _RAND_524[1:0];
  _RAND_525 = {1{`RANDOM}};
  rob_ingress_id_8 = _RAND_525[1:0];
  _RAND_526 = {1{`RANDOM}};
  rob_ingress_id_9 = _RAND_526[1:0];
  _RAND_527 = {1{`RANDOM}};
  rob_ingress_id_10 = _RAND_527[1:0];
  _RAND_528 = {1{`RANDOM}};
  rob_ingress_id_11 = _RAND_528[1:0];
  _RAND_529 = {1{`RANDOM}};
  rob_ingress_id_12 = _RAND_529[1:0];
  _RAND_530 = {1{`RANDOM}};
  rob_ingress_id_13 = _RAND_530[1:0];
  _RAND_531 = {1{`RANDOM}};
  rob_ingress_id_14 = _RAND_531[1:0];
  _RAND_532 = {1{`RANDOM}};
  rob_ingress_id_15 = _RAND_532[1:0];
  _RAND_533 = {1{`RANDOM}};
  rob_ingress_id_16 = _RAND_533[1:0];
  _RAND_534 = {1{`RANDOM}};
  rob_ingress_id_17 = _RAND_534[1:0];
  _RAND_535 = {1{`RANDOM}};
  rob_ingress_id_18 = _RAND_535[1:0];
  _RAND_536 = {1{`RANDOM}};
  rob_ingress_id_19 = _RAND_536[1:0];
  _RAND_537 = {1{`RANDOM}};
  rob_ingress_id_20 = _RAND_537[1:0];
  _RAND_538 = {1{`RANDOM}};
  rob_ingress_id_21 = _RAND_538[1:0];
  _RAND_539 = {1{`RANDOM}};
  rob_ingress_id_22 = _RAND_539[1:0];
  _RAND_540 = {1{`RANDOM}};
  rob_ingress_id_23 = _RAND_540[1:0];
  _RAND_541 = {1{`RANDOM}};
  rob_ingress_id_24 = _RAND_541[1:0];
  _RAND_542 = {1{`RANDOM}};
  rob_ingress_id_25 = _RAND_542[1:0];
  _RAND_543 = {1{`RANDOM}};
  rob_ingress_id_26 = _RAND_543[1:0];
  _RAND_544 = {1{`RANDOM}};
  rob_ingress_id_27 = _RAND_544[1:0];
  _RAND_545 = {1{`RANDOM}};
  rob_ingress_id_28 = _RAND_545[1:0];
  _RAND_546 = {1{`RANDOM}};
  rob_ingress_id_29 = _RAND_546[1:0];
  _RAND_547 = {1{`RANDOM}};
  rob_ingress_id_30 = _RAND_547[1:0];
  _RAND_548 = {1{`RANDOM}};
  rob_ingress_id_31 = _RAND_548[1:0];
  _RAND_549 = {1{`RANDOM}};
  rob_ingress_id_32 = _RAND_549[1:0];
  _RAND_550 = {1{`RANDOM}};
  rob_ingress_id_33 = _RAND_550[1:0];
  _RAND_551 = {1{`RANDOM}};
  rob_ingress_id_34 = _RAND_551[1:0];
  _RAND_552 = {1{`RANDOM}};
  rob_ingress_id_35 = _RAND_552[1:0];
  _RAND_553 = {1{`RANDOM}};
  rob_ingress_id_36 = _RAND_553[1:0];
  _RAND_554 = {1{`RANDOM}};
  rob_ingress_id_37 = _RAND_554[1:0];
  _RAND_555 = {1{`RANDOM}};
  rob_ingress_id_38 = _RAND_555[1:0];
  _RAND_556 = {1{`RANDOM}};
  rob_ingress_id_39 = _RAND_556[1:0];
  _RAND_557 = {1{`RANDOM}};
  rob_ingress_id_40 = _RAND_557[1:0];
  _RAND_558 = {1{`RANDOM}};
  rob_ingress_id_41 = _RAND_558[1:0];
  _RAND_559 = {1{`RANDOM}};
  rob_ingress_id_42 = _RAND_559[1:0];
  _RAND_560 = {1{`RANDOM}};
  rob_ingress_id_43 = _RAND_560[1:0];
  _RAND_561 = {1{`RANDOM}};
  rob_ingress_id_44 = _RAND_561[1:0];
  _RAND_562 = {1{`RANDOM}};
  rob_ingress_id_45 = _RAND_562[1:0];
  _RAND_563 = {1{`RANDOM}};
  rob_ingress_id_46 = _RAND_563[1:0];
  _RAND_564 = {1{`RANDOM}};
  rob_ingress_id_47 = _RAND_564[1:0];
  _RAND_565 = {1{`RANDOM}};
  rob_ingress_id_48 = _RAND_565[1:0];
  _RAND_566 = {1{`RANDOM}};
  rob_ingress_id_49 = _RAND_566[1:0];
  _RAND_567 = {1{`RANDOM}};
  rob_ingress_id_50 = _RAND_567[1:0];
  _RAND_568 = {1{`RANDOM}};
  rob_ingress_id_51 = _RAND_568[1:0];
  _RAND_569 = {1{`RANDOM}};
  rob_ingress_id_52 = _RAND_569[1:0];
  _RAND_570 = {1{`RANDOM}};
  rob_ingress_id_53 = _RAND_570[1:0];
  _RAND_571 = {1{`RANDOM}};
  rob_ingress_id_54 = _RAND_571[1:0];
  _RAND_572 = {1{`RANDOM}};
  rob_ingress_id_55 = _RAND_572[1:0];
  _RAND_573 = {1{`RANDOM}};
  rob_ingress_id_56 = _RAND_573[1:0];
  _RAND_574 = {1{`RANDOM}};
  rob_ingress_id_57 = _RAND_574[1:0];
  _RAND_575 = {1{`RANDOM}};
  rob_ingress_id_58 = _RAND_575[1:0];
  _RAND_576 = {1{`RANDOM}};
  rob_ingress_id_59 = _RAND_576[1:0];
  _RAND_577 = {1{`RANDOM}};
  rob_ingress_id_60 = _RAND_577[1:0];
  _RAND_578 = {1{`RANDOM}};
  rob_ingress_id_61 = _RAND_578[1:0];
  _RAND_579 = {1{`RANDOM}};
  rob_ingress_id_62 = _RAND_579[1:0];
  _RAND_580 = {1{`RANDOM}};
  rob_ingress_id_63 = _RAND_580[1:0];
  _RAND_581 = {1{`RANDOM}};
  rob_ingress_id_64 = _RAND_581[1:0];
  _RAND_582 = {1{`RANDOM}};
  rob_ingress_id_65 = _RAND_582[1:0];
  _RAND_583 = {1{`RANDOM}};
  rob_ingress_id_66 = _RAND_583[1:0];
  _RAND_584 = {1{`RANDOM}};
  rob_ingress_id_67 = _RAND_584[1:0];
  _RAND_585 = {1{`RANDOM}};
  rob_ingress_id_68 = _RAND_585[1:0];
  _RAND_586 = {1{`RANDOM}};
  rob_ingress_id_69 = _RAND_586[1:0];
  _RAND_587 = {1{`RANDOM}};
  rob_ingress_id_70 = _RAND_587[1:0];
  _RAND_588 = {1{`RANDOM}};
  rob_ingress_id_71 = _RAND_588[1:0];
  _RAND_589 = {1{`RANDOM}};
  rob_ingress_id_72 = _RAND_589[1:0];
  _RAND_590 = {1{`RANDOM}};
  rob_ingress_id_73 = _RAND_590[1:0];
  _RAND_591 = {1{`RANDOM}};
  rob_ingress_id_74 = _RAND_591[1:0];
  _RAND_592 = {1{`RANDOM}};
  rob_ingress_id_75 = _RAND_592[1:0];
  _RAND_593 = {1{`RANDOM}};
  rob_ingress_id_76 = _RAND_593[1:0];
  _RAND_594 = {1{`RANDOM}};
  rob_ingress_id_77 = _RAND_594[1:0];
  _RAND_595 = {1{`RANDOM}};
  rob_ingress_id_78 = _RAND_595[1:0];
  _RAND_596 = {1{`RANDOM}};
  rob_ingress_id_79 = _RAND_596[1:0];
  _RAND_597 = {1{`RANDOM}};
  rob_ingress_id_80 = _RAND_597[1:0];
  _RAND_598 = {1{`RANDOM}};
  rob_ingress_id_81 = _RAND_598[1:0];
  _RAND_599 = {1{`RANDOM}};
  rob_ingress_id_82 = _RAND_599[1:0];
  _RAND_600 = {1{`RANDOM}};
  rob_ingress_id_83 = _RAND_600[1:0];
  _RAND_601 = {1{`RANDOM}};
  rob_ingress_id_84 = _RAND_601[1:0];
  _RAND_602 = {1{`RANDOM}};
  rob_ingress_id_85 = _RAND_602[1:0];
  _RAND_603 = {1{`RANDOM}};
  rob_ingress_id_86 = _RAND_603[1:0];
  _RAND_604 = {1{`RANDOM}};
  rob_ingress_id_87 = _RAND_604[1:0];
  _RAND_605 = {1{`RANDOM}};
  rob_ingress_id_88 = _RAND_605[1:0];
  _RAND_606 = {1{`RANDOM}};
  rob_ingress_id_89 = _RAND_606[1:0];
  _RAND_607 = {1{`RANDOM}};
  rob_ingress_id_90 = _RAND_607[1:0];
  _RAND_608 = {1{`RANDOM}};
  rob_ingress_id_91 = _RAND_608[1:0];
  _RAND_609 = {1{`RANDOM}};
  rob_ingress_id_92 = _RAND_609[1:0];
  _RAND_610 = {1{`RANDOM}};
  rob_ingress_id_93 = _RAND_610[1:0];
  _RAND_611 = {1{`RANDOM}};
  rob_ingress_id_94 = _RAND_611[1:0];
  _RAND_612 = {1{`RANDOM}};
  rob_ingress_id_95 = _RAND_612[1:0];
  _RAND_613 = {1{`RANDOM}};
  rob_ingress_id_96 = _RAND_613[1:0];
  _RAND_614 = {1{`RANDOM}};
  rob_ingress_id_97 = _RAND_614[1:0];
  _RAND_615 = {1{`RANDOM}};
  rob_ingress_id_98 = _RAND_615[1:0];
  _RAND_616 = {1{`RANDOM}};
  rob_ingress_id_99 = _RAND_616[1:0];
  _RAND_617 = {1{`RANDOM}};
  rob_ingress_id_100 = _RAND_617[1:0];
  _RAND_618 = {1{`RANDOM}};
  rob_ingress_id_101 = _RAND_618[1:0];
  _RAND_619 = {1{`RANDOM}};
  rob_ingress_id_102 = _RAND_619[1:0];
  _RAND_620 = {1{`RANDOM}};
  rob_ingress_id_103 = _RAND_620[1:0];
  _RAND_621 = {1{`RANDOM}};
  rob_ingress_id_104 = _RAND_621[1:0];
  _RAND_622 = {1{`RANDOM}};
  rob_ingress_id_105 = _RAND_622[1:0];
  _RAND_623 = {1{`RANDOM}};
  rob_ingress_id_106 = _RAND_623[1:0];
  _RAND_624 = {1{`RANDOM}};
  rob_ingress_id_107 = _RAND_624[1:0];
  _RAND_625 = {1{`RANDOM}};
  rob_ingress_id_108 = _RAND_625[1:0];
  _RAND_626 = {1{`RANDOM}};
  rob_ingress_id_109 = _RAND_626[1:0];
  _RAND_627 = {1{`RANDOM}};
  rob_ingress_id_110 = _RAND_627[1:0];
  _RAND_628 = {1{`RANDOM}};
  rob_ingress_id_111 = _RAND_628[1:0];
  _RAND_629 = {1{`RANDOM}};
  rob_ingress_id_112 = _RAND_629[1:0];
  _RAND_630 = {1{`RANDOM}};
  rob_ingress_id_113 = _RAND_630[1:0];
  _RAND_631 = {1{`RANDOM}};
  rob_ingress_id_114 = _RAND_631[1:0];
  _RAND_632 = {1{`RANDOM}};
  rob_ingress_id_115 = _RAND_632[1:0];
  _RAND_633 = {1{`RANDOM}};
  rob_ingress_id_116 = _RAND_633[1:0];
  _RAND_634 = {1{`RANDOM}};
  rob_ingress_id_117 = _RAND_634[1:0];
  _RAND_635 = {1{`RANDOM}};
  rob_ingress_id_118 = _RAND_635[1:0];
  _RAND_636 = {1{`RANDOM}};
  rob_ingress_id_119 = _RAND_636[1:0];
  _RAND_637 = {1{`RANDOM}};
  rob_ingress_id_120 = _RAND_637[1:0];
  _RAND_638 = {1{`RANDOM}};
  rob_ingress_id_121 = _RAND_638[1:0];
  _RAND_639 = {1{`RANDOM}};
  rob_ingress_id_122 = _RAND_639[1:0];
  _RAND_640 = {1{`RANDOM}};
  rob_ingress_id_123 = _RAND_640[1:0];
  _RAND_641 = {1{`RANDOM}};
  rob_ingress_id_124 = _RAND_641[1:0];
  _RAND_642 = {1{`RANDOM}};
  rob_ingress_id_125 = _RAND_642[1:0];
  _RAND_643 = {1{`RANDOM}};
  rob_ingress_id_126 = _RAND_643[1:0];
  _RAND_644 = {1{`RANDOM}};
  rob_ingress_id_127 = _RAND_644[1:0];
  _RAND_645 = {1{`RANDOM}};
  rob_n_flits_0 = _RAND_645[3:0];
  _RAND_646 = {1{`RANDOM}};
  rob_n_flits_1 = _RAND_646[3:0];
  _RAND_647 = {1{`RANDOM}};
  rob_n_flits_2 = _RAND_647[3:0];
  _RAND_648 = {1{`RANDOM}};
  rob_n_flits_3 = _RAND_648[3:0];
  _RAND_649 = {1{`RANDOM}};
  rob_n_flits_4 = _RAND_649[3:0];
  _RAND_650 = {1{`RANDOM}};
  rob_n_flits_5 = _RAND_650[3:0];
  _RAND_651 = {1{`RANDOM}};
  rob_n_flits_6 = _RAND_651[3:0];
  _RAND_652 = {1{`RANDOM}};
  rob_n_flits_7 = _RAND_652[3:0];
  _RAND_653 = {1{`RANDOM}};
  rob_n_flits_8 = _RAND_653[3:0];
  _RAND_654 = {1{`RANDOM}};
  rob_n_flits_9 = _RAND_654[3:0];
  _RAND_655 = {1{`RANDOM}};
  rob_n_flits_10 = _RAND_655[3:0];
  _RAND_656 = {1{`RANDOM}};
  rob_n_flits_11 = _RAND_656[3:0];
  _RAND_657 = {1{`RANDOM}};
  rob_n_flits_12 = _RAND_657[3:0];
  _RAND_658 = {1{`RANDOM}};
  rob_n_flits_13 = _RAND_658[3:0];
  _RAND_659 = {1{`RANDOM}};
  rob_n_flits_14 = _RAND_659[3:0];
  _RAND_660 = {1{`RANDOM}};
  rob_n_flits_15 = _RAND_660[3:0];
  _RAND_661 = {1{`RANDOM}};
  rob_n_flits_16 = _RAND_661[3:0];
  _RAND_662 = {1{`RANDOM}};
  rob_n_flits_17 = _RAND_662[3:0];
  _RAND_663 = {1{`RANDOM}};
  rob_n_flits_18 = _RAND_663[3:0];
  _RAND_664 = {1{`RANDOM}};
  rob_n_flits_19 = _RAND_664[3:0];
  _RAND_665 = {1{`RANDOM}};
  rob_n_flits_20 = _RAND_665[3:0];
  _RAND_666 = {1{`RANDOM}};
  rob_n_flits_21 = _RAND_666[3:0];
  _RAND_667 = {1{`RANDOM}};
  rob_n_flits_22 = _RAND_667[3:0];
  _RAND_668 = {1{`RANDOM}};
  rob_n_flits_23 = _RAND_668[3:0];
  _RAND_669 = {1{`RANDOM}};
  rob_n_flits_24 = _RAND_669[3:0];
  _RAND_670 = {1{`RANDOM}};
  rob_n_flits_25 = _RAND_670[3:0];
  _RAND_671 = {1{`RANDOM}};
  rob_n_flits_26 = _RAND_671[3:0];
  _RAND_672 = {1{`RANDOM}};
  rob_n_flits_27 = _RAND_672[3:0];
  _RAND_673 = {1{`RANDOM}};
  rob_n_flits_28 = _RAND_673[3:0];
  _RAND_674 = {1{`RANDOM}};
  rob_n_flits_29 = _RAND_674[3:0];
  _RAND_675 = {1{`RANDOM}};
  rob_n_flits_30 = _RAND_675[3:0];
  _RAND_676 = {1{`RANDOM}};
  rob_n_flits_31 = _RAND_676[3:0];
  _RAND_677 = {1{`RANDOM}};
  rob_n_flits_32 = _RAND_677[3:0];
  _RAND_678 = {1{`RANDOM}};
  rob_n_flits_33 = _RAND_678[3:0];
  _RAND_679 = {1{`RANDOM}};
  rob_n_flits_34 = _RAND_679[3:0];
  _RAND_680 = {1{`RANDOM}};
  rob_n_flits_35 = _RAND_680[3:0];
  _RAND_681 = {1{`RANDOM}};
  rob_n_flits_36 = _RAND_681[3:0];
  _RAND_682 = {1{`RANDOM}};
  rob_n_flits_37 = _RAND_682[3:0];
  _RAND_683 = {1{`RANDOM}};
  rob_n_flits_38 = _RAND_683[3:0];
  _RAND_684 = {1{`RANDOM}};
  rob_n_flits_39 = _RAND_684[3:0];
  _RAND_685 = {1{`RANDOM}};
  rob_n_flits_40 = _RAND_685[3:0];
  _RAND_686 = {1{`RANDOM}};
  rob_n_flits_41 = _RAND_686[3:0];
  _RAND_687 = {1{`RANDOM}};
  rob_n_flits_42 = _RAND_687[3:0];
  _RAND_688 = {1{`RANDOM}};
  rob_n_flits_43 = _RAND_688[3:0];
  _RAND_689 = {1{`RANDOM}};
  rob_n_flits_44 = _RAND_689[3:0];
  _RAND_690 = {1{`RANDOM}};
  rob_n_flits_45 = _RAND_690[3:0];
  _RAND_691 = {1{`RANDOM}};
  rob_n_flits_46 = _RAND_691[3:0];
  _RAND_692 = {1{`RANDOM}};
  rob_n_flits_47 = _RAND_692[3:0];
  _RAND_693 = {1{`RANDOM}};
  rob_n_flits_48 = _RAND_693[3:0];
  _RAND_694 = {1{`RANDOM}};
  rob_n_flits_49 = _RAND_694[3:0];
  _RAND_695 = {1{`RANDOM}};
  rob_n_flits_50 = _RAND_695[3:0];
  _RAND_696 = {1{`RANDOM}};
  rob_n_flits_51 = _RAND_696[3:0];
  _RAND_697 = {1{`RANDOM}};
  rob_n_flits_52 = _RAND_697[3:0];
  _RAND_698 = {1{`RANDOM}};
  rob_n_flits_53 = _RAND_698[3:0];
  _RAND_699 = {1{`RANDOM}};
  rob_n_flits_54 = _RAND_699[3:0];
  _RAND_700 = {1{`RANDOM}};
  rob_n_flits_55 = _RAND_700[3:0];
  _RAND_701 = {1{`RANDOM}};
  rob_n_flits_56 = _RAND_701[3:0];
  _RAND_702 = {1{`RANDOM}};
  rob_n_flits_57 = _RAND_702[3:0];
  _RAND_703 = {1{`RANDOM}};
  rob_n_flits_58 = _RAND_703[3:0];
  _RAND_704 = {1{`RANDOM}};
  rob_n_flits_59 = _RAND_704[3:0];
  _RAND_705 = {1{`RANDOM}};
  rob_n_flits_60 = _RAND_705[3:0];
  _RAND_706 = {1{`RANDOM}};
  rob_n_flits_61 = _RAND_706[3:0];
  _RAND_707 = {1{`RANDOM}};
  rob_n_flits_62 = _RAND_707[3:0];
  _RAND_708 = {1{`RANDOM}};
  rob_n_flits_63 = _RAND_708[3:0];
  _RAND_709 = {1{`RANDOM}};
  rob_n_flits_64 = _RAND_709[3:0];
  _RAND_710 = {1{`RANDOM}};
  rob_n_flits_65 = _RAND_710[3:0];
  _RAND_711 = {1{`RANDOM}};
  rob_n_flits_66 = _RAND_711[3:0];
  _RAND_712 = {1{`RANDOM}};
  rob_n_flits_67 = _RAND_712[3:0];
  _RAND_713 = {1{`RANDOM}};
  rob_n_flits_68 = _RAND_713[3:0];
  _RAND_714 = {1{`RANDOM}};
  rob_n_flits_69 = _RAND_714[3:0];
  _RAND_715 = {1{`RANDOM}};
  rob_n_flits_70 = _RAND_715[3:0];
  _RAND_716 = {1{`RANDOM}};
  rob_n_flits_71 = _RAND_716[3:0];
  _RAND_717 = {1{`RANDOM}};
  rob_n_flits_72 = _RAND_717[3:0];
  _RAND_718 = {1{`RANDOM}};
  rob_n_flits_73 = _RAND_718[3:0];
  _RAND_719 = {1{`RANDOM}};
  rob_n_flits_74 = _RAND_719[3:0];
  _RAND_720 = {1{`RANDOM}};
  rob_n_flits_75 = _RAND_720[3:0];
  _RAND_721 = {1{`RANDOM}};
  rob_n_flits_76 = _RAND_721[3:0];
  _RAND_722 = {1{`RANDOM}};
  rob_n_flits_77 = _RAND_722[3:0];
  _RAND_723 = {1{`RANDOM}};
  rob_n_flits_78 = _RAND_723[3:0];
  _RAND_724 = {1{`RANDOM}};
  rob_n_flits_79 = _RAND_724[3:0];
  _RAND_725 = {1{`RANDOM}};
  rob_n_flits_80 = _RAND_725[3:0];
  _RAND_726 = {1{`RANDOM}};
  rob_n_flits_81 = _RAND_726[3:0];
  _RAND_727 = {1{`RANDOM}};
  rob_n_flits_82 = _RAND_727[3:0];
  _RAND_728 = {1{`RANDOM}};
  rob_n_flits_83 = _RAND_728[3:0];
  _RAND_729 = {1{`RANDOM}};
  rob_n_flits_84 = _RAND_729[3:0];
  _RAND_730 = {1{`RANDOM}};
  rob_n_flits_85 = _RAND_730[3:0];
  _RAND_731 = {1{`RANDOM}};
  rob_n_flits_86 = _RAND_731[3:0];
  _RAND_732 = {1{`RANDOM}};
  rob_n_flits_87 = _RAND_732[3:0];
  _RAND_733 = {1{`RANDOM}};
  rob_n_flits_88 = _RAND_733[3:0];
  _RAND_734 = {1{`RANDOM}};
  rob_n_flits_89 = _RAND_734[3:0];
  _RAND_735 = {1{`RANDOM}};
  rob_n_flits_90 = _RAND_735[3:0];
  _RAND_736 = {1{`RANDOM}};
  rob_n_flits_91 = _RAND_736[3:0];
  _RAND_737 = {1{`RANDOM}};
  rob_n_flits_92 = _RAND_737[3:0];
  _RAND_738 = {1{`RANDOM}};
  rob_n_flits_93 = _RAND_738[3:0];
  _RAND_739 = {1{`RANDOM}};
  rob_n_flits_94 = _RAND_739[3:0];
  _RAND_740 = {1{`RANDOM}};
  rob_n_flits_95 = _RAND_740[3:0];
  _RAND_741 = {1{`RANDOM}};
  rob_n_flits_96 = _RAND_741[3:0];
  _RAND_742 = {1{`RANDOM}};
  rob_n_flits_97 = _RAND_742[3:0];
  _RAND_743 = {1{`RANDOM}};
  rob_n_flits_98 = _RAND_743[3:0];
  _RAND_744 = {1{`RANDOM}};
  rob_n_flits_99 = _RAND_744[3:0];
  _RAND_745 = {1{`RANDOM}};
  rob_n_flits_100 = _RAND_745[3:0];
  _RAND_746 = {1{`RANDOM}};
  rob_n_flits_101 = _RAND_746[3:0];
  _RAND_747 = {1{`RANDOM}};
  rob_n_flits_102 = _RAND_747[3:0];
  _RAND_748 = {1{`RANDOM}};
  rob_n_flits_103 = _RAND_748[3:0];
  _RAND_749 = {1{`RANDOM}};
  rob_n_flits_104 = _RAND_749[3:0];
  _RAND_750 = {1{`RANDOM}};
  rob_n_flits_105 = _RAND_750[3:0];
  _RAND_751 = {1{`RANDOM}};
  rob_n_flits_106 = _RAND_751[3:0];
  _RAND_752 = {1{`RANDOM}};
  rob_n_flits_107 = _RAND_752[3:0];
  _RAND_753 = {1{`RANDOM}};
  rob_n_flits_108 = _RAND_753[3:0];
  _RAND_754 = {1{`RANDOM}};
  rob_n_flits_109 = _RAND_754[3:0];
  _RAND_755 = {1{`RANDOM}};
  rob_n_flits_110 = _RAND_755[3:0];
  _RAND_756 = {1{`RANDOM}};
  rob_n_flits_111 = _RAND_756[3:0];
  _RAND_757 = {1{`RANDOM}};
  rob_n_flits_112 = _RAND_757[3:0];
  _RAND_758 = {1{`RANDOM}};
  rob_n_flits_113 = _RAND_758[3:0];
  _RAND_759 = {1{`RANDOM}};
  rob_n_flits_114 = _RAND_759[3:0];
  _RAND_760 = {1{`RANDOM}};
  rob_n_flits_115 = _RAND_760[3:0];
  _RAND_761 = {1{`RANDOM}};
  rob_n_flits_116 = _RAND_761[3:0];
  _RAND_762 = {1{`RANDOM}};
  rob_n_flits_117 = _RAND_762[3:0];
  _RAND_763 = {1{`RANDOM}};
  rob_n_flits_118 = _RAND_763[3:0];
  _RAND_764 = {1{`RANDOM}};
  rob_n_flits_119 = _RAND_764[3:0];
  _RAND_765 = {1{`RANDOM}};
  rob_n_flits_120 = _RAND_765[3:0];
  _RAND_766 = {1{`RANDOM}};
  rob_n_flits_121 = _RAND_766[3:0];
  _RAND_767 = {1{`RANDOM}};
  rob_n_flits_122 = _RAND_767[3:0];
  _RAND_768 = {1{`RANDOM}};
  rob_n_flits_123 = _RAND_768[3:0];
  _RAND_769 = {1{`RANDOM}};
  rob_n_flits_124 = _RAND_769[3:0];
  _RAND_770 = {1{`RANDOM}};
  rob_n_flits_125 = _RAND_770[3:0];
  _RAND_771 = {1{`RANDOM}};
  rob_n_flits_126 = _RAND_771[3:0];
  _RAND_772 = {1{`RANDOM}};
  rob_n_flits_127 = _RAND_772[3:0];
  _RAND_773 = {1{`RANDOM}};
  rob_flits_returned_0 = _RAND_773[3:0];
  _RAND_774 = {1{`RANDOM}};
  rob_flits_returned_1 = _RAND_774[3:0];
  _RAND_775 = {1{`RANDOM}};
  rob_flits_returned_2 = _RAND_775[3:0];
  _RAND_776 = {1{`RANDOM}};
  rob_flits_returned_3 = _RAND_776[3:0];
  _RAND_777 = {1{`RANDOM}};
  rob_flits_returned_4 = _RAND_777[3:0];
  _RAND_778 = {1{`RANDOM}};
  rob_flits_returned_5 = _RAND_778[3:0];
  _RAND_779 = {1{`RANDOM}};
  rob_flits_returned_6 = _RAND_779[3:0];
  _RAND_780 = {1{`RANDOM}};
  rob_flits_returned_7 = _RAND_780[3:0];
  _RAND_781 = {1{`RANDOM}};
  rob_flits_returned_8 = _RAND_781[3:0];
  _RAND_782 = {1{`RANDOM}};
  rob_flits_returned_9 = _RAND_782[3:0];
  _RAND_783 = {1{`RANDOM}};
  rob_flits_returned_10 = _RAND_783[3:0];
  _RAND_784 = {1{`RANDOM}};
  rob_flits_returned_11 = _RAND_784[3:0];
  _RAND_785 = {1{`RANDOM}};
  rob_flits_returned_12 = _RAND_785[3:0];
  _RAND_786 = {1{`RANDOM}};
  rob_flits_returned_13 = _RAND_786[3:0];
  _RAND_787 = {1{`RANDOM}};
  rob_flits_returned_14 = _RAND_787[3:0];
  _RAND_788 = {1{`RANDOM}};
  rob_flits_returned_15 = _RAND_788[3:0];
  _RAND_789 = {1{`RANDOM}};
  rob_flits_returned_16 = _RAND_789[3:0];
  _RAND_790 = {1{`RANDOM}};
  rob_flits_returned_17 = _RAND_790[3:0];
  _RAND_791 = {1{`RANDOM}};
  rob_flits_returned_18 = _RAND_791[3:0];
  _RAND_792 = {1{`RANDOM}};
  rob_flits_returned_19 = _RAND_792[3:0];
  _RAND_793 = {1{`RANDOM}};
  rob_flits_returned_20 = _RAND_793[3:0];
  _RAND_794 = {1{`RANDOM}};
  rob_flits_returned_21 = _RAND_794[3:0];
  _RAND_795 = {1{`RANDOM}};
  rob_flits_returned_22 = _RAND_795[3:0];
  _RAND_796 = {1{`RANDOM}};
  rob_flits_returned_23 = _RAND_796[3:0];
  _RAND_797 = {1{`RANDOM}};
  rob_flits_returned_24 = _RAND_797[3:0];
  _RAND_798 = {1{`RANDOM}};
  rob_flits_returned_25 = _RAND_798[3:0];
  _RAND_799 = {1{`RANDOM}};
  rob_flits_returned_26 = _RAND_799[3:0];
  _RAND_800 = {1{`RANDOM}};
  rob_flits_returned_27 = _RAND_800[3:0];
  _RAND_801 = {1{`RANDOM}};
  rob_flits_returned_28 = _RAND_801[3:0];
  _RAND_802 = {1{`RANDOM}};
  rob_flits_returned_29 = _RAND_802[3:0];
  _RAND_803 = {1{`RANDOM}};
  rob_flits_returned_30 = _RAND_803[3:0];
  _RAND_804 = {1{`RANDOM}};
  rob_flits_returned_31 = _RAND_804[3:0];
  _RAND_805 = {1{`RANDOM}};
  rob_flits_returned_32 = _RAND_805[3:0];
  _RAND_806 = {1{`RANDOM}};
  rob_flits_returned_33 = _RAND_806[3:0];
  _RAND_807 = {1{`RANDOM}};
  rob_flits_returned_34 = _RAND_807[3:0];
  _RAND_808 = {1{`RANDOM}};
  rob_flits_returned_35 = _RAND_808[3:0];
  _RAND_809 = {1{`RANDOM}};
  rob_flits_returned_36 = _RAND_809[3:0];
  _RAND_810 = {1{`RANDOM}};
  rob_flits_returned_37 = _RAND_810[3:0];
  _RAND_811 = {1{`RANDOM}};
  rob_flits_returned_38 = _RAND_811[3:0];
  _RAND_812 = {1{`RANDOM}};
  rob_flits_returned_39 = _RAND_812[3:0];
  _RAND_813 = {1{`RANDOM}};
  rob_flits_returned_40 = _RAND_813[3:0];
  _RAND_814 = {1{`RANDOM}};
  rob_flits_returned_41 = _RAND_814[3:0];
  _RAND_815 = {1{`RANDOM}};
  rob_flits_returned_42 = _RAND_815[3:0];
  _RAND_816 = {1{`RANDOM}};
  rob_flits_returned_43 = _RAND_816[3:0];
  _RAND_817 = {1{`RANDOM}};
  rob_flits_returned_44 = _RAND_817[3:0];
  _RAND_818 = {1{`RANDOM}};
  rob_flits_returned_45 = _RAND_818[3:0];
  _RAND_819 = {1{`RANDOM}};
  rob_flits_returned_46 = _RAND_819[3:0];
  _RAND_820 = {1{`RANDOM}};
  rob_flits_returned_47 = _RAND_820[3:0];
  _RAND_821 = {1{`RANDOM}};
  rob_flits_returned_48 = _RAND_821[3:0];
  _RAND_822 = {1{`RANDOM}};
  rob_flits_returned_49 = _RAND_822[3:0];
  _RAND_823 = {1{`RANDOM}};
  rob_flits_returned_50 = _RAND_823[3:0];
  _RAND_824 = {1{`RANDOM}};
  rob_flits_returned_51 = _RAND_824[3:0];
  _RAND_825 = {1{`RANDOM}};
  rob_flits_returned_52 = _RAND_825[3:0];
  _RAND_826 = {1{`RANDOM}};
  rob_flits_returned_53 = _RAND_826[3:0];
  _RAND_827 = {1{`RANDOM}};
  rob_flits_returned_54 = _RAND_827[3:0];
  _RAND_828 = {1{`RANDOM}};
  rob_flits_returned_55 = _RAND_828[3:0];
  _RAND_829 = {1{`RANDOM}};
  rob_flits_returned_56 = _RAND_829[3:0];
  _RAND_830 = {1{`RANDOM}};
  rob_flits_returned_57 = _RAND_830[3:0];
  _RAND_831 = {1{`RANDOM}};
  rob_flits_returned_58 = _RAND_831[3:0];
  _RAND_832 = {1{`RANDOM}};
  rob_flits_returned_59 = _RAND_832[3:0];
  _RAND_833 = {1{`RANDOM}};
  rob_flits_returned_60 = _RAND_833[3:0];
  _RAND_834 = {1{`RANDOM}};
  rob_flits_returned_61 = _RAND_834[3:0];
  _RAND_835 = {1{`RANDOM}};
  rob_flits_returned_62 = _RAND_835[3:0];
  _RAND_836 = {1{`RANDOM}};
  rob_flits_returned_63 = _RAND_836[3:0];
  _RAND_837 = {1{`RANDOM}};
  rob_flits_returned_64 = _RAND_837[3:0];
  _RAND_838 = {1{`RANDOM}};
  rob_flits_returned_65 = _RAND_838[3:0];
  _RAND_839 = {1{`RANDOM}};
  rob_flits_returned_66 = _RAND_839[3:0];
  _RAND_840 = {1{`RANDOM}};
  rob_flits_returned_67 = _RAND_840[3:0];
  _RAND_841 = {1{`RANDOM}};
  rob_flits_returned_68 = _RAND_841[3:0];
  _RAND_842 = {1{`RANDOM}};
  rob_flits_returned_69 = _RAND_842[3:0];
  _RAND_843 = {1{`RANDOM}};
  rob_flits_returned_70 = _RAND_843[3:0];
  _RAND_844 = {1{`RANDOM}};
  rob_flits_returned_71 = _RAND_844[3:0];
  _RAND_845 = {1{`RANDOM}};
  rob_flits_returned_72 = _RAND_845[3:0];
  _RAND_846 = {1{`RANDOM}};
  rob_flits_returned_73 = _RAND_846[3:0];
  _RAND_847 = {1{`RANDOM}};
  rob_flits_returned_74 = _RAND_847[3:0];
  _RAND_848 = {1{`RANDOM}};
  rob_flits_returned_75 = _RAND_848[3:0];
  _RAND_849 = {1{`RANDOM}};
  rob_flits_returned_76 = _RAND_849[3:0];
  _RAND_850 = {1{`RANDOM}};
  rob_flits_returned_77 = _RAND_850[3:0];
  _RAND_851 = {1{`RANDOM}};
  rob_flits_returned_78 = _RAND_851[3:0];
  _RAND_852 = {1{`RANDOM}};
  rob_flits_returned_79 = _RAND_852[3:0];
  _RAND_853 = {1{`RANDOM}};
  rob_flits_returned_80 = _RAND_853[3:0];
  _RAND_854 = {1{`RANDOM}};
  rob_flits_returned_81 = _RAND_854[3:0];
  _RAND_855 = {1{`RANDOM}};
  rob_flits_returned_82 = _RAND_855[3:0];
  _RAND_856 = {1{`RANDOM}};
  rob_flits_returned_83 = _RAND_856[3:0];
  _RAND_857 = {1{`RANDOM}};
  rob_flits_returned_84 = _RAND_857[3:0];
  _RAND_858 = {1{`RANDOM}};
  rob_flits_returned_85 = _RAND_858[3:0];
  _RAND_859 = {1{`RANDOM}};
  rob_flits_returned_86 = _RAND_859[3:0];
  _RAND_860 = {1{`RANDOM}};
  rob_flits_returned_87 = _RAND_860[3:0];
  _RAND_861 = {1{`RANDOM}};
  rob_flits_returned_88 = _RAND_861[3:0];
  _RAND_862 = {1{`RANDOM}};
  rob_flits_returned_89 = _RAND_862[3:0];
  _RAND_863 = {1{`RANDOM}};
  rob_flits_returned_90 = _RAND_863[3:0];
  _RAND_864 = {1{`RANDOM}};
  rob_flits_returned_91 = _RAND_864[3:0];
  _RAND_865 = {1{`RANDOM}};
  rob_flits_returned_92 = _RAND_865[3:0];
  _RAND_866 = {1{`RANDOM}};
  rob_flits_returned_93 = _RAND_866[3:0];
  _RAND_867 = {1{`RANDOM}};
  rob_flits_returned_94 = _RAND_867[3:0];
  _RAND_868 = {1{`RANDOM}};
  rob_flits_returned_95 = _RAND_868[3:0];
  _RAND_869 = {1{`RANDOM}};
  rob_flits_returned_96 = _RAND_869[3:0];
  _RAND_870 = {1{`RANDOM}};
  rob_flits_returned_97 = _RAND_870[3:0];
  _RAND_871 = {1{`RANDOM}};
  rob_flits_returned_98 = _RAND_871[3:0];
  _RAND_872 = {1{`RANDOM}};
  rob_flits_returned_99 = _RAND_872[3:0];
  _RAND_873 = {1{`RANDOM}};
  rob_flits_returned_100 = _RAND_873[3:0];
  _RAND_874 = {1{`RANDOM}};
  rob_flits_returned_101 = _RAND_874[3:0];
  _RAND_875 = {1{`RANDOM}};
  rob_flits_returned_102 = _RAND_875[3:0];
  _RAND_876 = {1{`RANDOM}};
  rob_flits_returned_103 = _RAND_876[3:0];
  _RAND_877 = {1{`RANDOM}};
  rob_flits_returned_104 = _RAND_877[3:0];
  _RAND_878 = {1{`RANDOM}};
  rob_flits_returned_105 = _RAND_878[3:0];
  _RAND_879 = {1{`RANDOM}};
  rob_flits_returned_106 = _RAND_879[3:0];
  _RAND_880 = {1{`RANDOM}};
  rob_flits_returned_107 = _RAND_880[3:0];
  _RAND_881 = {1{`RANDOM}};
  rob_flits_returned_108 = _RAND_881[3:0];
  _RAND_882 = {1{`RANDOM}};
  rob_flits_returned_109 = _RAND_882[3:0];
  _RAND_883 = {1{`RANDOM}};
  rob_flits_returned_110 = _RAND_883[3:0];
  _RAND_884 = {1{`RANDOM}};
  rob_flits_returned_111 = _RAND_884[3:0];
  _RAND_885 = {1{`RANDOM}};
  rob_flits_returned_112 = _RAND_885[3:0];
  _RAND_886 = {1{`RANDOM}};
  rob_flits_returned_113 = _RAND_886[3:0];
  _RAND_887 = {1{`RANDOM}};
  rob_flits_returned_114 = _RAND_887[3:0];
  _RAND_888 = {1{`RANDOM}};
  rob_flits_returned_115 = _RAND_888[3:0];
  _RAND_889 = {1{`RANDOM}};
  rob_flits_returned_116 = _RAND_889[3:0];
  _RAND_890 = {1{`RANDOM}};
  rob_flits_returned_117 = _RAND_890[3:0];
  _RAND_891 = {1{`RANDOM}};
  rob_flits_returned_118 = _RAND_891[3:0];
  _RAND_892 = {1{`RANDOM}};
  rob_flits_returned_119 = _RAND_892[3:0];
  _RAND_893 = {1{`RANDOM}};
  rob_flits_returned_120 = _RAND_893[3:0];
  _RAND_894 = {1{`RANDOM}};
  rob_flits_returned_121 = _RAND_894[3:0];
  _RAND_895 = {1{`RANDOM}};
  rob_flits_returned_122 = _RAND_895[3:0];
  _RAND_896 = {1{`RANDOM}};
  rob_flits_returned_123 = _RAND_896[3:0];
  _RAND_897 = {1{`RANDOM}};
  rob_flits_returned_124 = _RAND_897[3:0];
  _RAND_898 = {1{`RANDOM}};
  rob_flits_returned_125 = _RAND_898[3:0];
  _RAND_899 = {1{`RANDOM}};
  rob_flits_returned_126 = _RAND_899[3:0];
  _RAND_900 = {1{`RANDOM}};
  rob_flits_returned_127 = _RAND_900[3:0];
  _RAND_901 = {2{`RANDOM}};
  rob_tscs_0 = _RAND_901[63:0];
  _RAND_902 = {2{`RANDOM}};
  rob_tscs_1 = _RAND_902[63:0];
  _RAND_903 = {2{`RANDOM}};
  rob_tscs_2 = _RAND_903[63:0];
  _RAND_904 = {2{`RANDOM}};
  rob_tscs_3 = _RAND_904[63:0];
  _RAND_905 = {2{`RANDOM}};
  rob_tscs_4 = _RAND_905[63:0];
  _RAND_906 = {2{`RANDOM}};
  rob_tscs_5 = _RAND_906[63:0];
  _RAND_907 = {2{`RANDOM}};
  rob_tscs_6 = _RAND_907[63:0];
  _RAND_908 = {2{`RANDOM}};
  rob_tscs_7 = _RAND_908[63:0];
  _RAND_909 = {2{`RANDOM}};
  rob_tscs_8 = _RAND_909[63:0];
  _RAND_910 = {2{`RANDOM}};
  rob_tscs_9 = _RAND_910[63:0];
  _RAND_911 = {2{`RANDOM}};
  rob_tscs_10 = _RAND_911[63:0];
  _RAND_912 = {2{`RANDOM}};
  rob_tscs_11 = _RAND_912[63:0];
  _RAND_913 = {2{`RANDOM}};
  rob_tscs_12 = _RAND_913[63:0];
  _RAND_914 = {2{`RANDOM}};
  rob_tscs_13 = _RAND_914[63:0];
  _RAND_915 = {2{`RANDOM}};
  rob_tscs_14 = _RAND_915[63:0];
  _RAND_916 = {2{`RANDOM}};
  rob_tscs_15 = _RAND_916[63:0];
  _RAND_917 = {2{`RANDOM}};
  rob_tscs_16 = _RAND_917[63:0];
  _RAND_918 = {2{`RANDOM}};
  rob_tscs_17 = _RAND_918[63:0];
  _RAND_919 = {2{`RANDOM}};
  rob_tscs_18 = _RAND_919[63:0];
  _RAND_920 = {2{`RANDOM}};
  rob_tscs_19 = _RAND_920[63:0];
  _RAND_921 = {2{`RANDOM}};
  rob_tscs_20 = _RAND_921[63:0];
  _RAND_922 = {2{`RANDOM}};
  rob_tscs_21 = _RAND_922[63:0];
  _RAND_923 = {2{`RANDOM}};
  rob_tscs_22 = _RAND_923[63:0];
  _RAND_924 = {2{`RANDOM}};
  rob_tscs_23 = _RAND_924[63:0];
  _RAND_925 = {2{`RANDOM}};
  rob_tscs_24 = _RAND_925[63:0];
  _RAND_926 = {2{`RANDOM}};
  rob_tscs_25 = _RAND_926[63:0];
  _RAND_927 = {2{`RANDOM}};
  rob_tscs_26 = _RAND_927[63:0];
  _RAND_928 = {2{`RANDOM}};
  rob_tscs_27 = _RAND_928[63:0];
  _RAND_929 = {2{`RANDOM}};
  rob_tscs_28 = _RAND_929[63:0];
  _RAND_930 = {2{`RANDOM}};
  rob_tscs_29 = _RAND_930[63:0];
  _RAND_931 = {2{`RANDOM}};
  rob_tscs_30 = _RAND_931[63:0];
  _RAND_932 = {2{`RANDOM}};
  rob_tscs_31 = _RAND_932[63:0];
  _RAND_933 = {2{`RANDOM}};
  rob_tscs_32 = _RAND_933[63:0];
  _RAND_934 = {2{`RANDOM}};
  rob_tscs_33 = _RAND_934[63:0];
  _RAND_935 = {2{`RANDOM}};
  rob_tscs_34 = _RAND_935[63:0];
  _RAND_936 = {2{`RANDOM}};
  rob_tscs_35 = _RAND_936[63:0];
  _RAND_937 = {2{`RANDOM}};
  rob_tscs_36 = _RAND_937[63:0];
  _RAND_938 = {2{`RANDOM}};
  rob_tscs_37 = _RAND_938[63:0];
  _RAND_939 = {2{`RANDOM}};
  rob_tscs_38 = _RAND_939[63:0];
  _RAND_940 = {2{`RANDOM}};
  rob_tscs_39 = _RAND_940[63:0];
  _RAND_941 = {2{`RANDOM}};
  rob_tscs_40 = _RAND_941[63:0];
  _RAND_942 = {2{`RANDOM}};
  rob_tscs_41 = _RAND_942[63:0];
  _RAND_943 = {2{`RANDOM}};
  rob_tscs_42 = _RAND_943[63:0];
  _RAND_944 = {2{`RANDOM}};
  rob_tscs_43 = _RAND_944[63:0];
  _RAND_945 = {2{`RANDOM}};
  rob_tscs_44 = _RAND_945[63:0];
  _RAND_946 = {2{`RANDOM}};
  rob_tscs_45 = _RAND_946[63:0];
  _RAND_947 = {2{`RANDOM}};
  rob_tscs_46 = _RAND_947[63:0];
  _RAND_948 = {2{`RANDOM}};
  rob_tscs_47 = _RAND_948[63:0];
  _RAND_949 = {2{`RANDOM}};
  rob_tscs_48 = _RAND_949[63:0];
  _RAND_950 = {2{`RANDOM}};
  rob_tscs_49 = _RAND_950[63:0];
  _RAND_951 = {2{`RANDOM}};
  rob_tscs_50 = _RAND_951[63:0];
  _RAND_952 = {2{`RANDOM}};
  rob_tscs_51 = _RAND_952[63:0];
  _RAND_953 = {2{`RANDOM}};
  rob_tscs_52 = _RAND_953[63:0];
  _RAND_954 = {2{`RANDOM}};
  rob_tscs_53 = _RAND_954[63:0];
  _RAND_955 = {2{`RANDOM}};
  rob_tscs_54 = _RAND_955[63:0];
  _RAND_956 = {2{`RANDOM}};
  rob_tscs_55 = _RAND_956[63:0];
  _RAND_957 = {2{`RANDOM}};
  rob_tscs_56 = _RAND_957[63:0];
  _RAND_958 = {2{`RANDOM}};
  rob_tscs_57 = _RAND_958[63:0];
  _RAND_959 = {2{`RANDOM}};
  rob_tscs_58 = _RAND_959[63:0];
  _RAND_960 = {2{`RANDOM}};
  rob_tscs_59 = _RAND_960[63:0];
  _RAND_961 = {2{`RANDOM}};
  rob_tscs_60 = _RAND_961[63:0];
  _RAND_962 = {2{`RANDOM}};
  rob_tscs_61 = _RAND_962[63:0];
  _RAND_963 = {2{`RANDOM}};
  rob_tscs_62 = _RAND_963[63:0];
  _RAND_964 = {2{`RANDOM}};
  rob_tscs_63 = _RAND_964[63:0];
  _RAND_965 = {2{`RANDOM}};
  rob_tscs_64 = _RAND_965[63:0];
  _RAND_966 = {2{`RANDOM}};
  rob_tscs_65 = _RAND_966[63:0];
  _RAND_967 = {2{`RANDOM}};
  rob_tscs_66 = _RAND_967[63:0];
  _RAND_968 = {2{`RANDOM}};
  rob_tscs_67 = _RAND_968[63:0];
  _RAND_969 = {2{`RANDOM}};
  rob_tscs_68 = _RAND_969[63:0];
  _RAND_970 = {2{`RANDOM}};
  rob_tscs_69 = _RAND_970[63:0];
  _RAND_971 = {2{`RANDOM}};
  rob_tscs_70 = _RAND_971[63:0];
  _RAND_972 = {2{`RANDOM}};
  rob_tscs_71 = _RAND_972[63:0];
  _RAND_973 = {2{`RANDOM}};
  rob_tscs_72 = _RAND_973[63:0];
  _RAND_974 = {2{`RANDOM}};
  rob_tscs_73 = _RAND_974[63:0];
  _RAND_975 = {2{`RANDOM}};
  rob_tscs_74 = _RAND_975[63:0];
  _RAND_976 = {2{`RANDOM}};
  rob_tscs_75 = _RAND_976[63:0];
  _RAND_977 = {2{`RANDOM}};
  rob_tscs_76 = _RAND_977[63:0];
  _RAND_978 = {2{`RANDOM}};
  rob_tscs_77 = _RAND_978[63:0];
  _RAND_979 = {2{`RANDOM}};
  rob_tscs_78 = _RAND_979[63:0];
  _RAND_980 = {2{`RANDOM}};
  rob_tscs_79 = _RAND_980[63:0];
  _RAND_981 = {2{`RANDOM}};
  rob_tscs_80 = _RAND_981[63:0];
  _RAND_982 = {2{`RANDOM}};
  rob_tscs_81 = _RAND_982[63:0];
  _RAND_983 = {2{`RANDOM}};
  rob_tscs_82 = _RAND_983[63:0];
  _RAND_984 = {2{`RANDOM}};
  rob_tscs_83 = _RAND_984[63:0];
  _RAND_985 = {2{`RANDOM}};
  rob_tscs_84 = _RAND_985[63:0];
  _RAND_986 = {2{`RANDOM}};
  rob_tscs_85 = _RAND_986[63:0];
  _RAND_987 = {2{`RANDOM}};
  rob_tscs_86 = _RAND_987[63:0];
  _RAND_988 = {2{`RANDOM}};
  rob_tscs_87 = _RAND_988[63:0];
  _RAND_989 = {2{`RANDOM}};
  rob_tscs_88 = _RAND_989[63:0];
  _RAND_990 = {2{`RANDOM}};
  rob_tscs_89 = _RAND_990[63:0];
  _RAND_991 = {2{`RANDOM}};
  rob_tscs_90 = _RAND_991[63:0];
  _RAND_992 = {2{`RANDOM}};
  rob_tscs_91 = _RAND_992[63:0];
  _RAND_993 = {2{`RANDOM}};
  rob_tscs_92 = _RAND_993[63:0];
  _RAND_994 = {2{`RANDOM}};
  rob_tscs_93 = _RAND_994[63:0];
  _RAND_995 = {2{`RANDOM}};
  rob_tscs_94 = _RAND_995[63:0];
  _RAND_996 = {2{`RANDOM}};
  rob_tscs_95 = _RAND_996[63:0];
  _RAND_997 = {2{`RANDOM}};
  rob_tscs_96 = _RAND_997[63:0];
  _RAND_998 = {2{`RANDOM}};
  rob_tscs_97 = _RAND_998[63:0];
  _RAND_999 = {2{`RANDOM}};
  rob_tscs_98 = _RAND_999[63:0];
  _RAND_1000 = {2{`RANDOM}};
  rob_tscs_99 = _RAND_1000[63:0];
  _RAND_1001 = {2{`RANDOM}};
  rob_tscs_100 = _RAND_1001[63:0];
  _RAND_1002 = {2{`RANDOM}};
  rob_tscs_101 = _RAND_1002[63:0];
  _RAND_1003 = {2{`RANDOM}};
  rob_tscs_102 = _RAND_1003[63:0];
  _RAND_1004 = {2{`RANDOM}};
  rob_tscs_103 = _RAND_1004[63:0];
  _RAND_1005 = {2{`RANDOM}};
  rob_tscs_104 = _RAND_1005[63:0];
  _RAND_1006 = {2{`RANDOM}};
  rob_tscs_105 = _RAND_1006[63:0];
  _RAND_1007 = {2{`RANDOM}};
  rob_tscs_106 = _RAND_1007[63:0];
  _RAND_1008 = {2{`RANDOM}};
  rob_tscs_107 = _RAND_1008[63:0];
  _RAND_1009 = {2{`RANDOM}};
  rob_tscs_108 = _RAND_1009[63:0];
  _RAND_1010 = {2{`RANDOM}};
  rob_tscs_109 = _RAND_1010[63:0];
  _RAND_1011 = {2{`RANDOM}};
  rob_tscs_110 = _RAND_1011[63:0];
  _RAND_1012 = {2{`RANDOM}};
  rob_tscs_111 = _RAND_1012[63:0];
  _RAND_1013 = {2{`RANDOM}};
  rob_tscs_112 = _RAND_1013[63:0];
  _RAND_1014 = {2{`RANDOM}};
  rob_tscs_113 = _RAND_1014[63:0];
  _RAND_1015 = {2{`RANDOM}};
  rob_tscs_114 = _RAND_1015[63:0];
  _RAND_1016 = {2{`RANDOM}};
  rob_tscs_115 = _RAND_1016[63:0];
  _RAND_1017 = {2{`RANDOM}};
  rob_tscs_116 = _RAND_1017[63:0];
  _RAND_1018 = {2{`RANDOM}};
  rob_tscs_117 = _RAND_1018[63:0];
  _RAND_1019 = {2{`RANDOM}};
  rob_tscs_118 = _RAND_1019[63:0];
  _RAND_1020 = {2{`RANDOM}};
  rob_tscs_119 = _RAND_1020[63:0];
  _RAND_1021 = {2{`RANDOM}};
  rob_tscs_120 = _RAND_1021[63:0];
  _RAND_1022 = {2{`RANDOM}};
  rob_tscs_121 = _RAND_1022[63:0];
  _RAND_1023 = {2{`RANDOM}};
  rob_tscs_122 = _RAND_1023[63:0];
  _RAND_1024 = {2{`RANDOM}};
  rob_tscs_123 = _RAND_1024[63:0];
  _RAND_1025 = {2{`RANDOM}};
  rob_tscs_124 = _RAND_1025[63:0];
  _RAND_1026 = {2{`RANDOM}};
  rob_tscs_125 = _RAND_1026[63:0];
  _RAND_1027 = {2{`RANDOM}};
  rob_tscs_126 = _RAND_1027[63:0];
  _RAND_1028 = {2{`RANDOM}};
  rob_tscs_127 = _RAND_1028[63:0];
  _RAND_1029 = {1{`RANDOM}};
  io_success_REG = _RAND_1029[0:0];
  _RAND_1030 = {1{`RANDOM}};
  packet_valid = _RAND_1030[0:0];
  _RAND_1031 = {1{`RANDOM}};
  packet_rob_idx = _RAND_1031[6:0];
  _RAND_1032 = {1{`RANDOM}};
  packet_valid_1 = _RAND_1032[0:0];
  _RAND_1033 = {1{`RANDOM}};
  packet_rob_idx_1 = _RAND_1033[6:0];
  _RAND_1034 = {1{`RANDOM}};
  packet_valid_2 = _RAND_1034[0:0];
  _RAND_1035 = {1{`RANDOM}};
  packet_rob_idx_2 = _RAND_1035[6:0];
  _RAND_1036 = {1{`RANDOM}};
  packet_valid_3 = _RAND_1036[0:0];
  _RAND_1037 = {1{`RANDOM}};
  packet_rob_idx_3 = _RAND_1037[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(~idle_counter[10]); // @[TestHarness.scala 148:9]
    end
    //
    if (_T_118 & _T_3) begin
      assert(_T_76[0]); // @[TestHarness.scala 201:13]
    end
    //
    if (_T_118 & _T_3) begin
      assert(_T_82 == io_from_noc_0_flit_bits_payload); // @[TestHarness.scala 202:13]
    end
    //
    if (_T_118 & _T_3) begin
      assert(io_from_noc_0_flit_bits_ingress_id == _GEN_8704); // @[TestHarness.scala 203:13]
    end
    //
    if (_T_118 & _T_3) begin
      assert(2'h0 == _GEN_8832); // @[TestHarness.scala 204:13]
    end
    //
    if (_T_118 & _T_3) begin
      assert(_GEN_8960 < _GEN_9088); // @[TestHarness.scala 205:13]
    end
    //
    if (_T_118 & _T_3) begin
      assert(~packet_valid & io_from_noc_0_flit_bits_head | out_payload_rob_idx == _GEN_15381); // @[TestHarness.scala 206:13]
    end
    //
    if (_T_165 & _T_3) begin
      assert(_T_123[0]); // @[TestHarness.scala 201:13]
    end
    //
    if (_T_165 & _T_3) begin
      assert(_T_129 == io_from_noc_1_flit_bits_payload); // @[TestHarness.scala 202:13]
    end
    //
    if (_T_165 & _T_3) begin
      assert(io_from_noc_1_flit_bits_ingress_id == _GEN_10501); // @[TestHarness.scala 203:13]
    end
    //
    if (_T_165 & _T_3) begin
      assert(2'h1 == _GEN_10629); // @[TestHarness.scala 204:13]
    end
    //
    if (_T_165 & _T_3) begin
      assert(_GEN_10757 < _GEN_10885); // @[TestHarness.scala 205:13]
    end
    //
    if (_T_165 & _T_3) begin
      assert(~packet_valid_1 & io_from_noc_1_flit_bits_head | out_payload_1_rob_idx == _GEN_15382); // @[TestHarness.scala 206:13]
    end
    //
    if (_T_212 & _T_3) begin
      assert(_T_170[0]); // @[TestHarness.scala 201:13]
    end
    //
    if (_T_212 & _T_3) begin
      assert(_T_176 == io_from_noc_2_flit_bits_payload); // @[TestHarness.scala 202:13]
    end
    //
    if (_T_212 & _T_3) begin
      assert(io_from_noc_2_flit_bits_ingress_id == _GEN_12298); // @[TestHarness.scala 203:13]
    end
    //
    if (_T_212 & _T_3) begin
      assert(2'h2 == _GEN_12426); // @[TestHarness.scala 204:13]
    end
    //
    if (_T_212 & _T_3) begin
      assert(_GEN_12554 < _GEN_12682); // @[TestHarness.scala 205:13]
    end
    //
    if (_T_212 & _T_3) begin
      assert(~packet_valid_2 & io_from_noc_2_flit_bits_head | out_payload_2_rob_idx == _GEN_15383); // @[TestHarness.scala 206:13]
    end
    //
    if (_T_259 & _T_3) begin
      assert(_T_217[0]); // @[TestHarness.scala 201:13]
    end
    //
    if (_T_259 & _T_3) begin
      assert(_T_223 == io_from_noc_3_flit_bits_payload); // @[TestHarness.scala 202:13]
    end
    //
    if (_T_259 & _T_3) begin
      assert(io_from_noc_3_flit_bits_ingress_id == _GEN_14095); // @[TestHarness.scala 203:13]
    end
    //
    if (_T_259 & _T_3) begin
      assert(2'h3 == _GEN_14223); // @[TestHarness.scala 204:13]
    end
    //
    if (_T_259 & _T_3) begin
      assert(_GEN_14351 < _GEN_14479); // @[TestHarness.scala 205:13]
    end
    //
    if (_T_259 & _T_3) begin
      assert(~packet_valid_3 & io_from_noc_3_flit_bits_head | out_payload_3_rob_idx == _GEN_15384); // @[TestHarness.scala 206:13]
    end
    //
    if (rob_valids[0] & _T_3) begin
      assert(_T_264 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[1] & _T_3) begin
      assert(_T_271 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[2] & _T_3) begin
      assert(_T_278 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[3] & _T_3) begin
      assert(_T_285 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[4] & _T_3) begin
      assert(_T_292 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[5] & _T_3) begin
      assert(_T_299 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[6] & _T_3) begin
      assert(_T_306 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[7] & _T_3) begin
      assert(_T_313 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[8] & _T_3) begin
      assert(_T_320 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[9] & _T_3) begin
      assert(_T_327 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[10] & _T_3) begin
      assert(_T_334 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[11] & _T_3) begin
      assert(_T_341 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[12] & _T_3) begin
      assert(_T_348 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[13] & _T_3) begin
      assert(_T_355 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[14] & _T_3) begin
      assert(_T_362 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[15] & _T_3) begin
      assert(_T_369 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[16] & _T_3) begin
      assert(_T_376 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[17] & _T_3) begin
      assert(_T_383 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[18] & _T_3) begin
      assert(_T_390 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[19] & _T_3) begin
      assert(_T_397 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[20] & _T_3) begin
      assert(_T_404 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[21] & _T_3) begin
      assert(_T_411 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[22] & _T_3) begin
      assert(_T_418 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[23] & _T_3) begin
      assert(_T_425 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[24] & _T_3) begin
      assert(_T_432 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[25] & _T_3) begin
      assert(_T_439 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[26] & _T_3) begin
      assert(_T_446 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[27] & _T_3) begin
      assert(_T_453 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[28] & _T_3) begin
      assert(_T_460 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[29] & _T_3) begin
      assert(_T_467 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[30] & _T_3) begin
      assert(_T_474 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[31] & _T_3) begin
      assert(_T_481 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[32] & _T_3) begin
      assert(_T_488 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[33] & _T_3) begin
      assert(_T_495 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[34] & _T_3) begin
      assert(_T_502 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[35] & _T_3) begin
      assert(_T_509 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[36] & _T_3) begin
      assert(_T_516 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[37] & _T_3) begin
      assert(_T_523 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[38] & _T_3) begin
      assert(_T_530 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[39] & _T_3) begin
      assert(_T_537 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[40] & _T_3) begin
      assert(_T_544 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[41] & _T_3) begin
      assert(_T_551 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[42] & _T_3) begin
      assert(_T_558 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[43] & _T_3) begin
      assert(_T_565 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[44] & _T_3) begin
      assert(_T_572 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[45] & _T_3) begin
      assert(_T_579 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[46] & _T_3) begin
      assert(_T_586 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[47] & _T_3) begin
      assert(_T_593 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[48] & _T_3) begin
      assert(_T_600 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[49] & _T_3) begin
      assert(_T_607 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[50] & _T_3) begin
      assert(_T_614 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[51] & _T_3) begin
      assert(_T_621 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[52] & _T_3) begin
      assert(_T_628 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[53] & _T_3) begin
      assert(_T_635 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[54] & _T_3) begin
      assert(_T_642 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[55] & _T_3) begin
      assert(_T_649 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[56] & _T_3) begin
      assert(_T_656 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[57] & _T_3) begin
      assert(_T_663 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[58] & _T_3) begin
      assert(_T_670 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[59] & _T_3) begin
      assert(_T_677 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[60] & _T_3) begin
      assert(_T_684 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[61] & _T_3) begin
      assert(_T_691 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[62] & _T_3) begin
      assert(_T_698 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[63] & _T_3) begin
      assert(_T_705 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[64] & _T_3) begin
      assert(_T_712 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[65] & _T_3) begin
      assert(_T_719 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[66] & _T_3) begin
      assert(_T_726 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[67] & _T_3) begin
      assert(_T_733 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[68] & _T_3) begin
      assert(_T_740 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[69] & _T_3) begin
      assert(_T_747 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[70] & _T_3) begin
      assert(_T_754 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[71] & _T_3) begin
      assert(_T_761 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[72] & _T_3) begin
      assert(_T_768 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[73] & _T_3) begin
      assert(_T_775 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[74] & _T_3) begin
      assert(_T_782 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[75] & _T_3) begin
      assert(_T_789 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[76] & _T_3) begin
      assert(_T_796 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[77] & _T_3) begin
      assert(_T_803 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[78] & _T_3) begin
      assert(_T_810 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[79] & _T_3) begin
      assert(_T_817 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[80] & _T_3) begin
      assert(_T_824 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[81] & _T_3) begin
      assert(_T_831 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[82] & _T_3) begin
      assert(_T_838 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[83] & _T_3) begin
      assert(_T_845 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[84] & _T_3) begin
      assert(_T_852 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[85] & _T_3) begin
      assert(_T_859 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[86] & _T_3) begin
      assert(_T_866 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[87] & _T_3) begin
      assert(_T_873 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[88] & _T_3) begin
      assert(_T_880 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[89] & _T_3) begin
      assert(_T_887 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[90] & _T_3) begin
      assert(_T_894 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[91] & _T_3) begin
      assert(_T_901 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[92] & _T_3) begin
      assert(_T_908 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[93] & _T_3) begin
      assert(_T_915 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[94] & _T_3) begin
      assert(_T_922 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[95] & _T_3) begin
      assert(_T_929 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[96] & _T_3) begin
      assert(_T_936 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[97] & _T_3) begin
      assert(_T_943 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[98] & _T_3) begin
      assert(_T_950 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[99] & _T_3) begin
      assert(_T_957 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[100] & _T_3) begin
      assert(_T_964 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[101] & _T_3) begin
      assert(_T_971 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[102] & _T_3) begin
      assert(_T_978 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[103] & _T_3) begin
      assert(_T_985 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[104] & _T_3) begin
      assert(_T_992 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[105] & _T_3) begin
      assert(_T_999 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[106] & _T_3) begin
      assert(_T_1006 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[107] & _T_3) begin
      assert(_T_1013 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[108] & _T_3) begin
      assert(_T_1020 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[109] & _T_3) begin
      assert(_T_1027 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[110] & _T_3) begin
      assert(_T_1034 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[111] & _T_3) begin
      assert(_T_1041 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[112] & _T_3) begin
      assert(_T_1048 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[113] & _T_3) begin
      assert(_T_1055 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[114] & _T_3) begin
      assert(_T_1062 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[115] & _T_3) begin
      assert(_T_1069 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[116] & _T_3) begin
      assert(_T_1076 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[117] & _T_3) begin
      assert(_T_1083 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[118] & _T_3) begin
      assert(_T_1090 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[119] & _T_3) begin
      assert(_T_1097 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[120] & _T_3) begin
      assert(_T_1104 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[121] & _T_3) begin
      assert(_T_1111 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[122] & _T_3) begin
      assert(_T_1118 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[123] & _T_3) begin
      assert(_T_1125 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[124] & _T_3) begin
      assert(_T_1132 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[125] & _T_3) begin
      assert(_T_1139 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[126] & _T_3) begin
      assert(_T_1146 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[127] & _T_3) begin
      assert(_T_1153 < 64'h4000); // @[TestHarness.scala 229:13]
    end
  end
endmodule
module TestHarness(
  input   clock,
  input   reset,
  output  io_success
);
  wire  lazyNoC_clock; // @[TestHarness.scala 238:19]
  wire  lazyNoC_reset; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_ingress_3_flit_ready; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_ingress_3_flit_valid; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_ingress_3_flit_bits_head; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_ingress_3_flit_bits_tail; // @[TestHarness.scala 238:19]
  wire [63:0] lazyNoC_io_ingress_3_flit_bits_payload; // @[TestHarness.scala 238:19]
  wire [1:0] lazyNoC_io_ingress_3_flit_bits_egress_id; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_ingress_2_flit_ready; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_ingress_2_flit_valid; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_ingress_2_flit_bits_head; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_ingress_2_flit_bits_tail; // @[TestHarness.scala 238:19]
  wire [63:0] lazyNoC_io_ingress_2_flit_bits_payload; // @[TestHarness.scala 238:19]
  wire [1:0] lazyNoC_io_ingress_2_flit_bits_egress_id; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_ingress_1_flit_ready; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_ingress_1_flit_valid; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_ingress_1_flit_bits_head; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_ingress_1_flit_bits_tail; // @[TestHarness.scala 238:19]
  wire [63:0] lazyNoC_io_ingress_1_flit_bits_payload; // @[TestHarness.scala 238:19]
  wire [1:0] lazyNoC_io_ingress_1_flit_bits_egress_id; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_ingress_0_flit_ready; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_ingress_0_flit_valid; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_ingress_0_flit_bits_head; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_ingress_0_flit_bits_tail; // @[TestHarness.scala 238:19]
  wire [63:0] lazyNoC_io_ingress_0_flit_bits_payload; // @[TestHarness.scala 238:19]
  wire [1:0] lazyNoC_io_ingress_0_flit_bits_egress_id; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_egress_3_flit_valid; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_egress_3_flit_bits_head; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_egress_3_flit_bits_tail; // @[TestHarness.scala 238:19]
  wire [63:0] lazyNoC_io_egress_3_flit_bits_payload; // @[TestHarness.scala 238:19]
  wire [1:0] lazyNoC_io_egress_3_flit_bits_ingress_id; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_egress_2_flit_valid; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_egress_2_flit_bits_head; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_egress_2_flit_bits_tail; // @[TestHarness.scala 238:19]
  wire [63:0] lazyNoC_io_egress_2_flit_bits_payload; // @[TestHarness.scala 238:19]
  wire [1:0] lazyNoC_io_egress_2_flit_bits_ingress_id; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_egress_1_flit_valid; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_egress_1_flit_bits_head; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_egress_1_flit_bits_tail; // @[TestHarness.scala 238:19]
  wire [63:0] lazyNoC_io_egress_1_flit_bits_payload; // @[TestHarness.scala 238:19]
  wire [1:0] lazyNoC_io_egress_1_flit_bits_ingress_id; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_egress_0_flit_valid; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_egress_0_flit_bits_head; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_egress_0_flit_bits_tail; // @[TestHarness.scala 238:19]
  wire [63:0] lazyNoC_io_egress_0_flit_bits_payload; // @[TestHarness.scala 238:19]
  wire [1:0] lazyNoC_io_egress_0_flit_bits_ingress_id; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_router_clocks_0_clock; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_router_clocks_0_reset; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_router_clocks_1_clock; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_router_clocks_1_reset; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_router_clocks_2_clock; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_router_clocks_2_reset; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_router_clocks_3_clock; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_router_clocks_3_reset; // @[TestHarness.scala 238:19]
  wire  noc_tester_clock; // @[TestHarness.scala 269:26]
  wire  noc_tester_reset; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_to_noc_3_flit_ready; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_to_noc_3_flit_valid; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_to_noc_3_flit_bits_head; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_to_noc_3_flit_bits_tail; // @[TestHarness.scala 269:26]
  wire [63:0] noc_tester_io_to_noc_3_flit_bits_payload; // @[TestHarness.scala 269:26]
  wire [1:0] noc_tester_io_to_noc_3_flit_bits_egress_id; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_to_noc_2_flit_ready; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_to_noc_2_flit_valid; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_to_noc_2_flit_bits_head; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_to_noc_2_flit_bits_tail; // @[TestHarness.scala 269:26]
  wire [63:0] noc_tester_io_to_noc_2_flit_bits_payload; // @[TestHarness.scala 269:26]
  wire [1:0] noc_tester_io_to_noc_2_flit_bits_egress_id; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_to_noc_1_flit_ready; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_to_noc_1_flit_valid; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_to_noc_1_flit_bits_head; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_to_noc_1_flit_bits_tail; // @[TestHarness.scala 269:26]
  wire [63:0] noc_tester_io_to_noc_1_flit_bits_payload; // @[TestHarness.scala 269:26]
  wire [1:0] noc_tester_io_to_noc_1_flit_bits_egress_id; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_to_noc_0_flit_ready; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_to_noc_0_flit_valid; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_to_noc_0_flit_bits_head; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_to_noc_0_flit_bits_tail; // @[TestHarness.scala 269:26]
  wire [63:0] noc_tester_io_to_noc_0_flit_bits_payload; // @[TestHarness.scala 269:26]
  wire [1:0] noc_tester_io_to_noc_0_flit_bits_egress_id; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_from_noc_3_flit_ready; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_from_noc_3_flit_valid; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_from_noc_3_flit_bits_head; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_from_noc_3_flit_bits_tail; // @[TestHarness.scala 269:26]
  wire [63:0] noc_tester_io_from_noc_3_flit_bits_payload; // @[TestHarness.scala 269:26]
  wire [1:0] noc_tester_io_from_noc_3_flit_bits_ingress_id; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_from_noc_2_flit_ready; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_from_noc_2_flit_valid; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_from_noc_2_flit_bits_head; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_from_noc_2_flit_bits_tail; // @[TestHarness.scala 269:26]
  wire [63:0] noc_tester_io_from_noc_2_flit_bits_payload; // @[TestHarness.scala 269:26]
  wire [1:0] noc_tester_io_from_noc_2_flit_bits_ingress_id; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_from_noc_1_flit_ready; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_from_noc_1_flit_valid; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_from_noc_1_flit_bits_head; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_from_noc_1_flit_bits_tail; // @[TestHarness.scala 269:26]
  wire [63:0] noc_tester_io_from_noc_1_flit_bits_payload; // @[TestHarness.scala 269:26]
  wire [1:0] noc_tester_io_from_noc_1_flit_bits_ingress_id; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_from_noc_0_flit_ready; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_from_noc_0_flit_valid; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_from_noc_0_flit_bits_head; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_from_noc_0_flit_bits_tail; // @[TestHarness.scala 269:26]
  wire [63:0] noc_tester_io_from_noc_0_flit_bits_payload; // @[TestHarness.scala 269:26]
  wire [1:0] noc_tester_io_from_noc_0_flit_bits_ingress_id; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_success; // @[TestHarness.scala 269:26]
  NoC lazyNoC ( // @[TestHarness.scala 238:19]
    .clock(lazyNoC_clock),
    .reset(lazyNoC_reset),
    .io_ingress_3_flit_ready(lazyNoC_io_ingress_3_flit_ready),
    .io_ingress_3_flit_valid(lazyNoC_io_ingress_3_flit_valid),
    .io_ingress_3_flit_bits_head(lazyNoC_io_ingress_3_flit_bits_head),
    .io_ingress_3_flit_bits_tail(lazyNoC_io_ingress_3_flit_bits_tail),
    .io_ingress_3_flit_bits_payload(lazyNoC_io_ingress_3_flit_bits_payload),
    .io_ingress_3_flit_bits_egress_id(lazyNoC_io_ingress_3_flit_bits_egress_id),
    .io_ingress_2_flit_ready(lazyNoC_io_ingress_2_flit_ready),
    .io_ingress_2_flit_valid(lazyNoC_io_ingress_2_flit_valid),
    .io_ingress_2_flit_bits_head(lazyNoC_io_ingress_2_flit_bits_head),
    .io_ingress_2_flit_bits_tail(lazyNoC_io_ingress_2_flit_bits_tail),
    .io_ingress_2_flit_bits_payload(lazyNoC_io_ingress_2_flit_bits_payload),
    .io_ingress_2_flit_bits_egress_id(lazyNoC_io_ingress_2_flit_bits_egress_id),
    .io_ingress_1_flit_ready(lazyNoC_io_ingress_1_flit_ready),
    .io_ingress_1_flit_valid(lazyNoC_io_ingress_1_flit_valid),
    .io_ingress_1_flit_bits_head(lazyNoC_io_ingress_1_flit_bits_head),
    .io_ingress_1_flit_bits_tail(lazyNoC_io_ingress_1_flit_bits_tail),
    .io_ingress_1_flit_bits_payload(lazyNoC_io_ingress_1_flit_bits_payload),
    .io_ingress_1_flit_bits_egress_id(lazyNoC_io_ingress_1_flit_bits_egress_id),
    .io_ingress_0_flit_ready(lazyNoC_io_ingress_0_flit_ready),
    .io_ingress_0_flit_valid(lazyNoC_io_ingress_0_flit_valid),
    .io_ingress_0_flit_bits_head(lazyNoC_io_ingress_0_flit_bits_head),
    .io_ingress_0_flit_bits_tail(lazyNoC_io_ingress_0_flit_bits_tail),
    .io_ingress_0_flit_bits_payload(lazyNoC_io_ingress_0_flit_bits_payload),
    .io_ingress_0_flit_bits_egress_id(lazyNoC_io_ingress_0_flit_bits_egress_id),
    .io_egress_3_flit_valid(lazyNoC_io_egress_3_flit_valid),
    .io_egress_3_flit_bits_head(lazyNoC_io_egress_3_flit_bits_head),
    .io_egress_3_flit_bits_tail(lazyNoC_io_egress_3_flit_bits_tail),
    .io_egress_3_flit_bits_payload(lazyNoC_io_egress_3_flit_bits_payload),
    .io_egress_3_flit_bits_ingress_id(lazyNoC_io_egress_3_flit_bits_ingress_id),
    .io_egress_2_flit_valid(lazyNoC_io_egress_2_flit_valid),
    .io_egress_2_flit_bits_head(lazyNoC_io_egress_2_flit_bits_head),
    .io_egress_2_flit_bits_tail(lazyNoC_io_egress_2_flit_bits_tail),
    .io_egress_2_flit_bits_payload(lazyNoC_io_egress_2_flit_bits_payload),
    .io_egress_2_flit_bits_ingress_id(lazyNoC_io_egress_2_flit_bits_ingress_id),
    .io_egress_1_flit_valid(lazyNoC_io_egress_1_flit_valid),
    .io_egress_1_flit_bits_head(lazyNoC_io_egress_1_flit_bits_head),
    .io_egress_1_flit_bits_tail(lazyNoC_io_egress_1_flit_bits_tail),
    .io_egress_1_flit_bits_payload(lazyNoC_io_egress_1_flit_bits_payload),
    .io_egress_1_flit_bits_ingress_id(lazyNoC_io_egress_1_flit_bits_ingress_id),
    .io_egress_0_flit_valid(lazyNoC_io_egress_0_flit_valid),
    .io_egress_0_flit_bits_head(lazyNoC_io_egress_0_flit_bits_head),
    .io_egress_0_flit_bits_tail(lazyNoC_io_egress_0_flit_bits_tail),
    .io_egress_0_flit_bits_payload(lazyNoC_io_egress_0_flit_bits_payload),
    .io_egress_0_flit_bits_ingress_id(lazyNoC_io_egress_0_flit_bits_ingress_id),
    .io_router_clocks_0_clock(lazyNoC_io_router_clocks_0_clock),
    .io_router_clocks_0_reset(lazyNoC_io_router_clocks_0_reset),
    .io_router_clocks_1_clock(lazyNoC_io_router_clocks_1_clock),
    .io_router_clocks_1_reset(lazyNoC_io_router_clocks_1_reset),
    .io_router_clocks_2_clock(lazyNoC_io_router_clocks_2_clock),
    .io_router_clocks_2_reset(lazyNoC_io_router_clocks_2_reset),
    .io_router_clocks_3_clock(lazyNoC_io_router_clocks_3_clock),
    .io_router_clocks_3_reset(lazyNoC_io_router_clocks_3_reset)
  );
  NoCTester noc_tester ( // @[TestHarness.scala 269:26]
    .clock(noc_tester_clock),
    .reset(noc_tester_reset),
    .io_to_noc_3_flit_ready(noc_tester_io_to_noc_3_flit_ready),
    .io_to_noc_3_flit_valid(noc_tester_io_to_noc_3_flit_valid),
    .io_to_noc_3_flit_bits_head(noc_tester_io_to_noc_3_flit_bits_head),
    .io_to_noc_3_flit_bits_tail(noc_tester_io_to_noc_3_flit_bits_tail),
    .io_to_noc_3_flit_bits_payload(noc_tester_io_to_noc_3_flit_bits_payload),
    .io_to_noc_3_flit_bits_egress_id(noc_tester_io_to_noc_3_flit_bits_egress_id),
    .io_to_noc_2_flit_ready(noc_tester_io_to_noc_2_flit_ready),
    .io_to_noc_2_flit_valid(noc_tester_io_to_noc_2_flit_valid),
    .io_to_noc_2_flit_bits_head(noc_tester_io_to_noc_2_flit_bits_head),
    .io_to_noc_2_flit_bits_tail(noc_tester_io_to_noc_2_flit_bits_tail),
    .io_to_noc_2_flit_bits_payload(noc_tester_io_to_noc_2_flit_bits_payload),
    .io_to_noc_2_flit_bits_egress_id(noc_tester_io_to_noc_2_flit_bits_egress_id),
    .io_to_noc_1_flit_ready(noc_tester_io_to_noc_1_flit_ready),
    .io_to_noc_1_flit_valid(noc_tester_io_to_noc_1_flit_valid),
    .io_to_noc_1_flit_bits_head(noc_tester_io_to_noc_1_flit_bits_head),
    .io_to_noc_1_flit_bits_tail(noc_tester_io_to_noc_1_flit_bits_tail),
    .io_to_noc_1_flit_bits_payload(noc_tester_io_to_noc_1_flit_bits_payload),
    .io_to_noc_1_flit_bits_egress_id(noc_tester_io_to_noc_1_flit_bits_egress_id),
    .io_to_noc_0_flit_ready(noc_tester_io_to_noc_0_flit_ready),
    .io_to_noc_0_flit_valid(noc_tester_io_to_noc_0_flit_valid),
    .io_to_noc_0_flit_bits_head(noc_tester_io_to_noc_0_flit_bits_head),
    .io_to_noc_0_flit_bits_tail(noc_tester_io_to_noc_0_flit_bits_tail),
    .io_to_noc_0_flit_bits_payload(noc_tester_io_to_noc_0_flit_bits_payload),
    .io_to_noc_0_flit_bits_egress_id(noc_tester_io_to_noc_0_flit_bits_egress_id),
    .io_from_noc_3_flit_ready(noc_tester_io_from_noc_3_flit_ready),
    .io_from_noc_3_flit_valid(noc_tester_io_from_noc_3_flit_valid),
    .io_from_noc_3_flit_bits_head(noc_tester_io_from_noc_3_flit_bits_head),
    .io_from_noc_3_flit_bits_tail(noc_tester_io_from_noc_3_flit_bits_tail),
    .io_from_noc_3_flit_bits_payload(noc_tester_io_from_noc_3_flit_bits_payload),
    .io_from_noc_3_flit_bits_ingress_id(noc_tester_io_from_noc_3_flit_bits_ingress_id),
    .io_from_noc_2_flit_ready(noc_tester_io_from_noc_2_flit_ready),
    .io_from_noc_2_flit_valid(noc_tester_io_from_noc_2_flit_valid),
    .io_from_noc_2_flit_bits_head(noc_tester_io_from_noc_2_flit_bits_head),
    .io_from_noc_2_flit_bits_tail(noc_tester_io_from_noc_2_flit_bits_tail),
    .io_from_noc_2_flit_bits_payload(noc_tester_io_from_noc_2_flit_bits_payload),
    .io_from_noc_2_flit_bits_ingress_id(noc_tester_io_from_noc_2_flit_bits_ingress_id),
    .io_from_noc_1_flit_ready(noc_tester_io_from_noc_1_flit_ready),
    .io_from_noc_1_flit_valid(noc_tester_io_from_noc_1_flit_valid),
    .io_from_noc_1_flit_bits_head(noc_tester_io_from_noc_1_flit_bits_head),
    .io_from_noc_1_flit_bits_tail(noc_tester_io_from_noc_1_flit_bits_tail),
    .io_from_noc_1_flit_bits_payload(noc_tester_io_from_noc_1_flit_bits_payload),
    .io_from_noc_1_flit_bits_ingress_id(noc_tester_io_from_noc_1_flit_bits_ingress_id),
    .io_from_noc_0_flit_ready(noc_tester_io_from_noc_0_flit_ready),
    .io_from_noc_0_flit_valid(noc_tester_io_from_noc_0_flit_valid),
    .io_from_noc_0_flit_bits_head(noc_tester_io_from_noc_0_flit_bits_head),
    .io_from_noc_0_flit_bits_tail(noc_tester_io_from_noc_0_flit_bits_tail),
    .io_from_noc_0_flit_bits_payload(noc_tester_io_from_noc_0_flit_bits_payload),
    .io_from_noc_0_flit_bits_ingress_id(noc_tester_io_from_noc_0_flit_bits_ingress_id),
    .io_success(noc_tester_io_success)
  );
  assign io_success = noc_tester_io_success; // @[TestHarness.scala 272:14]
  assign lazyNoC_clock = clock;
  assign lazyNoC_reset = reset;
  assign lazyNoC_io_ingress_3_flit_valid = noc_tester_io_to_noc_3_flit_valid; // @[TestHarness.scala 270:18]
  assign lazyNoC_io_ingress_3_flit_bits_head = noc_tester_io_to_noc_3_flit_bits_head; // @[TestHarness.scala 270:18]
  assign lazyNoC_io_ingress_3_flit_bits_tail = noc_tester_io_to_noc_3_flit_bits_tail; // @[TestHarness.scala 270:18]
  assign lazyNoC_io_ingress_3_flit_bits_payload = noc_tester_io_to_noc_3_flit_bits_payload; // @[TestHarness.scala 270:18]
  assign lazyNoC_io_ingress_3_flit_bits_egress_id = noc_tester_io_to_noc_3_flit_bits_egress_id; // @[TestHarness.scala 270:18]
  assign lazyNoC_io_ingress_2_flit_valid = noc_tester_io_to_noc_2_flit_valid; // @[TestHarness.scala 270:18]
  assign lazyNoC_io_ingress_2_flit_bits_head = noc_tester_io_to_noc_2_flit_bits_head; // @[TestHarness.scala 270:18]
  assign lazyNoC_io_ingress_2_flit_bits_tail = noc_tester_io_to_noc_2_flit_bits_tail; // @[TestHarness.scala 270:18]
  assign lazyNoC_io_ingress_2_flit_bits_payload = noc_tester_io_to_noc_2_flit_bits_payload; // @[TestHarness.scala 270:18]
  assign lazyNoC_io_ingress_2_flit_bits_egress_id = noc_tester_io_to_noc_2_flit_bits_egress_id; // @[TestHarness.scala 270:18]
  assign lazyNoC_io_ingress_1_flit_valid = noc_tester_io_to_noc_1_flit_valid; // @[TestHarness.scala 270:18]
  assign lazyNoC_io_ingress_1_flit_bits_head = noc_tester_io_to_noc_1_flit_bits_head; // @[TestHarness.scala 270:18]
  assign lazyNoC_io_ingress_1_flit_bits_tail = noc_tester_io_to_noc_1_flit_bits_tail; // @[TestHarness.scala 270:18]
  assign lazyNoC_io_ingress_1_flit_bits_payload = noc_tester_io_to_noc_1_flit_bits_payload; // @[TestHarness.scala 270:18]
  assign lazyNoC_io_ingress_1_flit_bits_egress_id = noc_tester_io_to_noc_1_flit_bits_egress_id; // @[TestHarness.scala 270:18]
  assign lazyNoC_io_ingress_0_flit_valid = noc_tester_io_to_noc_0_flit_valid; // @[TestHarness.scala 270:18]
  assign lazyNoC_io_ingress_0_flit_bits_head = noc_tester_io_to_noc_0_flit_bits_head; // @[TestHarness.scala 270:18]
  assign lazyNoC_io_ingress_0_flit_bits_tail = noc_tester_io_to_noc_0_flit_bits_tail; // @[TestHarness.scala 270:18]
  assign lazyNoC_io_ingress_0_flit_bits_payload = noc_tester_io_to_noc_0_flit_bits_payload; // @[TestHarness.scala 270:18]
  assign lazyNoC_io_ingress_0_flit_bits_egress_id = noc_tester_io_to_noc_0_flit_bits_egress_id; // @[TestHarness.scala 270:18]
  assign lazyNoC_io_router_clocks_0_clock = clock; // @[TestHarness.scala 239:40]
  assign lazyNoC_io_router_clocks_0_reset = reset; // @[TestHarness.scala 240:40]
  assign lazyNoC_io_router_clocks_1_clock = clock; // @[TestHarness.scala 239:40]
  assign lazyNoC_io_router_clocks_1_reset = reset; // @[TestHarness.scala 240:40]
  assign lazyNoC_io_router_clocks_2_clock = clock; // @[TestHarness.scala 239:40]
  assign lazyNoC_io_router_clocks_2_reset = reset; // @[TestHarness.scala 240:40]
  assign lazyNoC_io_router_clocks_3_clock = clock; // @[TestHarness.scala 239:40]
  assign lazyNoC_io_router_clocks_3_reset = reset; // @[TestHarness.scala 240:40]
  assign noc_tester_clock = clock;
  assign noc_tester_reset = reset;
  assign noc_tester_io_to_noc_3_flit_ready = lazyNoC_io_ingress_3_flit_ready; // @[TestHarness.scala 270:18]
  assign noc_tester_io_to_noc_2_flit_ready = lazyNoC_io_ingress_2_flit_ready; // @[TestHarness.scala 270:18]
  assign noc_tester_io_to_noc_1_flit_ready = lazyNoC_io_ingress_1_flit_ready; // @[TestHarness.scala 270:18]
  assign noc_tester_io_to_noc_0_flit_ready = lazyNoC_io_ingress_0_flit_ready; // @[TestHarness.scala 270:18]
  assign noc_tester_io_from_noc_3_flit_valid = lazyNoC_io_egress_3_flit_valid; // @[TestHarness.scala 271:26]
  assign noc_tester_io_from_noc_3_flit_bits_head = lazyNoC_io_egress_3_flit_bits_head; // @[TestHarness.scala 271:26]
  assign noc_tester_io_from_noc_3_flit_bits_tail = lazyNoC_io_egress_3_flit_bits_tail; // @[TestHarness.scala 271:26]
  assign noc_tester_io_from_noc_3_flit_bits_payload = lazyNoC_io_egress_3_flit_bits_payload; // @[TestHarness.scala 271:26]
  assign noc_tester_io_from_noc_3_flit_bits_ingress_id = lazyNoC_io_egress_3_flit_bits_ingress_id; // @[TestHarness.scala 271:26]
  assign noc_tester_io_from_noc_2_flit_valid = lazyNoC_io_egress_2_flit_valid; // @[TestHarness.scala 271:26]
  assign noc_tester_io_from_noc_2_flit_bits_head = lazyNoC_io_egress_2_flit_bits_head; // @[TestHarness.scala 271:26]
  assign noc_tester_io_from_noc_2_flit_bits_tail = lazyNoC_io_egress_2_flit_bits_tail; // @[TestHarness.scala 271:26]
  assign noc_tester_io_from_noc_2_flit_bits_payload = lazyNoC_io_egress_2_flit_bits_payload; // @[TestHarness.scala 271:26]
  assign noc_tester_io_from_noc_2_flit_bits_ingress_id = lazyNoC_io_egress_2_flit_bits_ingress_id; // @[TestHarness.scala 271:26]
  assign noc_tester_io_from_noc_1_flit_valid = lazyNoC_io_egress_1_flit_valid; // @[TestHarness.scala 271:26]
  assign noc_tester_io_from_noc_1_flit_bits_head = lazyNoC_io_egress_1_flit_bits_head; // @[TestHarness.scala 271:26]
  assign noc_tester_io_from_noc_1_flit_bits_tail = lazyNoC_io_egress_1_flit_bits_tail; // @[TestHarness.scala 271:26]
  assign noc_tester_io_from_noc_1_flit_bits_payload = lazyNoC_io_egress_1_flit_bits_payload; // @[TestHarness.scala 271:26]
  assign noc_tester_io_from_noc_1_flit_bits_ingress_id = lazyNoC_io_egress_1_flit_bits_ingress_id; // @[TestHarness.scala 271:26]
  assign noc_tester_io_from_noc_0_flit_valid = lazyNoC_io_egress_0_flit_valid; // @[TestHarness.scala 271:26]
  assign noc_tester_io_from_noc_0_flit_bits_head = lazyNoC_io_egress_0_flit_bits_head; // @[TestHarness.scala 271:26]
  assign noc_tester_io_from_noc_0_flit_bits_tail = lazyNoC_io_egress_0_flit_bits_tail; // @[TestHarness.scala 271:26]
  assign noc_tester_io_from_noc_0_flit_bits_payload = lazyNoC_io_egress_0_flit_bits_payload; // @[TestHarness.scala 271:26]
  assign noc_tester_io_from_noc_0_flit_bits_ingress_id = lazyNoC_io_egress_0_flit_bits_ingress_id; // @[TestHarness.scala 271:26]
endmodule
module NoCChiselTester(
  input   clock,
  input   reset
);
  wire  th_clock; // @[NocTests.scala 11:18]
  wire  th_reset; // @[NocTests.scala 11:18]
  wire  th_io_success; // @[NocTests.scala 11:18]
  TestHarness th ( // @[NocTests.scala 11:18]
    .clock(th_clock),
    .reset(th_reset),
    .io_success(th_io_success)
  );
  assign th_clock = clock;
  assign th_reset = reset;
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (th_io_success & ~reset) begin
          $finish; // @[NocTests.scala 12:30]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
