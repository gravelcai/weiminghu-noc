//

module NoC_top 
(
    input           clock,
    input           reset,

    // XP0
    output          aw_ingress_0_flit_ready,
    input           aw_ingress_0_flit_valid,
    input           aw_ingress_0_flit_bits_head,
    input           aw_ingress_0_flit_bits_tail,
    input  [81:0]   aw_ingress_0_flit_bits_payload,
    input  [1:0]    aw_ingress_0_flit_bits_egress_id,
    output          aw_egress_0_flit_valid,
    output          aw_egress_0_flit_bits_head,
    output          aw_egress_0_flit_bits_tail,
    output [81:0]   aw_egress_0_flit_bits_payload,
    output [1:0]    aw_egress_0_flit_bits_ingress_id,

    output          w_ingress_0_flit_ready,
    input           w_ingress_0_flit_valid,
    input           w_ingress_0_flit_bits_head,
    input           w_ingress_0_flit_bits_tail,
    input  [81:0]   w_ingress_0_flit_bits_payload,
    input  [1:0]    w_ingress_0_flit_bits_egress_id,
    output          w_egress_0_flit_valid,
    output          w_egress_0_flit_bits_head,
    output          w_egress_0_flit_bits_tail,
    output [81:0]   w_egress_0_flit_bits_payload,
    output [1:0]    w_egress_0_flit_bits_ingress_id,

    output          b_ingress_0_flit_ready,
    input           b_ingress_0_flit_valid,
    input           b_ingress_0_flit_bits_head,
    input           b_ingress_0_flit_bits_tail,
    input  [19:0]   b_ingress_0_flit_bits_payload,
    input  [1:0]    b_ingress_0_flit_bits_egress_id,
    output          b_egress_0_flit_valid,
    output          b_egress_0_flit_bits_head,
    output          b_egress_0_flit_bits_tail,
    output [19:0]   b_egress_0_flit_bits_payload,
    output [1:0]    b_egress_0_flit_bits_ingress_id,

    output          ar_ingress_0_flit_ready,
    input           ar_ingress_0_flit_valid,
    input           ar_ingress_0_flit_bits_head,
    input           ar_ingress_0_flit_bits_tail,
    input  [81:0]   ar_ingress_0_flit_bits_payload,
    input  [1:0]    ar_ingress_0_flit_bits_egress_id,
    output          ar_egress_0_flit_valid,
    output          ar_egress_0_flit_bits_head,
    output          ar_egress_0_flit_bits_tail,
    output [81:0]   ar_egress_0_flit_bits_payload,
    output [1:0]    ar_egress_0_flit_bits_ingress_id,

    output          r_ingress_0_flit_ready,
    input           r_ingress_0_flit_valid,
    input           r_ingress_0_flit_bits_head,
    input           r_ingress_0_flit_bits_tail,
    input  [81:0]   r_ingress_0_flit_bits_payload,
    input  [1:0]    r_ingress_0_flit_bits_egress_id,
    output          r_egress_0_flit_valid,
    output          r_egress_0_flit_bits_head,
    output          r_egress_0_flit_bits_tail,
    output [81:0]   r_egress_0_flit_bits_payload,
    output [1:0]    r_egress_0_flit_bits_ingress_id,

    // XP1
    output          aw_ingress_1_flit_ready,
    input           aw_ingress_1_flit_valid,
    input           aw_ingress_1_flit_bits_head,
    input           aw_ingress_1_flit_bits_tail,
    input  [81:0]   aw_ingress_1_flit_bits_payload,
    input  [1:0]    aw_ingress_1_flit_bits_egress_id,
    output          aw_egress_1_flit_valid,
    output          aw_egress_1_flit_bits_head,
    output          aw_egress_1_flit_bits_tail,
    output [81:0]   aw_egress_1_flit_bits_payload,
    output [1:0]    aw_egress_1_flit_bits_ingress_id,

    output          w_ingress_1_flit_ready,
    input           w_ingress_1_flit_valid,
    input           w_ingress_1_flit_bits_head,
    input           w_ingress_1_flit_bits_tail,
    input  [81:0]   w_ingress_1_flit_bits_payload,
    input  [1:0]    w_ingress_1_flit_bits_egress_id,
    output          w_egress_1_flit_valid,
    output          w_egress_1_flit_bits_head,
    output          w_egress_1_flit_bits_tail,
    output [81:0]   w_egress_1_flit_bits_payload,
    output [1:0]    w_egress_1_flit_bits_ingress_id,

    output          b_ingress_1_flit_ready,
    input           b_ingress_1_flit_valid,
    input           b_ingress_1_flit_bits_head,
    input           b_ingress_1_flit_bits_tail,
    input  [19:0]   b_ingress_1_flit_bits_payload,
    input  [1:0]    b_ingress_1_flit_bits_egress_id,
    output          b_egress_1_flit_valid,
    output          b_egress_1_flit_bits_head,
    output          b_egress_1_flit_bits_tail,
    output [19:0]   b_egress_1_flit_bits_payload,
    output [1:0]    b_egress_1_flit_bits_ingress_id,

    output          ar_ingress_1_flit_ready,
    input           ar_ingress_1_flit_valid,
    input           ar_ingress_1_flit_bits_head,
    input           ar_ingress_1_flit_bits_tail,
    input  [81:0]   ar_ingress_1_flit_bits_payload,
    input  [1:0]    ar_ingress_1_flit_bits_egress_id,
    output          ar_egress_1_flit_valid,
    output          ar_egress_1_flit_bits_head,
    output          ar_egress_1_flit_bits_tail,
    output [81:0]   ar_egress_1_flit_bits_payload,
    output [1:0]    ar_egress_1_flit_bits_ingress_id,

    output          r_ingress_1_flit_ready,
    input           r_ingress_1_flit_valid,
    input           r_ingress_1_flit_bits_head,
    input           r_ingress_1_flit_bits_tail,
    input  [81:0]   r_ingress_1_flit_bits_payload,
    input  [1:0]    r_ingress_1_flit_bits_egress_id,
    output          r_egress_1_flit_valid,
    output          r_egress_1_flit_bits_head,
    output          r_egress_1_flit_bits_tail,
    output [81:0]   r_egress_1_flit_bits_payload,
    output [1:0]    r_egress_1_flit_bits_ingress_id,

    // XP2
    output          aw_ingress_2_flit_ready,
    input           aw_ingress_2_flit_valid,
    input           aw_ingress_2_flit_bits_head,
    input           aw_ingress_2_flit_bits_tail,
    input  [81:0]   aw_ingress_2_flit_bits_payload,
    input  [1:0]    aw_ingress_2_flit_bits_egress_id,
    output          aw_egress_2_flit_valid,
    output          aw_egress_2_flit_bits_head,
    output          aw_egress_2_flit_bits_tail,
    output [81:0]   aw_egress_2_flit_bits_payload,
    output [1:0]    aw_egress_2_flit_bits_ingress_id,

    output          w_ingress_2_flit_ready,
    input           w_ingress_2_flit_valid,
    input           w_ingress_2_flit_bits_head,
    input           w_ingress_2_flit_bits_tail,
    input  [81:0]   w_ingress_2_flit_bits_payload,
    input  [1:0]    w_ingress_2_flit_bits_egress_id,
    output          w_egress_2_flit_valid,
    output          w_egress_2_flit_bits_head,
    output          w_egress_2_flit_bits_tail,
    output [81:0]   w_egress_2_flit_bits_payload,
    output [1:0]    w_egress_2_flit_bits_ingress_id,

    output          b_ingress_2_flit_ready,
    input           b_ingress_2_flit_valid,
    input           b_ingress_2_flit_bits_head,
    input           b_ingress_2_flit_bits_tail,
    input  [19:0]   b_ingress_2_flit_bits_payload,
    input  [1:0]    b_ingress_2_flit_bits_egress_id,
    output          b_egress_2_flit_valid,
    output          b_egress_2_flit_bits_head,
    output          b_egress_2_flit_bits_tail,
    output [19:0]   b_egress_2_flit_bits_payload,
    output [1:0]    b_egress_2_flit_bits_ingress_id,

    output          ar_ingress_2_flit_ready,
    input           ar_ingress_2_flit_valid,
    input           ar_ingress_2_flit_bits_head,
    input           ar_ingress_2_flit_bits_tail,
    input  [81:0]   ar_ingress_2_flit_bits_payload,
    input  [1:0]    ar_ingress_2_flit_bits_egress_id,
    output          ar_egress_2_flit_valid,
    output          ar_egress_2_flit_bits_head,
    output          ar_egress_2_flit_bits_tail,
    output [81:0]   ar_egress_2_flit_bits_payload,
    output [1:0]    ar_egress_2_flit_bits_ingress_id,

    output          r_ingress_2_flit_ready,
    input           r_ingress_2_flit_valid,
    input           r_ingress_2_flit_bits_head,
    input           r_ingress_2_flit_bits_tail,
    input  [81:0]   r_ingress_2_flit_bits_payload,
    input  [1:0]    r_ingress_2_flit_bits_egress_id,
    output          r_egress_2_flit_valid,
    output          r_egress_2_flit_bits_head,
    output          r_egress_2_flit_bits_tail,
    output [81:0]   r_egress_2_flit_bits_payload,
    output [1:0]    r_egress_2_flit_bits_ingress_id,

    // XP3
    output          aw_ingress_3_flit_ready,
    input           aw_ingress_3_flit_valid,
    input           aw_ingress_3_flit_bits_head,
    input           aw_ingress_3_flit_bits_tail,
    input  [81:0]   aw_ingress_3_flit_bits_payload,
    input  [1:0]    aw_ingress_3_flit_bits_egress_id,
    output          aw_egress_3_flit_valid,
    output          aw_egress_3_flit_bits_head,
    output          aw_egress_3_flit_bits_tail,
    output [81:0]   aw_egress_3_flit_bits_payload,
    output [1:0]    aw_egress_3_flit_bits_ingress_id,

    output          w_ingress_3_flit_ready,
    input           w_ingress_3_flit_valid,
    input           w_ingress_3_flit_bits_head,
    input           w_ingress_3_flit_bits_tail,
    input  [81:0]   w_ingress_3_flit_bits_payload,
    input  [1:0]    w_ingress_3_flit_bits_egress_id,
    output          w_egress_3_flit_valid,
    output          w_egress_3_flit_bits_head,
    output          w_egress_3_flit_bits_tail,
    output [81:0]   w_egress_3_flit_bits_payload,
    output [1:0]    w_egress_3_flit_bits_ingress_id,

    output          b_ingress_3_flit_ready,
    input           b_ingress_3_flit_valid,
    input           b_ingress_3_flit_bits_head,
    input           b_ingress_3_flit_bits_tail,
    input  [19:0]   b_ingress_3_flit_bits_payload,
    input  [1:0]    b_ingress_3_flit_bits_egress_id,
    output          b_egress_3_flit_valid,
    output          b_egress_3_flit_bits_head,
    output          b_egress_3_flit_bits_tail,
    output [19:0]   b_egress_3_flit_bits_payload,
    output [1:0]    b_egress_3_flit_bits_ingress_id,

    output          ar_ingress_3_flit_ready,
    input           ar_ingress_3_flit_valid,
    input           ar_ingress_3_flit_bits_head,
    input           ar_ingress_3_flit_bits_tail,
    input  [81:0]   ar_ingress_3_flit_bits_payload,
    input  [1:0]    ar_ingress_3_flit_bits_egress_id,
    output          ar_egress_3_flit_valid,
    output          ar_egress_3_flit_bits_head,
    output          ar_egress_3_flit_bits_tail,
    output [81:0]   ar_egress_3_flit_bits_payload,
    output [1:0]    ar_egress_3_flit_bits_ingress_id,

    output          r_ingress_3_flit_ready,
    input           r_ingress_3_flit_valid,
    input           r_ingress_3_flit_bits_head,
    input           r_ingress_3_flit_bits_tail,
    input  [81:0]   r_ingress_3_flit_bits_payload,
    input  [1:0]    r_ingress_3_flit_bits_egress_id,
    output          r_egress_3_flit_valid,
    output          r_egress_3_flit_bits_head,
    output          r_egress_3_flit_bits_tail,
    output [81:0]   r_egress_3_flit_bits_payload,
    output [1:0]    r_egress_3_flit_bits_ingress_id

);

//---------------------------------------------------------------------
// NoC instantiate.
//---------------------------------------------------------------------

    // AW
    NoC_82b u_aw_channel (
        .clock                                  ( clock ),
        .reset                                  ( reset ),
        .io_ingress_3_flit_ready                ( aw_ingress_3_flit_ready ),
        .io_ingress_3_flit_valid                ( aw_ingress_3_flit_valid ),
        .io_ingress_3_flit_bits_head            ( aw_ingress_3_flit_bits_head ),
        .io_ingress_3_flit_bits_tail            ( aw_ingress_3_flit_bits_tail ),
        .io_ingress_3_flit_bits_payload         ( aw_ingress_3_flit_bits_payload ),
        .io_ingress_3_flit_bits_egress_id       ( aw_ingress_3_flit_bits_egress_id ),
        .io_ingress_2_flit_ready                ( aw_ingress_2_flit_ready ),
        .io_ingress_2_flit_valid                ( aw_ingress_2_flit_valid ),
        .io_ingress_2_flit_bits_head            ( aw_ingress_2_flit_bits_head ),
        .io_ingress_2_flit_bits_tail            ( aw_ingress_2_flit_bits_tail ),
        .io_ingress_2_flit_bits_payload         ( aw_ingress_2_flit_bits_payload ),
        .io_ingress_2_flit_bits_egress_id       ( aw_ingress_2_flit_bits_egress_id ),
        .io_ingress_1_flit_ready                ( aw_ingress_1_flit_ready ),
        .io_ingress_1_flit_valid                ( aw_ingress_1_flit_valid ),
        .io_ingress_1_flit_bits_head            ( aw_ingress_1_flit_bits_head ),
        .io_ingress_1_flit_bits_tail            ( aw_ingress_1_flit_bits_tail ),
        .io_ingress_1_flit_bits_payload         ( aw_ingress_1_flit_bits_payload ),
        .io_ingress_1_flit_bits_egress_id       ( aw_ingress_1_flit_bits_egress_id ),
        .io_ingress_0_flit_ready                ( aw_ingress_0_flit_ready ),
        .io_ingress_0_flit_valid                ( aw_ingress_0_flit_valid ),
        .io_ingress_0_flit_bits_head            ( aw_ingress_0_flit_bits_head ),
        .io_ingress_0_flit_bits_tail            ( aw_ingress_0_flit_bits_tail ),
        .io_ingress_0_flit_bits_payload         ( aw_ingress_0_flit_bits_payload ),
        .io_ingress_0_flit_bits_egress_id       ( aw_ingress_0_flit_bits_egress_id ),
        .io_egress_3_flit_valid                 ( aw_egress_3_flit_valid ),
        .io_egress_3_flit_bits_head             ( aw_egress_3_flit_bits_head ),
        .io_egress_3_flit_bits_tail             ( aw_egress_3_flit_bits_tail ),
        .io_egress_3_flit_bits_payload          ( aw_egress_3_flit_bits_payload ),
        .io_egress_3_flit_bits_ingress_id       ( aw_egress_3_flit_bits_ingress_id ),
        .io_egress_2_flit_valid                 ( aw_egress_2_flit_valid ),
        .io_egress_2_flit_bits_head             ( aw_egress_2_flit_bits_head ),
        .io_egress_2_flit_bits_tail             ( aw_egress_2_flit_bits_tail ),
        .io_egress_2_flit_bits_payload          ( aw_egress_2_flit_bits_payload ),
        .io_egress_2_flit_bits_ingress_id       ( aw_egress_2_flit_bits_ingress_id ),
        .io_egress_1_flit_valid                 ( aw_egress_1_flit_valid ),
        .io_egress_1_flit_bits_head             ( aw_egress_1_flit_bits_head ),
        .io_egress_1_flit_bits_tail             ( aw_egress_1_flit_bits_tail ),
        .io_egress_1_flit_bits_payload          ( aw_egress_1_flit_bits_payload ),
        .io_egress_1_flit_bits_ingress_id       ( aw_egress_1_flit_bits_ingress_id ),
        .io_egress_0_flit_valid                 ( aw_egress_0_flit_valid ),
        .io_egress_0_flit_bits_head             ( aw_egress_0_flit_bits_head ),
        .io_egress_0_flit_bits_tail             ( aw_egress_0_flit_bits_tail ),
        .io_egress_0_flit_bits_payload          ( aw_egress_0_flit_bits_payload ),
        .io_egress_0_flit_bits_ingress_id       ( aw_egress_0_flit_bits_ingress_id ),
        .io_router_clocks_0_clock               ( clock ),
        .io_router_clocks_0_reset               ( reset ),
        .io_router_clocks_1_clock               ( clock ),
        .io_router_clocks_1_reset               ( reset ),
        .io_router_clocks_2_clock               ( clock ),
        .io_router_clocks_2_reset               ( reset ),
        .io_router_clocks_3_clock               ( clock ),
        .io_router_clocks_3_reset               ( reset )
    );

    // W
    NoC_82b u_w_channel (
        .clock                                  ( clock ),
        .reset                                  ( reset ),
        .io_ingress_3_flit_ready                ( w_ingress_3_flit_ready ),
        .io_ingress_3_flit_valid                ( w_ingress_3_flit_valid ),
        .io_ingress_3_flit_bits_head            ( w_ingress_3_flit_bits_head ),
        .io_ingress_3_flit_bits_tail            ( w_ingress_3_flit_bits_tail ),
        .io_ingress_3_flit_bits_payload         ( w_ingress_3_flit_bits_payload ),
        .io_ingress_3_flit_bits_egress_id       ( w_ingress_3_flit_bits_egress_id ),
        .io_ingress_2_flit_ready                ( w_ingress_2_flit_ready ),
        .io_ingress_2_flit_valid                ( w_ingress_2_flit_valid ),
        .io_ingress_2_flit_bits_head            ( w_ingress_2_flit_bits_head ),
        .io_ingress_2_flit_bits_tail            ( w_ingress_2_flit_bits_tail ),
        .io_ingress_2_flit_bits_payload         ( w_ingress_2_flit_bits_payload ),
        .io_ingress_2_flit_bits_egress_id       ( w_ingress_2_flit_bits_egress_id ),
        .io_ingress_1_flit_ready                ( w_ingress_1_flit_ready ),
        .io_ingress_1_flit_valid                ( w_ingress_1_flit_valid ),
        .io_ingress_1_flit_bits_head            ( w_ingress_1_flit_bits_head ),
        .io_ingress_1_flit_bits_tail            ( w_ingress_1_flit_bits_tail ),
        .io_ingress_1_flit_bits_payload         ( w_ingress_1_flit_bits_payload ),
        .io_ingress_1_flit_bits_egress_id       ( w_ingress_1_flit_bits_egress_id ),
        .io_ingress_0_flit_ready                ( w_ingress_0_flit_ready ),
        .io_ingress_0_flit_valid                ( w_ingress_0_flit_valid ),
        .io_ingress_0_flit_bits_head            ( w_ingress_0_flit_bits_head ),
        .io_ingress_0_flit_bits_tail            ( w_ingress_0_flit_bits_tail ),
        .io_ingress_0_flit_bits_payload         ( w_ingress_0_flit_bits_payload ),
        .io_ingress_0_flit_bits_egress_id       ( w_ingress_0_flit_bits_egress_id ),
        .io_egress_3_flit_valid                 ( w_egress_3_flit_valid ),
        .io_egress_3_flit_bits_head             ( w_egress_3_flit_bits_head ),
        .io_egress_3_flit_bits_tail             ( w_egress_3_flit_bits_tail ),
        .io_egress_3_flit_bits_payload          ( w_egress_3_flit_bits_payload ),
        .io_egress_3_flit_bits_ingress_id       ( w_egress_3_flit_bits_ingress_id ),
        .io_egress_2_flit_valid                 ( w_egress_2_flit_valid ),
        .io_egress_2_flit_bits_head             ( w_egress_2_flit_bits_head ),
        .io_egress_2_flit_bits_tail             ( w_egress_2_flit_bits_tail ),
        .io_egress_2_flit_bits_payload          ( w_egress_2_flit_bits_payload ),
        .io_egress_2_flit_bits_ingress_id       ( w_egress_2_flit_bits_ingress_id ),
        .io_egress_1_flit_valid                 ( w_egress_1_flit_valid ),
        .io_egress_1_flit_bits_head             ( w_egress_1_flit_bits_head ),
        .io_egress_1_flit_bits_tail             ( w_egress_1_flit_bits_tail ),
        .io_egress_1_flit_bits_payload          ( w_egress_1_flit_bits_payload ),
        .io_egress_1_flit_bits_ingress_id       ( w_egress_1_flit_bits_ingress_id ),
        .io_egress_0_flit_valid                 ( w_egress_0_flit_valid ),
        .io_egress_0_flit_bits_head             ( w_egress_0_flit_bits_head ),
        .io_egress_0_flit_bits_tail             ( w_egress_0_flit_bits_tail ),
        .io_egress_0_flit_bits_payload          ( w_egress_0_flit_bits_payload ),
        .io_egress_0_flit_bits_ingress_id       ( w_egress_0_flit_bits_ingress_id ),
        .io_router_clocks_0_clock               ( clock ),
        .io_router_clocks_0_reset               ( reset ),
        .io_router_clocks_1_clock               ( clock ),
        .io_router_clocks_1_reset               ( reset ),
        .io_router_clocks_2_clock               ( clock ),
        .io_router_clocks_2_reset               ( reset ),
        .io_router_clocks_3_clock               ( clock ),
        .io_router_clocks_3_reset               ( reset )
    );


    // B
    NoC_82b u_b_channel (
        .clock                                  ( clock ),
        .reset                                  ( reset ),
        .io_ingress_3_flit_ready                ( b_ingress_3_flit_ready ),
        .io_ingress_3_flit_valid                ( b_ingress_3_flit_valid ),
        .io_ingress_3_flit_bits_head            ( b_ingress_3_flit_bits_head ),
        .io_ingress_3_flit_bits_tail            ( b_ingress_3_flit_bits_tail ),
        .io_ingress_3_flit_bits_payload         ( b_ingress_3_flit_bits_payload ),
        .io_ingress_3_flit_bits_egress_id       ( b_ingress_3_flit_bits_egress_id ),
        .io_ingress_2_flit_ready                ( b_ingress_2_flit_ready ),
        .io_ingress_2_flit_valid                ( b_ingress_2_flit_valid ),
        .io_ingress_2_flit_bits_head            ( b_ingress_2_flit_bits_head ),
        .io_ingress_2_flit_bits_tail            ( b_ingress_2_flit_bits_tail ),
        .io_ingress_2_flit_bits_payload         ( b_ingress_2_flit_bits_payload ),
        .io_ingress_2_flit_bits_egress_id       ( b_ingress_2_flit_bits_egress_id ),
        .io_ingress_1_flit_ready                ( b_ingress_1_flit_ready ),
        .io_ingress_1_flit_valid                ( b_ingress_1_flit_valid ),
        .io_ingress_1_flit_bits_head            ( b_ingress_1_flit_bits_head ),
        .io_ingress_1_flit_bits_tail            ( b_ingress_1_flit_bits_tail ),
        .io_ingress_1_flit_bits_payload         ( b_ingress_1_flit_bits_payload ),
        .io_ingress_1_flit_bits_egress_id       ( b_ingress_1_flit_bits_egress_id ),
        .io_ingress_0_flit_ready                ( b_ingress_0_flit_ready ),
        .io_ingress_0_flit_valid                ( b_ingress_0_flit_valid ),
        .io_ingress_0_flit_bits_head            ( b_ingress_0_flit_bits_head ),
        .io_ingress_0_flit_bits_tail            ( b_ingress_0_flit_bits_tail ),
        .io_ingress_0_flit_bits_payload         ( b_ingress_0_flit_bits_payload ),
        .io_ingress_0_flit_bits_egress_id       ( b_ingress_0_flit_bits_egress_id ),
        .io_egress_3_flit_valid                 ( b_egress_3_flit_valid ),
        .io_egress_3_flit_bits_head             ( b_egress_3_flit_bits_head ),
        .io_egress_3_flit_bits_tail             ( b_egress_3_flit_bits_tail ),
        .io_egress_3_flit_bits_payload          ( b_egress_3_flit_bits_payload ),
        .io_egress_3_flit_bits_ingress_id       ( b_egress_3_flit_bits_ingress_id ),
        .io_egress_2_flit_valid                 ( b_egress_2_flit_valid ),
        .io_egress_2_flit_bits_head             ( b_egress_2_flit_bits_head ),
        .io_egress_2_flit_bits_tail             ( b_egress_2_flit_bits_tail ),
        .io_egress_2_flit_bits_payload          ( b_egress_2_flit_bits_payload ),
        .io_egress_2_flit_bits_ingress_id       ( b_egress_2_flit_bits_ingress_id ),
        .io_egress_1_flit_valid                 ( b_egress_1_flit_valid ),
        .io_egress_1_flit_bits_head             ( b_egress_1_flit_bits_head ),
        .io_egress_1_flit_bits_tail             ( b_egress_1_flit_bits_tail ),
        .io_egress_1_flit_bits_payload          ( b_egress_1_flit_bits_payload ),
        .io_egress_1_flit_bits_ingress_id       ( b_egress_1_flit_bits_ingress_id ),
        .io_egress_0_flit_valid                 ( b_egress_0_flit_valid ),
        .io_egress_0_flit_bits_head             ( b_egress_0_flit_bits_head ),
        .io_egress_0_flit_bits_tail             ( b_egress_0_flit_bits_tail ),
        .io_egress_0_flit_bits_payload          ( b_egress_0_flit_bits_payload ),
        .io_egress_0_flit_bits_ingress_id       ( b_egress_0_flit_bits_ingress_id ),
        .io_router_clocks_0_clock               ( clock ),
        .io_router_clocks_0_reset               ( reset ),
        .io_router_clocks_1_clock               ( clock ),
        .io_router_clocks_1_reset               ( reset ),
        .io_router_clocks_2_clock               ( clock ),
        .io_router_clocks_2_reset               ( reset ),
        .io_router_clocks_3_clock               ( clock ),
        .io_router_clocks_3_reset               ( reset )
    );

    // AR
    NoC_82b u_ar_channel (
        .clock                                  ( clock ),
        .reset                                  ( reset ),
        .io_ingress_3_flit_ready                ( ar_ingress_3_flit_ready ),
        .io_ingress_3_flit_valid                ( ar_ingress_3_flit_valid ),
        .io_ingress_3_flit_bits_head            ( ar_ingress_3_flit_bits_head ),
        .io_ingress_3_flit_bits_tail            ( ar_ingress_3_flit_bits_tail ),
        .io_ingress_3_flit_bits_payload         ( ar_ingress_3_flit_bits_payload ),
        .io_ingress_3_flit_bits_egress_id       ( ar_ingress_3_flit_bits_egress_id ),
        .io_ingress_2_flit_ready                ( ar_ingress_2_flit_ready ),
        .io_ingress_2_flit_valid                ( ar_ingress_2_flit_valid ),
        .io_ingress_2_flit_bits_head            ( ar_ingress_2_flit_bits_head ),
        .io_ingress_2_flit_bits_tail            ( ar_ingress_2_flit_bits_tail ),
        .io_ingress_2_flit_bits_payload         ( ar_ingress_2_flit_bits_payload ),
        .io_ingress_2_flit_bits_egress_id       ( ar_ingress_2_flit_bits_egress_id ),
        .io_ingress_1_flit_ready                ( ar_ingress_1_flit_ready ),
        .io_ingress_1_flit_valid                ( ar_ingress_1_flit_valid ),
        .io_ingress_1_flit_bits_head            ( ar_ingress_1_flit_bits_head ),
        .io_ingress_1_flit_bits_tail            ( ar_ingress_1_flit_bits_tail ),
        .io_ingress_1_flit_bits_payload         ( ar_ingress_1_flit_bits_payload ),
        .io_ingress_1_flit_bits_egress_id       ( ar_ingress_1_flit_bits_egress_id ),
        .io_ingress_0_flit_ready                ( ar_ingress_0_flit_ready ),
        .io_ingress_0_flit_valid                ( ar_ingress_0_flit_valid ),
        .io_ingress_0_flit_bits_head            ( ar_ingress_0_flit_bits_head ),
        .io_ingress_0_flit_bits_tail            ( ar_ingress_0_flit_bits_tail ),
        .io_ingress_0_flit_bits_payload         ( ar_ingress_0_flit_bits_payload ),
        .io_ingress_0_flit_bits_egress_id       ( ar_ingress_0_flit_bits_egress_id ),
        .io_egress_3_flit_valid                 ( ar_egress_3_flit_valid ),
        .io_egress_3_flit_bits_head             ( ar_egress_3_flit_bits_head ),
        .io_egress_3_flit_bits_tail             ( ar_egress_3_flit_bits_tail ),
        .io_egress_3_flit_bits_payload          ( ar_egress_3_flit_bits_payload ),
        .io_egress_3_flit_bits_ingress_id       ( ar_egress_3_flit_bits_ingress_id ),
        .io_egress_2_flit_valid                 ( ar_egress_2_flit_valid ),
        .io_egress_2_flit_bits_head             ( ar_egress_2_flit_bits_head ),
        .io_egress_2_flit_bits_tail             ( ar_egress_2_flit_bits_tail ),
        .io_egress_2_flit_bits_payload          ( ar_egress_2_flit_bits_payload ),
        .io_egress_2_flit_bits_ingress_id       ( ar_egress_2_flit_bits_ingress_id ),
        .io_egress_1_flit_valid                 ( ar_egress_1_flit_valid ),
        .io_egress_1_flit_bits_head             ( ar_egress_1_flit_bits_head ),
        .io_egress_1_flit_bits_tail             ( ar_egress_1_flit_bits_tail ),
        .io_egress_1_flit_bits_payload          ( ar_egress_1_flit_bits_payload ),
        .io_egress_1_flit_bits_ingress_id       ( ar_egress_1_flit_bits_ingress_id ),
        .io_egress_0_flit_valid                 ( ar_egress_0_flit_valid ),
        .io_egress_0_flit_bits_head             ( ar_egress_0_flit_bits_head ),
        .io_egress_0_flit_bits_tail             ( ar_egress_0_flit_bits_tail ),
        .io_egress_0_flit_bits_payload          ( ar_egress_0_flit_bits_payload ),
        .io_egress_0_flit_bits_ingress_id       ( ar_egress_0_flit_bits_ingress_id ),
        .io_router_clocks_0_clock               ( clock ),
        .io_router_clocks_0_reset               ( reset ),
        .io_router_clocks_1_clock               ( clock ),
        .io_router_clocks_1_reset               ( reset ),
        .io_router_clocks_2_clock               ( clock ),
        .io_router_clocks_2_reset               ( reset ),
        .io_router_clocks_3_clock               ( clock ),
        .io_router_clocks_3_reset               ( reset )
    );


    // R
    NoC_82b u_r_channel (
        .clock                                  ( clock ),
        .reset                                  ( reset ),
        .io_ingress_3_flit_ready                ( r_ingress_3_flit_ready ),
        .io_ingress_3_flit_valid                ( r_ingress_3_flit_valid ),
        .io_ingress_3_flit_bits_head            ( r_ingress_3_flit_bits_head ),
        .io_ingress_3_flit_bits_tail            ( r_ingress_3_flit_bits_tail ),
        .io_ingress_3_flit_bits_payload         ( r_ingress_3_flit_bits_payload ),
        .io_ingress_3_flit_bits_egress_id       ( r_ingress_3_flit_bits_egress_id ),
        .io_ingress_2_flit_ready                ( r_ingress_2_flit_ready ),
        .io_ingress_2_flit_valid                ( r_ingress_2_flit_valid ),
        .io_ingress_2_flit_bits_head            ( r_ingress_2_flit_bits_head ),
        .io_ingress_2_flit_bits_tail            ( r_ingress_2_flit_bits_tail ),
        .io_ingress_2_flit_bits_payload         ( r_ingress_2_flit_bits_payload ),
        .io_ingress_2_flit_bits_egress_id       ( r_ingress_2_flit_bits_egress_id ),
        .io_ingress_1_flit_ready                ( r_ingress_1_flit_ready ),
        .io_ingress_1_flit_valid                ( r_ingress_1_flit_valid ),
        .io_ingress_1_flit_bits_head            ( r_ingress_1_flit_bits_head ),
        .io_ingress_1_flit_bits_tail            ( r_ingress_1_flit_bits_tail ),
        .io_ingress_1_flit_bits_payload         ( r_ingress_1_flit_bits_payload ),
        .io_ingress_1_flit_bits_egress_id       ( r_ingress_1_flit_bits_egress_id ),
        .io_ingress_0_flit_ready                ( r_ingress_0_flit_ready ),
        .io_ingress_0_flit_valid                ( r_ingress_0_flit_valid ),
        .io_ingress_0_flit_bits_head            ( r_ingress_0_flit_bits_head ),
        .io_ingress_0_flit_bits_tail            ( r_ingress_0_flit_bits_tail ),
        .io_ingress_0_flit_bits_payload         ( r_ingress_0_flit_bits_payload ),
        .io_ingress_0_flit_bits_egress_id       ( r_ingress_0_flit_bits_egress_id ),
        .io_egress_3_flit_valid                 ( r_egress_3_flit_valid ),
        .io_egress_3_flit_bits_head             ( r_egress_3_flit_bits_head ),
        .io_egress_3_flit_bits_tail             ( r_egress_3_flit_bits_tail ),
        .io_egress_3_flit_bits_payload          ( r_egress_3_flit_bits_payload ),
        .io_egress_3_flit_bits_ingress_id       ( r_egress_3_flit_bits_ingress_id ),
        .io_egress_2_flit_valid                 ( r_egress_2_flit_valid ),
        .io_egress_2_flit_bits_head             ( r_egress_2_flit_bits_head ),
        .io_egress_2_flit_bits_tail             ( r_egress_2_flit_bits_tail ),
        .io_egress_2_flit_bits_payload          ( r_egress_2_flit_bits_payload ),
        .io_egress_2_flit_bits_ingress_id       ( r_egress_2_flit_bits_ingress_id ),
        .io_egress_1_flit_valid                 ( r_egress_1_flit_valid ),
        .io_egress_1_flit_bits_head             ( r_egress_1_flit_bits_head ),
        .io_egress_1_flit_bits_tail             ( r_egress_1_flit_bits_tail ),
        .io_egress_1_flit_bits_payload          ( r_egress_1_flit_bits_payload ),
        .io_egress_1_flit_bits_ingress_id       ( r_egress_1_flit_bits_ingress_id ),
        .io_egress_0_flit_valid                 ( r_egress_0_flit_valid ),
        .io_egress_0_flit_bits_head             ( r_egress_0_flit_bits_head ),
        .io_egress_0_flit_bits_tail             ( r_egress_0_flit_bits_tail ),
        .io_egress_0_flit_bits_payload          ( r_egress_0_flit_bits_payload ),
        .io_egress_0_flit_bits_ingress_id       ( r_egress_0_flit_bits_ingress_id ),
        .io_router_clocks_0_clock               ( clock ),
        .io_router_clocks_0_reset               ( reset ),
        .io_router_clocks_1_clock               ( clock ),
        .io_router_clocks_1_reset               ( reset ),
        .io_router_clocks_2_clock               ( clock ),
        .io_router_clocks_2_reset               ( reset ),
        .io_router_clocks_3_clock               ( clock ),
        .io_router_clocks_3_reset               ( reset )
    );



endmodule
