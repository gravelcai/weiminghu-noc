module tb_SoC;





endmodule