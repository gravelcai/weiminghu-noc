module Queue(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_head,
  input         io_enq_bits_tail,
  input  [63:0] io_enq_bits_payload,
  input  [1:0]  io_enq_bits_flow_ingress_node,
  input  [1:0]  io_enq_bits_flow_egress_node,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_head,
  output        io_deq_bits_tail,
  output [63:0] io_deq_bits_payload,
  output [1:0]  io_deq_bits_flow_ingress_node,
  output [1:0]  io_deq_bits_flow_egress_node
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg  ram_head [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_head_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_head_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_head_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_tail [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_tail_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_tail_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_tail_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_en; // @[Decoupled.scala 273:95]
  reg [63:0] ram_payload [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_payload_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_payload_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [63:0] ram_payload_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [63:0] ram_payload_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_payload_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_payload_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_payload_MPORT_en; // @[Decoupled.scala 273:95]
  reg [1:0] ram_flow_ingress_node [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_flow_ingress_node_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_flow_ingress_node_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [1:0] ram_flow_ingress_node_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_flow_ingress_node_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_flow_ingress_node_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_flow_ingress_node_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_flow_ingress_node_MPORT_en; // @[Decoupled.scala 273:95]
  reg [1:0] ram_flow_egress_node [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_flow_egress_node_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_flow_egress_node_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [1:0] ram_flow_egress_node_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_flow_egress_node_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_flow_egress_node_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_flow_egress_node_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_flow_egress_node_MPORT_en; // @[Decoupled.scala 273:95]
  reg  enq_ptr_value; // @[Counter.scala 61:40]
  reg  deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  assign ram_head_io_deq_bits_MPORT_en = 1'h1;
  assign ram_head_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_head_io_deq_bits_MPORT_data = ram_head[ram_head_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_head_MPORT_data = io_enq_bits_head;
  assign ram_head_MPORT_addr = enq_ptr_value;
  assign ram_head_MPORT_mask = 1'h1;
  assign ram_head_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tail_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tail_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_tail_io_deq_bits_MPORT_data = ram_tail[ram_tail_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_tail_MPORT_data = io_enq_bits_tail;
  assign ram_tail_MPORT_addr = enq_ptr_value;
  assign ram_tail_MPORT_mask = 1'h1;
  assign ram_tail_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_payload_io_deq_bits_MPORT_en = 1'h1;
  assign ram_payload_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_payload_io_deq_bits_MPORT_data = ram_payload[ram_payload_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_payload_MPORT_data = io_enq_bits_payload;
  assign ram_payload_MPORT_addr = enq_ptr_value;
  assign ram_payload_MPORT_mask = 1'h1;
  assign ram_payload_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_flow_ingress_node_io_deq_bits_MPORT_en = 1'h1;
  assign ram_flow_ingress_node_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_flow_ingress_node_io_deq_bits_MPORT_data =
    ram_flow_ingress_node[ram_flow_ingress_node_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_flow_ingress_node_MPORT_data = io_enq_bits_flow_ingress_node;
  assign ram_flow_ingress_node_MPORT_addr = enq_ptr_value;
  assign ram_flow_ingress_node_MPORT_mask = 1'h1;
  assign ram_flow_ingress_node_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_flow_egress_node_io_deq_bits_MPORT_en = 1'h1;
  assign ram_flow_egress_node_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_flow_egress_node_io_deq_bits_MPORT_data = ram_flow_egress_node[ram_flow_egress_node_io_deq_bits_MPORT_addr]
    ; // @[Decoupled.scala 273:95]
  assign ram_flow_egress_node_MPORT_data = io_enq_bits_flow_egress_node;
  assign ram_flow_egress_node_MPORT_addr = enq_ptr_value;
  assign ram_flow_egress_node_MPORT_mask = 1'h1;
  assign ram_flow_egress_node_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_head = ram_head_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_tail = ram_tail_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_payload = ram_payload_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_flow_ingress_node = ram_flow_ingress_node_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_flow_egress_node = ram_flow_egress_node_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  always @(posedge clock) begin
    if (ram_head_MPORT_en & ram_head_MPORT_mask) begin
      ram_head[ram_head_MPORT_addr] <= ram_head_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_tail_MPORT_en & ram_tail_MPORT_mask) begin
      ram_tail[ram_tail_MPORT_addr] <= ram_tail_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_payload_MPORT_en & ram_payload_MPORT_mask) begin
      ram_payload[ram_payload_MPORT_addr] <= ram_payload_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_flow_ingress_node_MPORT_en & ram_flow_ingress_node_MPORT_mask) begin
      ram_flow_ingress_node[ram_flow_ingress_node_MPORT_addr] <= ram_flow_ingress_node_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_flow_egress_node_MPORT_en & ram_flow_egress_node_MPORT_mask) begin
      ram_flow_egress_node[ram_flow_egress_node_MPORT_addr] <= ram_flow_egress_node_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_head[initvar] = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_tail[initvar] = _RAND_1[0:0];
  _RAND_2 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload[initvar] = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_flow_ingress_node[initvar] = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_flow_egress_node[initvar] = _RAND_4[1:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  enq_ptr_value = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  deq_ptr_value = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  maybe_full = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_1(
  input   clock,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input   io_enq_bits_vc_sel_1_0,
  input   io_enq_bits_vc_sel_1_1,
  input   io_enq_bits_vc_sel_1_2,
  input   io_enq_bits_vc_sel_1_3,
  input   io_enq_bits_vc_sel_0_0,
  input   io_enq_bits_vc_sel_0_1,
  input   io_enq_bits_vc_sel_0_2,
  input   io_enq_bits_vc_sel_0_3,
  input   io_deq_ready,
  output  io_deq_valid,
  output  io_deq_bits_vc_sel_1_0,
  output  io_deq_bits_vc_sel_1_1,
  output  io_deq_bits_vc_sel_1_2,
  output  io_deq_bits_vc_sel_1_3,
  output  io_deq_bits_vc_sel_0_0,
  output  io_deq_bits_vc_sel_0_1,
  output  io_deq_bits_vc_sel_0_2,
  output  io_deq_bits_vc_sel_0_3
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg  ram_vc_sel_1_0 [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_0_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_0_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_0_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_0_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_0_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_0_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_vc_sel_1_1 [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_1_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_1_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_1_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_1_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_1_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_1_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_vc_sel_1_2 [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_2_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_2_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_2_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_2_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_2_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_2_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_vc_sel_1_3 [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_3_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_3_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_3_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_3_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_3_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_3_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_vc_sel_0_0 [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_0_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_0_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_0_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_0_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_0_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_0_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_vc_sel_0_1 [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_1_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_1_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_1_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_1_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_1_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_1_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_vc_sel_0_2 [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_2_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_2_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_2_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_2_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_2_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_2_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_vc_sel_0_3 [0:1]; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_3_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_3_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_3_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_3_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_3_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_3_MPORT_en; // @[Decoupled.scala 273:95]
  reg  enq_ptr_value; // @[Counter.scala 61:40]
  reg  deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  assign ram_vc_sel_1_0_io_deq_bits_MPORT_en = 1'h1;
  assign ram_vc_sel_1_0_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_vc_sel_1_0_io_deq_bits_MPORT_data = ram_vc_sel_1_0[ram_vc_sel_1_0_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_vc_sel_1_0_MPORT_data = io_enq_bits_vc_sel_1_0;
  assign ram_vc_sel_1_0_MPORT_addr = enq_ptr_value;
  assign ram_vc_sel_1_0_MPORT_mask = 1'h1;
  assign ram_vc_sel_1_0_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_vc_sel_1_1_io_deq_bits_MPORT_en = 1'h1;
  assign ram_vc_sel_1_1_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_vc_sel_1_1_io_deq_bits_MPORT_data = ram_vc_sel_1_1[ram_vc_sel_1_1_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_vc_sel_1_1_MPORT_data = io_enq_bits_vc_sel_1_1;
  assign ram_vc_sel_1_1_MPORT_addr = enq_ptr_value;
  assign ram_vc_sel_1_1_MPORT_mask = 1'h1;
  assign ram_vc_sel_1_1_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_vc_sel_1_2_io_deq_bits_MPORT_en = 1'h1;
  assign ram_vc_sel_1_2_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_vc_sel_1_2_io_deq_bits_MPORT_data = ram_vc_sel_1_2[ram_vc_sel_1_2_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_vc_sel_1_2_MPORT_data = io_enq_bits_vc_sel_1_2;
  assign ram_vc_sel_1_2_MPORT_addr = enq_ptr_value;
  assign ram_vc_sel_1_2_MPORT_mask = 1'h1;
  assign ram_vc_sel_1_2_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_vc_sel_1_3_io_deq_bits_MPORT_en = 1'h1;
  assign ram_vc_sel_1_3_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_vc_sel_1_3_io_deq_bits_MPORT_data = ram_vc_sel_1_3[ram_vc_sel_1_3_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_vc_sel_1_3_MPORT_data = io_enq_bits_vc_sel_1_3;
  assign ram_vc_sel_1_3_MPORT_addr = enq_ptr_value;
  assign ram_vc_sel_1_3_MPORT_mask = 1'h1;
  assign ram_vc_sel_1_3_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_vc_sel_0_0_io_deq_bits_MPORT_en = 1'h1;
  assign ram_vc_sel_0_0_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_vc_sel_0_0_io_deq_bits_MPORT_data = ram_vc_sel_0_0[ram_vc_sel_0_0_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_vc_sel_0_0_MPORT_data = io_enq_bits_vc_sel_0_0;
  assign ram_vc_sel_0_0_MPORT_addr = enq_ptr_value;
  assign ram_vc_sel_0_0_MPORT_mask = 1'h1;
  assign ram_vc_sel_0_0_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_vc_sel_0_1_io_deq_bits_MPORT_en = 1'h1;
  assign ram_vc_sel_0_1_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_vc_sel_0_1_io_deq_bits_MPORT_data = ram_vc_sel_0_1[ram_vc_sel_0_1_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_vc_sel_0_1_MPORT_data = io_enq_bits_vc_sel_0_1;
  assign ram_vc_sel_0_1_MPORT_addr = enq_ptr_value;
  assign ram_vc_sel_0_1_MPORT_mask = 1'h1;
  assign ram_vc_sel_0_1_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_vc_sel_0_2_io_deq_bits_MPORT_en = 1'h1;
  assign ram_vc_sel_0_2_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_vc_sel_0_2_io_deq_bits_MPORT_data = ram_vc_sel_0_2[ram_vc_sel_0_2_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_vc_sel_0_2_MPORT_data = io_enq_bits_vc_sel_0_2;
  assign ram_vc_sel_0_2_MPORT_addr = enq_ptr_value;
  assign ram_vc_sel_0_2_MPORT_mask = 1'h1;
  assign ram_vc_sel_0_2_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_vc_sel_0_3_io_deq_bits_MPORT_en = 1'h1;
  assign ram_vc_sel_0_3_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_vc_sel_0_3_io_deq_bits_MPORT_data = ram_vc_sel_0_3[ram_vc_sel_0_3_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_vc_sel_0_3_MPORT_data = io_enq_bits_vc_sel_0_3;
  assign ram_vc_sel_0_3_MPORT_addr = enq_ptr_value;
  assign ram_vc_sel_0_3_MPORT_mask = 1'h1;
  assign ram_vc_sel_0_3_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_vc_sel_1_0 = ram_vc_sel_1_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_vc_sel_1_1 = ram_vc_sel_1_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_vc_sel_1_2 = ram_vc_sel_1_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_vc_sel_1_3 = ram_vc_sel_1_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_vc_sel_0_0 = ram_vc_sel_0_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_vc_sel_0_1 = ram_vc_sel_0_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_vc_sel_0_2 = ram_vc_sel_0_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_vc_sel_0_3 = ram_vc_sel_0_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  always @(posedge clock) begin
    if (ram_vc_sel_1_0_MPORT_en & ram_vc_sel_1_0_MPORT_mask) begin
      ram_vc_sel_1_0[ram_vc_sel_1_0_MPORT_addr] <= ram_vc_sel_1_0_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_vc_sel_1_1_MPORT_en & ram_vc_sel_1_1_MPORT_mask) begin
      ram_vc_sel_1_1[ram_vc_sel_1_1_MPORT_addr] <= ram_vc_sel_1_1_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_vc_sel_1_2_MPORT_en & ram_vc_sel_1_2_MPORT_mask) begin
      ram_vc_sel_1_2[ram_vc_sel_1_2_MPORT_addr] <= ram_vc_sel_1_2_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_vc_sel_1_3_MPORT_en & ram_vc_sel_1_3_MPORT_mask) begin
      ram_vc_sel_1_3[ram_vc_sel_1_3_MPORT_addr] <= ram_vc_sel_1_3_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_vc_sel_0_0_MPORT_en & ram_vc_sel_0_0_MPORT_mask) begin
      ram_vc_sel_0_0[ram_vc_sel_0_0_MPORT_addr] <= ram_vc_sel_0_0_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_vc_sel_0_1_MPORT_en & ram_vc_sel_0_1_MPORT_mask) begin
      ram_vc_sel_0_1[ram_vc_sel_0_1_MPORT_addr] <= ram_vc_sel_0_1_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_vc_sel_0_2_MPORT_en & ram_vc_sel_0_2_MPORT_mask) begin
      ram_vc_sel_0_2[ram_vc_sel_0_2_MPORT_addr] <= ram_vc_sel_0_2_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_vc_sel_0_3_MPORT_en & ram_vc_sel_0_3_MPORT_mask) begin
      ram_vc_sel_0_3[ram_vc_sel_0_3_MPORT_addr] <= ram_vc_sel_0_3_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 1'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_vc_sel_1_0[initvar] = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_vc_sel_1_1[initvar] = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_vc_sel_1_2[initvar] = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_vc_sel_1_3[initvar] = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_vc_sel_0_0[initvar] = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_vc_sel_0_1[initvar] = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_vc_sel_0_2[initvar] = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_vc_sel_0_3[initvar] = _RAND_7[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  enq_ptr_value = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  deq_ptr_value = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  maybe_full = _RAND_10[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_3(
  input   clock,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input   io_enq_bits_vc_sel_1_0,
  input   io_enq_bits_vc_sel_1_1,
  input   io_enq_bits_vc_sel_1_2,
  input   io_enq_bits_vc_sel_1_3,
  input   io_enq_bits_vc_sel_0_0,
  input   io_enq_bits_vc_sel_0_1,
  input   io_enq_bits_vc_sel_0_2,
  input   io_enq_bits_vc_sel_0_3,
  input   io_deq_ready,
  output  io_deq_valid,
  output  io_deq_bits_vc_sel_1_0,
  output  io_deq_bits_vc_sel_1_1,
  output  io_deq_bits_vc_sel_1_2,
  output  io_deq_bits_vc_sel_1_3,
  output  io_deq_bits_vc_sel_0_0,
  output  io_deq_bits_vc_sel_0_1,
  output  io_deq_bits_vc_sel_0_2,
  output  io_deq_bits_vc_sel_0_3
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg  ram_vc_sel_1_0 [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_0_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_0_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_0_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_0_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_0_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_0_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_vc_sel_1_1 [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_1_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_1_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_1_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_1_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_1_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_1_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_vc_sel_1_2 [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_2_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_2_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_2_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_2_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_2_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_2_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_vc_sel_1_3 [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_3_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_3_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_3_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_3_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_3_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_1_3_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_vc_sel_0_0 [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_0_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_0_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_0_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_0_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_0_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_0_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_vc_sel_0_1 [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_1_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_1_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_1_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_1_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_1_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_1_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_vc_sel_0_2 [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_2_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_2_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_2_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_2_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_2_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_2_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_vc_sel_0_3 [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_3_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_3_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_3_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_3_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_3_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_vc_sel_0_3_MPORT_en; // @[Decoupled.scala 273:95]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 278:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  assign ram_vc_sel_1_0_io_deq_bits_MPORT_en = 1'h1;
  assign ram_vc_sel_1_0_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_vc_sel_1_0_io_deq_bits_MPORT_data = ram_vc_sel_1_0[ram_vc_sel_1_0_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_vc_sel_1_0_MPORT_data = io_enq_bits_vc_sel_1_0;
  assign ram_vc_sel_1_0_MPORT_addr = 1'h0;
  assign ram_vc_sel_1_0_MPORT_mask = 1'h1;
  assign ram_vc_sel_1_0_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_vc_sel_1_1_io_deq_bits_MPORT_en = 1'h1;
  assign ram_vc_sel_1_1_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_vc_sel_1_1_io_deq_bits_MPORT_data = ram_vc_sel_1_1[ram_vc_sel_1_1_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_vc_sel_1_1_MPORT_data = io_enq_bits_vc_sel_1_1;
  assign ram_vc_sel_1_1_MPORT_addr = 1'h0;
  assign ram_vc_sel_1_1_MPORT_mask = 1'h1;
  assign ram_vc_sel_1_1_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_vc_sel_1_2_io_deq_bits_MPORT_en = 1'h1;
  assign ram_vc_sel_1_2_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_vc_sel_1_2_io_deq_bits_MPORT_data = ram_vc_sel_1_2[ram_vc_sel_1_2_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_vc_sel_1_2_MPORT_data = io_enq_bits_vc_sel_1_2;
  assign ram_vc_sel_1_2_MPORT_addr = 1'h0;
  assign ram_vc_sel_1_2_MPORT_mask = 1'h1;
  assign ram_vc_sel_1_2_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_vc_sel_1_3_io_deq_bits_MPORT_en = 1'h1;
  assign ram_vc_sel_1_3_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_vc_sel_1_3_io_deq_bits_MPORT_data = ram_vc_sel_1_3[ram_vc_sel_1_3_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_vc_sel_1_3_MPORT_data = io_enq_bits_vc_sel_1_3;
  assign ram_vc_sel_1_3_MPORT_addr = 1'h0;
  assign ram_vc_sel_1_3_MPORT_mask = 1'h1;
  assign ram_vc_sel_1_3_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_vc_sel_0_0_io_deq_bits_MPORT_en = 1'h1;
  assign ram_vc_sel_0_0_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_vc_sel_0_0_io_deq_bits_MPORT_data = ram_vc_sel_0_0[ram_vc_sel_0_0_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_vc_sel_0_0_MPORT_data = io_enq_bits_vc_sel_0_0;
  assign ram_vc_sel_0_0_MPORT_addr = 1'h0;
  assign ram_vc_sel_0_0_MPORT_mask = 1'h1;
  assign ram_vc_sel_0_0_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_vc_sel_0_1_io_deq_bits_MPORT_en = 1'h1;
  assign ram_vc_sel_0_1_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_vc_sel_0_1_io_deq_bits_MPORT_data = ram_vc_sel_0_1[ram_vc_sel_0_1_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_vc_sel_0_1_MPORT_data = io_enq_bits_vc_sel_0_1;
  assign ram_vc_sel_0_1_MPORT_addr = 1'h0;
  assign ram_vc_sel_0_1_MPORT_mask = 1'h1;
  assign ram_vc_sel_0_1_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_vc_sel_0_2_io_deq_bits_MPORT_en = 1'h1;
  assign ram_vc_sel_0_2_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_vc_sel_0_2_io_deq_bits_MPORT_data = ram_vc_sel_0_2[ram_vc_sel_0_2_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_vc_sel_0_2_MPORT_data = io_enq_bits_vc_sel_0_2;
  assign ram_vc_sel_0_2_MPORT_addr = 1'h0;
  assign ram_vc_sel_0_2_MPORT_mask = 1'h1;
  assign ram_vc_sel_0_2_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_vc_sel_0_3_io_deq_bits_MPORT_en = 1'h1;
  assign ram_vc_sel_0_3_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_vc_sel_0_3_io_deq_bits_MPORT_data = ram_vc_sel_0_3[ram_vc_sel_0_3_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_vc_sel_0_3_MPORT_data = io_enq_bits_vc_sel_0_3;
  assign ram_vc_sel_0_3_MPORT_addr = 1'h0;
  assign ram_vc_sel_0_3_MPORT_mask = 1'h1;
  assign ram_vc_sel_0_3_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = io_deq_ready | empty; // @[Decoupled.scala 303:16 323:{24,39}]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_vc_sel_1_0 = ram_vc_sel_1_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_vc_sel_1_1 = ram_vc_sel_1_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_vc_sel_1_2 = ram_vc_sel_1_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_vc_sel_1_3 = ram_vc_sel_1_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_vc_sel_0_0 = ram_vc_sel_0_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_vc_sel_0_1 = ram_vc_sel_0_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_vc_sel_0_2 = ram_vc_sel_0_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_vc_sel_0_3 = ram_vc_sel_0_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  always @(posedge clock) begin
    if (ram_vc_sel_1_0_MPORT_en & ram_vc_sel_1_0_MPORT_mask) begin
      ram_vc_sel_1_0[ram_vc_sel_1_0_MPORT_addr] <= ram_vc_sel_1_0_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_vc_sel_1_1_MPORT_en & ram_vc_sel_1_1_MPORT_mask) begin
      ram_vc_sel_1_1[ram_vc_sel_1_1_MPORT_addr] <= ram_vc_sel_1_1_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_vc_sel_1_2_MPORT_en & ram_vc_sel_1_2_MPORT_mask) begin
      ram_vc_sel_1_2[ram_vc_sel_1_2_MPORT_addr] <= ram_vc_sel_1_2_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_vc_sel_1_3_MPORT_en & ram_vc_sel_1_3_MPORT_mask) begin
      ram_vc_sel_1_3[ram_vc_sel_1_3_MPORT_addr] <= ram_vc_sel_1_3_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_vc_sel_0_0_MPORT_en & ram_vc_sel_0_0_MPORT_mask) begin
      ram_vc_sel_0_0[ram_vc_sel_0_0_MPORT_addr] <= ram_vc_sel_0_0_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_vc_sel_0_1_MPORT_en & ram_vc_sel_0_1_MPORT_mask) begin
      ram_vc_sel_0_1[ram_vc_sel_0_1_MPORT_addr] <= ram_vc_sel_0_1_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_vc_sel_0_2_MPORT_en & ram_vc_sel_0_2_MPORT_mask) begin
      ram_vc_sel_0_2[ram_vc_sel_0_2_MPORT_addr] <= ram_vc_sel_0_2_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_vc_sel_0_3_MPORT_en & ram_vc_sel_0_3_MPORT_mask) begin
      ram_vc_sel_0_3[ram_vc_sel_0_3_MPORT_addr] <= ram_vc_sel_0_3_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_vc_sel_1_0[initvar] = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_vc_sel_1_1[initvar] = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_vc_sel_1_2[initvar] = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_vc_sel_1_3[initvar] = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_vc_sel_0_0[initvar] = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_vc_sel_0_1[initvar] = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_vc_sel_0_2[initvar] = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_vc_sel_0_3[initvar] = _RAND_7[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  maybe_full = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IngressUnit(
  input         clock,
  input         reset,
  output        io_router_req_valid,
  output [1:0]  io_router_req_bits_flow_ingress_node,
  output [1:0]  io_router_req_bits_flow_egress_node,
  input         io_router_resp_vc_sel_1_0,
  input         io_router_resp_vc_sel_1_1,
  input         io_router_resp_vc_sel_1_2,
  input         io_router_resp_vc_sel_1_3,
  input         io_router_resp_vc_sel_0_0,
  input         io_router_resp_vc_sel_0_1,
  input         io_router_resp_vc_sel_0_2,
  input         io_router_resp_vc_sel_0_3,
  input         io_vcalloc_req_ready,
  output        io_vcalloc_req_valid,
  output        io_vcalloc_req_bits_vc_sel_1_0,
  output        io_vcalloc_req_bits_vc_sel_1_1,
  output        io_vcalloc_req_bits_vc_sel_1_2,
  output        io_vcalloc_req_bits_vc_sel_1_3,
  output        io_vcalloc_req_bits_vc_sel_0_0,
  output        io_vcalloc_req_bits_vc_sel_0_1,
  output        io_vcalloc_req_bits_vc_sel_0_2,
  output        io_vcalloc_req_bits_vc_sel_0_3,
  input         io_vcalloc_resp_vc_sel_1_0,
  input         io_vcalloc_resp_vc_sel_1_1,
  input         io_vcalloc_resp_vc_sel_1_2,
  input         io_vcalloc_resp_vc_sel_1_3,
  input         io_vcalloc_resp_vc_sel_0_0,
  input         io_vcalloc_resp_vc_sel_0_1,
  input         io_vcalloc_resp_vc_sel_0_2,
  input         io_vcalloc_resp_vc_sel_0_3,
  input         io_out_credit_available_1_1,
  input         io_out_credit_available_1_2,
  input         io_out_credit_available_1_3,
  input         io_out_credit_available_0_1,
  input         io_out_credit_available_0_2,
  input         io_out_credit_available_0_3,
  input         io_salloc_req_0_ready,
  output        io_salloc_req_0_valid,
  output        io_salloc_req_0_bits_vc_sel_1_0,
  output        io_salloc_req_0_bits_vc_sel_1_1,
  output        io_salloc_req_0_bits_vc_sel_1_2,
  output        io_salloc_req_0_bits_vc_sel_1_3,
  output        io_salloc_req_0_bits_vc_sel_0_0,
  output        io_salloc_req_0_bits_vc_sel_0_1,
  output        io_salloc_req_0_bits_vc_sel_0_2,
  output        io_salloc_req_0_bits_vc_sel_0_3,
  output        io_salloc_req_0_bits_tail,
  output        io_out_0_valid,
  output        io_out_0_bits_flit_head,
  output        io_out_0_bits_flit_tail,
  output [63:0] io_out_0_bits_flit_payload,
  output [1:0]  io_out_0_bits_flit_flow_ingress_node,
  output [1:0]  io_out_0_bits_flit_flow_egress_node,
  output [1:0]  io_out_0_bits_out_virt_channel,
  output        io_in_ready,
  input         io_in_valid,
  input         io_in_bits_head,
  input         io_in_bits_tail,
  input  [63:0] io_in_bits_payload,
  input         io_in_bits_egress_id
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  route_buffer_clock; // @[IngressUnit.scala 26:28]
  wire  route_buffer_reset; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_enq_ready; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_enq_valid; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_enq_bits_head; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_enq_bits_tail; // @[IngressUnit.scala 26:28]
  wire [63:0] route_buffer_io_enq_bits_payload; // @[IngressUnit.scala 26:28]
  wire [1:0] route_buffer_io_enq_bits_flow_ingress_node; // @[IngressUnit.scala 26:28]
  wire [1:0] route_buffer_io_enq_bits_flow_egress_node; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_deq_ready; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_deq_valid; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_deq_bits_head; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_deq_bits_tail; // @[IngressUnit.scala 26:28]
  wire [63:0] route_buffer_io_deq_bits_payload; // @[IngressUnit.scala 26:28]
  wire [1:0] route_buffer_io_deq_bits_flow_ingress_node; // @[IngressUnit.scala 26:28]
  wire [1:0] route_buffer_io_deq_bits_flow_egress_node; // @[IngressUnit.scala 26:28]
  wire  route_q_clock; // @[IngressUnit.scala 27:23]
  wire  route_q_reset; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_ready; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_valid; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_1_0; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_1_1; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_1_2; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_1_3; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_0_0; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_0_1; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_0_2; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_0_3; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_ready; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_valid; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_1_0; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_1_1; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_1_2; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_1_3; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_0_0; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_0_1; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_0_2; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_0_3; // @[IngressUnit.scala 27:23]
  wire  vcalloc_buffer_clock; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_reset; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_enq_ready; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_enq_valid; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_enq_bits_head; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_enq_bits_tail; // @[IngressUnit.scala 75:30]
  wire [63:0] vcalloc_buffer_io_enq_bits_payload; // @[IngressUnit.scala 75:30]
  wire [1:0] vcalloc_buffer_io_enq_bits_flow_ingress_node; // @[IngressUnit.scala 75:30]
  wire [1:0] vcalloc_buffer_io_enq_bits_flow_egress_node; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_deq_ready; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_deq_valid; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_deq_bits_head; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_deq_bits_tail; // @[IngressUnit.scala 75:30]
  wire [63:0] vcalloc_buffer_io_deq_bits_payload; // @[IngressUnit.scala 75:30]
  wire [1:0] vcalloc_buffer_io_deq_bits_flow_ingress_node; // @[IngressUnit.scala 75:30]
  wire [1:0] vcalloc_buffer_io_deq_bits_flow_egress_node; // @[IngressUnit.scala 75:30]
  wire  vcalloc_q_clock; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_reset; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_ready; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_valid; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_1_0; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_1_1; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_1_2; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_1_3; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_0_0; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_0_1; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_0_2; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_0_3; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_ready; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_valid; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_1_0; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_1_1; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_1_2; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_1_3; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_0_0; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_0_1; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_0_2; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_0_3; // @[IngressUnit.scala 76:25]
  wire  _T = ~io_in_bits_egress_id; // @[IngressUnit.scala 30:72]
  wire  _T_2 = _T | io_in_bits_egress_id; // @[package.scala 73:59]
  wire  _T_7 = ~reset; // @[IngressUnit.scala 30:9]
  wire [1:0] _route_buffer_io_enq_bits_flow_egress_node_T_3 = io_in_bits_egress_id ? 2'h3 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _GEN_9 = {{1'd0}, _T}; // @[Mux.scala 27:73]
  wire  at_dest = route_buffer_io_enq_bits_flow_egress_node == 2'h0; // @[IngressUnit.scala 55:59]
  wire  _T_9 = io_in_ready & io_in_valid; // @[Decoupled.scala 51:35]
  wire  _vcalloc_buffer_io_enq_valid_T = ~route_buffer_io_deq_bits_head; // @[IngressUnit.scala 88:30]
  wire  _vcalloc_buffer_io_enq_valid_T_1 = route_q_io_deq_valid | ~route_buffer_io_deq_bits_head; // @[IngressUnit.scala 88:27]
  wire  _vcalloc_buffer_io_enq_valid_T_2 = route_buffer_io_deq_valid & _vcalloc_buffer_io_enq_valid_T_1; // @[IngressUnit.scala 87:61]
  wire  _vcalloc_buffer_io_enq_valid_T_4 = io_vcalloc_req_ready | _vcalloc_buffer_io_enq_valid_T; // @[IngressUnit.scala 89:27]
  wire  _io_vcalloc_req_valid_T_1 = route_buffer_io_deq_valid & route_q_io_deq_valid & route_buffer_io_deq_bits_head; // @[IngressUnit.scala 91:78]
  wire  _route_buffer_io_deq_ready_T_2 = vcalloc_buffer_io_enq_ready & _vcalloc_buffer_io_enq_valid_T_1; // @[IngressUnit.scala 93:61]
  wire  _route_buffer_io_deq_ready_T_5 = _route_buffer_io_deq_ready_T_2 & _vcalloc_buffer_io_enq_valid_T_4; // @[IngressUnit.scala 94:37]
  wire  _route_buffer_io_deq_ready_T_7 = vcalloc_q_io_enq_ready | _vcalloc_buffer_io_enq_valid_T; // @[IngressUnit.scala 96:29]
  wire  _route_q_io_deq_ready_T = route_buffer_io_deq_ready & route_buffer_io_deq_valid; // @[Decoupled.scala 51:35]
  wire [3:0] c_lo = {vcalloc_q_io_deq_bits_vc_sel_0_3,vcalloc_q_io_deq_bits_vc_sel_0_2,vcalloc_q_io_deq_bits_vc_sel_0_1,
    vcalloc_q_io_deq_bits_vc_sel_0_0}; // @[IngressUnit.scala 107:41]
  wire [3:0] c_hi = {vcalloc_q_io_deq_bits_vc_sel_1_3,vcalloc_q_io_deq_bits_vc_sel_1_2,vcalloc_q_io_deq_bits_vc_sel_1_1,
    vcalloc_q_io_deq_bits_vc_sel_1_0}; // @[IngressUnit.scala 107:41]
  wire [7:0] _c_T = {vcalloc_q_io_deq_bits_vc_sel_1_3,vcalloc_q_io_deq_bits_vc_sel_1_2,vcalloc_q_io_deq_bits_vc_sel_1_1,
    vcalloc_q_io_deq_bits_vc_sel_1_0,vcalloc_q_io_deq_bits_vc_sel_0_3,vcalloc_q_io_deq_bits_vc_sel_0_2,
    vcalloc_q_io_deq_bits_vc_sel_0_1,vcalloc_q_io_deq_bits_vc_sel_0_0}; // @[IngressUnit.scala 107:41]
  wire [7:0] _c_T_1 = {io_out_credit_available_1_3,io_out_credit_available_1_2,io_out_credit_available_1_1,1'h1,
    io_out_credit_available_0_3,io_out_credit_available_0_2,io_out_credit_available_0_1,1'h1}; // @[IngressUnit.scala 107:74]
  wire [7:0] _c_T_2 = _c_T & _c_T_1; // @[IngressUnit.scala 107:48]
  wire  c = _c_T_2 != 8'h0; // @[IngressUnit.scala 107:82]
  wire  _vcalloc_q_io_deq_ready_T = vcalloc_buffer_io_deq_ready & vcalloc_buffer_io_deq_valid; // @[Decoupled.scala 51:35]
  reg  out_bundle_valid; // @[IngressUnit.scala 116:8]
  reg  out_bundle_bits_flit_head; // @[IngressUnit.scala 116:8]
  reg  out_bundle_bits_flit_tail; // @[IngressUnit.scala 116:8]
  reg [63:0] out_bundle_bits_flit_payload; // @[IngressUnit.scala 116:8]
  reg [1:0] out_bundle_bits_flit_flow_ingress_node; // @[IngressUnit.scala 116:8]
  reg [1:0] out_bundle_bits_flit_flow_egress_node; // @[IngressUnit.scala 116:8]
  reg [1:0] out_bundle_bits_out_virt_channel; // @[IngressUnit.scala 116:8]
  wire  out_channel_oh_0 = vcalloc_q_io_deq_bits_vc_sel_0_0 | vcalloc_q_io_deq_bits_vc_sel_0_1 |
    vcalloc_q_io_deq_bits_vc_sel_0_2 | vcalloc_q_io_deq_bits_vc_sel_0_3; // @[IngressUnit.scala 123:67]
  wire  out_channel_oh_1 = vcalloc_q_io_deq_bits_vc_sel_1_0 | vcalloc_q_io_deq_bits_vc_sel_1_1 |
    vcalloc_q_io_deq_bits_vc_sel_1_2 | vcalloc_q_io_deq_bits_vc_sel_1_3; // @[IngressUnit.scala 123:67]
  wire [1:0] out_bundle_bits_out_virt_channel_hi_1 = c_lo[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] out_bundle_bits_out_virt_channel_lo_1 = c_lo[1:0]; // @[OneHot.scala 31:18]
  wire  _out_bundle_bits_out_virt_channel_T_1 = |out_bundle_bits_out_virt_channel_hi_1; // @[OneHot.scala 32:14]
  wire [1:0] _out_bundle_bits_out_virt_channel_T_2 = out_bundle_bits_out_virt_channel_hi_1 |
    out_bundle_bits_out_virt_channel_lo_1; // @[OneHot.scala 32:28]
  wire [1:0] _out_bundle_bits_out_virt_channel_T_4 = {_out_bundle_bits_out_virt_channel_T_1,
    _out_bundle_bits_out_virt_channel_T_2[1]}; // @[Cat.scala 33:92]
  wire [1:0] out_bundle_bits_out_virt_channel_hi_3 = c_hi[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] out_bundle_bits_out_virt_channel_lo_3 = c_hi[1:0]; // @[OneHot.scala 31:18]
  wire  _out_bundle_bits_out_virt_channel_T_6 = |out_bundle_bits_out_virt_channel_hi_3; // @[OneHot.scala 32:14]
  wire [1:0] _out_bundle_bits_out_virt_channel_T_7 = out_bundle_bits_out_virt_channel_hi_3 |
    out_bundle_bits_out_virt_channel_lo_3; // @[OneHot.scala 32:28]
  wire [1:0] _out_bundle_bits_out_virt_channel_T_9 = {_out_bundle_bits_out_virt_channel_T_6,
    _out_bundle_bits_out_virt_channel_T_7[1]}; // @[Cat.scala 33:92]
  wire [1:0] _out_bundle_bits_out_virt_channel_T_10 = out_channel_oh_0 ? _out_bundle_bits_out_virt_channel_T_4 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _out_bundle_bits_out_virt_channel_T_11 = out_channel_oh_1 ? _out_bundle_bits_out_virt_channel_T_9 : 2'h0; // @[Mux.scala 27:73]
  Queue route_buffer ( // @[IngressUnit.scala 26:28]
    .clock(route_buffer_clock),
    .reset(route_buffer_reset),
    .io_enq_ready(route_buffer_io_enq_ready),
    .io_enq_valid(route_buffer_io_enq_valid),
    .io_enq_bits_head(route_buffer_io_enq_bits_head),
    .io_enq_bits_tail(route_buffer_io_enq_bits_tail),
    .io_enq_bits_payload(route_buffer_io_enq_bits_payload),
    .io_enq_bits_flow_ingress_node(route_buffer_io_enq_bits_flow_ingress_node),
    .io_enq_bits_flow_egress_node(route_buffer_io_enq_bits_flow_egress_node),
    .io_deq_ready(route_buffer_io_deq_ready),
    .io_deq_valid(route_buffer_io_deq_valid),
    .io_deq_bits_head(route_buffer_io_deq_bits_head),
    .io_deq_bits_tail(route_buffer_io_deq_bits_tail),
    .io_deq_bits_payload(route_buffer_io_deq_bits_payload),
    .io_deq_bits_flow_ingress_node(route_buffer_io_deq_bits_flow_ingress_node),
    .io_deq_bits_flow_egress_node(route_buffer_io_deq_bits_flow_egress_node)
  );
  Queue_1 route_q ( // @[IngressUnit.scala 27:23]
    .clock(route_q_clock),
    .reset(route_q_reset),
    .io_enq_ready(route_q_io_enq_ready),
    .io_enq_valid(route_q_io_enq_valid),
    .io_enq_bits_vc_sel_1_0(route_q_io_enq_bits_vc_sel_1_0),
    .io_enq_bits_vc_sel_1_1(route_q_io_enq_bits_vc_sel_1_1),
    .io_enq_bits_vc_sel_1_2(route_q_io_enq_bits_vc_sel_1_2),
    .io_enq_bits_vc_sel_1_3(route_q_io_enq_bits_vc_sel_1_3),
    .io_enq_bits_vc_sel_0_0(route_q_io_enq_bits_vc_sel_0_0),
    .io_enq_bits_vc_sel_0_1(route_q_io_enq_bits_vc_sel_0_1),
    .io_enq_bits_vc_sel_0_2(route_q_io_enq_bits_vc_sel_0_2),
    .io_enq_bits_vc_sel_0_3(route_q_io_enq_bits_vc_sel_0_3),
    .io_deq_ready(route_q_io_deq_ready),
    .io_deq_valid(route_q_io_deq_valid),
    .io_deq_bits_vc_sel_1_0(route_q_io_deq_bits_vc_sel_1_0),
    .io_deq_bits_vc_sel_1_1(route_q_io_deq_bits_vc_sel_1_1),
    .io_deq_bits_vc_sel_1_2(route_q_io_deq_bits_vc_sel_1_2),
    .io_deq_bits_vc_sel_1_3(route_q_io_deq_bits_vc_sel_1_3),
    .io_deq_bits_vc_sel_0_0(route_q_io_deq_bits_vc_sel_0_0),
    .io_deq_bits_vc_sel_0_1(route_q_io_deq_bits_vc_sel_0_1),
    .io_deq_bits_vc_sel_0_2(route_q_io_deq_bits_vc_sel_0_2),
    .io_deq_bits_vc_sel_0_3(route_q_io_deq_bits_vc_sel_0_3)
  );
  Queue vcalloc_buffer ( // @[IngressUnit.scala 75:30]
    .clock(vcalloc_buffer_clock),
    .reset(vcalloc_buffer_reset),
    .io_enq_ready(vcalloc_buffer_io_enq_ready),
    .io_enq_valid(vcalloc_buffer_io_enq_valid),
    .io_enq_bits_head(vcalloc_buffer_io_enq_bits_head),
    .io_enq_bits_tail(vcalloc_buffer_io_enq_bits_tail),
    .io_enq_bits_payload(vcalloc_buffer_io_enq_bits_payload),
    .io_enq_bits_flow_ingress_node(vcalloc_buffer_io_enq_bits_flow_ingress_node),
    .io_enq_bits_flow_egress_node(vcalloc_buffer_io_enq_bits_flow_egress_node),
    .io_deq_ready(vcalloc_buffer_io_deq_ready),
    .io_deq_valid(vcalloc_buffer_io_deq_valid),
    .io_deq_bits_head(vcalloc_buffer_io_deq_bits_head),
    .io_deq_bits_tail(vcalloc_buffer_io_deq_bits_tail),
    .io_deq_bits_payload(vcalloc_buffer_io_deq_bits_payload),
    .io_deq_bits_flow_ingress_node(vcalloc_buffer_io_deq_bits_flow_ingress_node),
    .io_deq_bits_flow_egress_node(vcalloc_buffer_io_deq_bits_flow_egress_node)
  );
  Queue_3 vcalloc_q ( // @[IngressUnit.scala 76:25]
    .clock(vcalloc_q_clock),
    .reset(vcalloc_q_reset),
    .io_enq_ready(vcalloc_q_io_enq_ready),
    .io_enq_valid(vcalloc_q_io_enq_valid),
    .io_enq_bits_vc_sel_1_0(vcalloc_q_io_enq_bits_vc_sel_1_0),
    .io_enq_bits_vc_sel_1_1(vcalloc_q_io_enq_bits_vc_sel_1_1),
    .io_enq_bits_vc_sel_1_2(vcalloc_q_io_enq_bits_vc_sel_1_2),
    .io_enq_bits_vc_sel_1_3(vcalloc_q_io_enq_bits_vc_sel_1_3),
    .io_enq_bits_vc_sel_0_0(vcalloc_q_io_enq_bits_vc_sel_0_0),
    .io_enq_bits_vc_sel_0_1(vcalloc_q_io_enq_bits_vc_sel_0_1),
    .io_enq_bits_vc_sel_0_2(vcalloc_q_io_enq_bits_vc_sel_0_2),
    .io_enq_bits_vc_sel_0_3(vcalloc_q_io_enq_bits_vc_sel_0_3),
    .io_deq_ready(vcalloc_q_io_deq_ready),
    .io_deq_valid(vcalloc_q_io_deq_valid),
    .io_deq_bits_vc_sel_1_0(vcalloc_q_io_deq_bits_vc_sel_1_0),
    .io_deq_bits_vc_sel_1_1(vcalloc_q_io_deq_bits_vc_sel_1_1),
    .io_deq_bits_vc_sel_1_2(vcalloc_q_io_deq_bits_vc_sel_1_2),
    .io_deq_bits_vc_sel_1_3(vcalloc_q_io_deq_bits_vc_sel_1_3),
    .io_deq_bits_vc_sel_0_0(vcalloc_q_io_deq_bits_vc_sel_0_0),
    .io_deq_bits_vc_sel_0_1(vcalloc_q_io_deq_bits_vc_sel_0_1),
    .io_deq_bits_vc_sel_0_2(vcalloc_q_io_deq_bits_vc_sel_0_2),
    .io_deq_bits_vc_sel_0_3(vcalloc_q_io_deq_bits_vc_sel_0_3)
  );
  assign io_router_req_valid = io_in_valid & route_buffer_io_enq_ready & io_in_bits_head & ~at_dest; // @[IngressUnit.scala 58:86]
  assign io_router_req_bits_flow_ingress_node = route_buffer_io_enq_bits_flow_ingress_node; // @[IngressUnit.scala 53:27]
  assign io_router_req_bits_flow_egress_node = route_buffer_io_enq_bits_flow_egress_node; // @[IngressUnit.scala 53:27]
  assign io_vcalloc_req_valid = _io_vcalloc_req_valid_T_1 & vcalloc_buffer_io_enq_ready & vcalloc_q_io_enq_ready; // @[IngressUnit.scala 92:41]
  assign io_vcalloc_req_bits_vc_sel_1_0 = route_q_io_deq_bits_vc_sel_1_0; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_1_1 = route_q_io_deq_bits_vc_sel_1_1; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_1_2 = route_q_io_deq_bits_vc_sel_1_2; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_1_3 = route_q_io_deq_bits_vc_sel_1_3; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_0_0 = route_q_io_deq_bits_vc_sel_0_0; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_0_1 = route_q_io_deq_bits_vc_sel_0_1; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_0_2 = route_q_io_deq_bits_vc_sel_0_2; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_0_3 = route_q_io_deq_bits_vc_sel_0_3; // @[IngressUnit.scala 81:30]
  assign io_salloc_req_0_valid = vcalloc_buffer_io_deq_valid & vcalloc_q_io_deq_valid & c; // @[IngressUnit.scala 109:83]
  assign io_salloc_req_0_bits_vc_sel_1_0 = vcalloc_q_io_deq_bits_vc_sel_1_0; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_1_1 = vcalloc_q_io_deq_bits_vc_sel_1_1; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_1_2 = vcalloc_q_io_deq_bits_vc_sel_1_2; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_1_3 = vcalloc_q_io_deq_bits_vc_sel_1_3; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_0_0 = vcalloc_q_io_deq_bits_vc_sel_0_0; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_0_1 = vcalloc_q_io_deq_bits_vc_sel_0_1; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_0_2 = vcalloc_q_io_deq_bits_vc_sel_0_2; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_0_3 = vcalloc_q_io_deq_bits_vc_sel_0_3; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_tail = vcalloc_buffer_io_deq_bits_tail; // @[IngressUnit.scala 105:30]
  assign io_out_0_valid = out_bundle_valid; // @[IngressUnit.scala 118:13]
  assign io_out_0_bits_flit_head = out_bundle_bits_flit_head; // @[IngressUnit.scala 118:13]
  assign io_out_0_bits_flit_tail = out_bundle_bits_flit_tail; // @[IngressUnit.scala 118:13]
  assign io_out_0_bits_flit_payload = out_bundle_bits_flit_payload; // @[IngressUnit.scala 118:13]
  assign io_out_0_bits_flit_flow_ingress_node = out_bundle_bits_flit_flow_ingress_node; // @[IngressUnit.scala 118:13]
  assign io_out_0_bits_flit_flow_egress_node = out_bundle_bits_flit_flow_egress_node; // @[IngressUnit.scala 118:13]
  assign io_out_0_bits_out_virt_channel = out_bundle_bits_out_virt_channel; // @[IngressUnit.scala 118:13]
  assign io_in_ready = route_buffer_io_enq_ready; // @[IngressUnit.scala 59:44]
  assign route_buffer_clock = clock;
  assign route_buffer_reset = reset;
  assign route_buffer_io_enq_valid = io_in_valid; // @[IngressUnit.scala 56:44]
  assign route_buffer_io_enq_bits_head = io_in_bits_head; // @[IngressUnit.scala 32:33]
  assign route_buffer_io_enq_bits_tail = io_in_bits_tail; // @[IngressUnit.scala 33:33]
  assign route_buffer_io_enq_bits_payload = io_in_bits_payload; // @[IngressUnit.scala 50:36]
  assign route_buffer_io_enq_bits_flow_ingress_node = 2'h0; // @[IngressUnit.scala 38:51]
  assign route_buffer_io_enq_bits_flow_egress_node = _GEN_9 | _route_buffer_io_enq_bits_flow_egress_node_T_3; // @[Mux.scala 27:73]
  assign route_buffer_io_deq_ready = _route_buffer_io_deq_ready_T_5 & _route_buffer_io_deq_ready_T_7; // @[IngressUnit.scala 95:37]
  assign route_q_clock = clock;
  assign route_q_reset = reset;
  assign route_q_io_enq_valid = _T_9 & io_in_bits_head & at_dest | io_router_req_valid; // @[IngressUnit.scala 62:24 64:53 65:26]
  assign route_q_io_enq_bits_vc_sel_1_0 = _T_9 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_1_0; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_1_1 = _T_9 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_1_1; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_1_2 = _T_9 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_1_2; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_1_3 = _T_9 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_1_3; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_0_0 = _T_9 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_0_0; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_0_1 = _T_9 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_0_1; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_0_2 = _T_9 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_0_2; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_0_3 = _T_9 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_0_3; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_deq_ready = _route_q_io_deq_ready_T & route_buffer_io_deq_bits_tail; // @[IngressUnit.scala 97:55]
  assign vcalloc_buffer_clock = clock;
  assign vcalloc_buffer_reset = reset;
  assign vcalloc_buffer_io_enq_valid = _vcalloc_buffer_io_enq_valid_T_2 & _vcalloc_buffer_io_enq_valid_T_4; // @[IngressUnit.scala 88:37]
  assign vcalloc_buffer_io_enq_bits_head = route_buffer_io_deq_bits_head; // @[IngressUnit.scala 79:30]
  assign vcalloc_buffer_io_enq_bits_tail = route_buffer_io_deq_bits_tail; // @[IngressUnit.scala 79:30]
  assign vcalloc_buffer_io_enq_bits_payload = route_buffer_io_deq_bits_payload; // @[IngressUnit.scala 79:30]
  assign vcalloc_buffer_io_enq_bits_flow_ingress_node = route_buffer_io_deq_bits_flow_ingress_node; // @[IngressUnit.scala 79:30]
  assign vcalloc_buffer_io_enq_bits_flow_egress_node = route_buffer_io_deq_bits_flow_egress_node; // @[IngressUnit.scala 79:30]
  assign vcalloc_buffer_io_deq_ready = io_salloc_req_0_ready & vcalloc_q_io_deq_valid & c; // @[IngressUnit.scala 110:83]
  assign vcalloc_q_clock = clock;
  assign vcalloc_q_reset = reset;
  assign vcalloc_q_io_enq_valid = io_vcalloc_req_ready & io_vcalloc_req_valid; // @[Decoupled.scala 51:35]
  assign vcalloc_q_io_enq_bits_vc_sel_1_0 = io_vcalloc_resp_vc_sel_1_0; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_1_1 = io_vcalloc_resp_vc_sel_1_1; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_1_2 = io_vcalloc_resp_vc_sel_1_2; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_1_3 = io_vcalloc_resp_vc_sel_1_3; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_0_0 = io_vcalloc_resp_vc_sel_0_0; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_0_1 = io_vcalloc_resp_vc_sel_0_1; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_0_2 = io_vcalloc_resp_vc_sel_0_2; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_0_3 = io_vcalloc_resp_vc_sel_0_3; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_deq_ready = vcalloc_buffer_io_deq_bits_tail & _vcalloc_q_io_deq_ready_T; // @[IngressUnit.scala 111:42]
  always @(posedge clock) begin
    out_bundle_valid <= vcalloc_buffer_io_deq_ready & vcalloc_buffer_io_deq_valid; // @[Decoupled.scala 51:35]
    out_bundle_bits_flit_head <= vcalloc_buffer_io_deq_bits_head; // @[IngressUnit.scala 121:24]
    out_bundle_bits_flit_tail <= vcalloc_buffer_io_deq_bits_tail; // @[IngressUnit.scala 121:24]
    out_bundle_bits_flit_payload <= vcalloc_buffer_io_deq_bits_payload; // @[IngressUnit.scala 121:24]
    out_bundle_bits_flit_flow_ingress_node <= vcalloc_buffer_io_deq_bits_flow_ingress_node; // @[IngressUnit.scala 121:24]
    out_bundle_bits_flit_flow_egress_node <= vcalloc_buffer_io_deq_bits_flow_egress_node; // @[IngressUnit.scala 121:24]
    out_bundle_bits_out_virt_channel <= _out_bundle_bits_out_virt_channel_T_10 | _out_bundle_bits_out_virt_channel_T_11; // @[Mux.scala 27:73]
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~(io_in_valid & ~_T_2))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at IngressUnit.scala:30 assert(!(io.in.valid && !cParam.possibleFlows.toSeq.map(_.egressId.U === io.in.bits.egress_id).orR))\n"
            ); // @[IngressUnit.scala 30:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7 & ~(~(route_q_io_enq_valid & ~route_q_io_enq_ready))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at IngressUnit.scala:73 assert(!(route_q.io.enq.valid && !route_q.io.enq.ready))\n"); // @[IngressUnit.scala 73:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7 & ~(~(vcalloc_q_io_enq_valid & ~vcalloc_q_io_enq_ready))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at IngressUnit.scala:102 assert(!(vcalloc_q.io.enq.valid && !vcalloc_q.io.enq.ready))\n"
            ); // @[IngressUnit.scala 102:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  out_bundle_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  out_bundle_bits_flit_head = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  out_bundle_bits_flit_tail = _RAND_2[0:0];
  _RAND_3 = {2{`RANDOM}};
  out_bundle_bits_flit_payload = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  out_bundle_bits_flit_flow_ingress_node = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  out_bundle_bits_flit_flow_egress_node = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  out_bundle_bits_out_virt_channel = _RAND_6[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(~(io_in_valid & ~_T_2)); // @[IngressUnit.scala 30:9]
    end
    //
    if (_T_7) begin
      assert(~(route_q_io_enq_valid & ~route_q_io_enq_ready)); // @[IngressUnit.scala 73:9]
    end
    //
    if (_T_7) begin
      assert(~(vcalloc_q_io_enq_valid & ~vcalloc_q_io_enq_ready)); // @[IngressUnit.scala 102:9]
    end
  end
endmodule
module OutputUnit(
  input         clock,
  input         reset,
  input         io_in_0_valid,
  input         io_in_0_bits_head,
  input         io_in_0_bits_tail,
  input  [63:0] io_in_0_bits_payload,
  input  [1:0]  io_in_0_bits_flow_ingress_node,
  input  [1:0]  io_in_0_bits_flow_egress_node,
  input  [1:0]  io_in_0_bits_virt_channel_id,
  output        io_credit_available_1,
  output        io_credit_available_2,
  output        io_credit_available_3,
  output        io_channel_status_1_occupied,
  output        io_channel_status_2_occupied,
  output        io_channel_status_3_occupied,
  input         io_allocs_1_alloc,
  input         io_allocs_2_alloc,
  input         io_allocs_3_alloc,
  input         io_credit_alloc_1_alloc,
  input         io_credit_alloc_2_alloc,
  input         io_credit_alloc_3_alloc,
  output        io_out_flit_0_valid,
  output        io_out_flit_0_bits_head,
  output        io_out_flit_0_bits_tail,
  output [63:0] io_out_flit_0_bits_payload,
  output [1:0]  io_out_flit_0_bits_flow_ingress_node,
  output [1:0]  io_out_flit_0_bits_flow_egress_node,
  output [1:0]  io_out_flit_0_bits_virt_channel_id,
  input  [3:0]  io_out_credit_return,
  input  [3:0]  io_out_vc_free
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg  states_3_occupied; // @[OutputUnit.scala 66:19]
  reg [2:0] states_3_c; // @[OutputUnit.scala 66:19]
  reg  states_2_occupied; // @[OutputUnit.scala 66:19]
  reg [2:0] states_2_c; // @[OutputUnit.scala 66:19]
  reg  states_1_occupied; // @[OutputUnit.scala 66:19]
  reg [2:0] states_1_c; // @[OutputUnit.scala 66:19]
  wire  _GEN_0 = io_out_vc_free[1] ? 1'h0 : states_1_occupied; // @[OutputUnit.scala 74:30 76:18 66:19]
  wire  _GEN_1 = io_out_vc_free[2] ? 1'h0 : states_2_occupied; // @[OutputUnit.scala 74:30 76:18 66:19]
  wire  _GEN_2 = io_out_vc_free[3] ? 1'h0 : states_3_occupied; // @[OutputUnit.scala 74:30 76:18 66:19]
  wire  _GEN_3 = io_allocs_1_alloc | _GEN_0; // @[OutputUnit.scala 83:20 84:18]
  wire  _GEN_9 = io_allocs_2_alloc | _GEN_1; // @[OutputUnit.scala 83:20 84:18]
  wire  _GEN_15 = io_allocs_3_alloc | _GEN_2; // @[OutputUnit.scala 83:20 84:18]
  wire  free_1 = io_out_credit_return[1]; // @[OutputUnit.scala 94:36]
  wire [2:0] _GEN_4 = {{2'd0}, free_1}; // @[OutputUnit.scala 97:18]
  wire [3:0] _states_1_c_T = states_1_c + _GEN_4; // @[OutputUnit.scala 97:18]
  wire [3:0] _GEN_6 = {{3'd0}, io_credit_alloc_1_alloc}; // @[OutputUnit.scala 97:26]
  wire [3:0] _states_1_c_T_2 = _states_1_c_T - _GEN_6; // @[OutputUnit.scala 97:26]
  wire  free_2 = io_out_credit_return[2]; // @[OutputUnit.scala 94:36]
  wire [2:0] _GEN_8 = {{2'd0}, free_2}; // @[OutputUnit.scala 97:18]
  wire [3:0] _states_2_c_T = states_2_c + _GEN_8; // @[OutputUnit.scala 97:18]
  wire [3:0] _GEN_10 = {{3'd0}, io_credit_alloc_2_alloc}; // @[OutputUnit.scala 97:26]
  wire [3:0] _states_2_c_T_2 = _states_2_c_T - _GEN_10; // @[OutputUnit.scala 97:26]
  wire  free_3 = io_out_credit_return[3]; // @[OutputUnit.scala 94:36]
  wire [2:0] _GEN_12 = {{2'd0}, free_3}; // @[OutputUnit.scala 97:18]
  wire [3:0] _states_3_c_T = states_3_c + _GEN_12; // @[OutputUnit.scala 97:18]
  wire [3:0] _GEN_14 = {{3'd0}, io_credit_alloc_3_alloc}; // @[OutputUnit.scala 97:26]
  wire [3:0] _states_3_c_T_2 = _states_3_c_T - _GEN_14; // @[OutputUnit.scala 97:26]
  wire [3:0] _GEN_26 = reset ? 4'h5 : _states_1_c_T_2; // @[OutputUnit.scala 103:23 105:29 97:11]
  wire [3:0] _GEN_27 = reset ? 4'h5 : _states_2_c_T_2; // @[OutputUnit.scala 103:23 105:29 97:11]
  wire [3:0] _GEN_28 = reset ? 4'h5 : _states_3_c_T_2; // @[OutputUnit.scala 103:23 105:29 97:11]
  assign io_credit_available_1 = states_1_c != 3'h0; // @[OutputUnit.scala 90:14]
  assign io_credit_available_2 = states_2_c != 3'h0; // @[OutputUnit.scala 90:14]
  assign io_credit_available_3 = states_3_c != 3'h0; // @[OutputUnit.scala 90:14]
  assign io_channel_status_1_occupied = io_out_vc_free[1] ? 1'h0 : states_1_occupied; // @[OutputUnit.scala 74:30 76:18 66:19]
  assign io_channel_status_2_occupied = io_out_vc_free[2] ? 1'h0 : states_2_occupied; // @[OutputUnit.scala 74:30 76:18 66:19]
  assign io_channel_status_3_occupied = io_out_vc_free[3] ? 1'h0 : states_3_occupied; // @[OutputUnit.scala 74:30 76:18 66:19]
  assign io_out_flit_0_valid = io_in_0_valid; // @[OutputUnit.scala 71:15]
  assign io_out_flit_0_bits_head = io_in_0_bits_head; // @[OutputUnit.scala 71:15]
  assign io_out_flit_0_bits_tail = io_in_0_bits_tail; // @[OutputUnit.scala 71:15]
  assign io_out_flit_0_bits_payload = io_in_0_bits_payload; // @[OutputUnit.scala 71:15]
  assign io_out_flit_0_bits_flow_ingress_node = io_in_0_bits_flow_ingress_node; // @[OutputUnit.scala 71:15]
  assign io_out_flit_0_bits_flow_egress_node = io_in_0_bits_flow_egress_node; // @[OutputUnit.scala 71:15]
  assign io_out_flit_0_bits_virt_channel_id = io_in_0_bits_virt_channel_id; // @[OutputUnit.scala 71:15]
  always @(posedge clock) begin
    if (reset) begin // @[OutputUnit.scala 103:23]
      states_3_occupied <= 1'h0; // @[OutputUnit.scala 104:31]
    end else begin
      states_3_occupied <= _GEN_15;
    end
    states_3_c <= _GEN_28[2:0];
    if (reset) begin // @[OutputUnit.scala 103:23]
      states_2_occupied <= 1'h0; // @[OutputUnit.scala 104:31]
    end else begin
      states_2_occupied <= _GEN_9;
    end
    states_2_c <= _GEN_27[2:0];
    if (reset) begin // @[OutputUnit.scala 103:23]
      states_1_occupied <= 1'h0; // @[OutputUnit.scala 104:31]
    end else begin
      states_1_occupied <= _GEN_3;
    end
    states_1_c <= _GEN_26[2:0];
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_out_vc_free[1] & ~reset & ~states_1_occupied) begin
          $fwrite(32'h80000002,"Assertion failed\n    at OutputUnit.scala:75 assert(s.occupied)\n"); // @[OutputUnit.scala 75:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_out_vc_free[2] & ~reset & ~states_2_occupied) begin
          $fwrite(32'h80000002,"Assertion failed\n    at OutputUnit.scala:75 assert(s.occupied)\n"); // @[OutputUnit.scala 75:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_out_vc_free[3] & ~reset & ~states_3_occupied) begin
          $fwrite(32'h80000002,"Assertion failed\n    at OutputUnit.scala:75 assert(s.occupied)\n"); // @[OutputUnit.scala 75:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  states_3_occupied = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  states_3_c = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  states_2_occupied = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  states_2_c = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  states_1_occupied = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  states_1_c = _RAND_5[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (io_out_vc_free[1] & ~reset) begin
      assert(states_1_occupied); // @[OutputUnit.scala 75:13]
    end
    //
    if (io_out_vc_free[2] & ~reset) begin
      assert(states_2_occupied); // @[OutputUnit.scala 75:13]
    end
    //
    if (io_out_vc_free[3] & ~reset) begin
      assert(states_3_occupied); // @[OutputUnit.scala 75:13]
    end
  end
endmodule
module Switch(
  input         clock,
  input         reset,
  input         io_in_0_0_valid,
  input         io_in_0_0_bits_flit_head,
  input         io_in_0_0_bits_flit_tail,
  input  [63:0] io_in_0_0_bits_flit_payload,
  input  [1:0]  io_in_0_0_bits_flit_flow_ingress_node,
  input  [1:0]  io_in_0_0_bits_flit_flow_egress_node,
  input  [1:0]  io_in_0_0_bits_out_virt_channel,
  output        io_out_1_0_valid,
  output        io_out_1_0_bits_head,
  output        io_out_1_0_bits_tail,
  output [63:0] io_out_1_0_bits_payload,
  output [1:0]  io_out_1_0_bits_flow_ingress_node,
  output [1:0]  io_out_1_0_bits_flow_egress_node,
  output [1:0]  io_out_1_0_bits_virt_channel_id,
  output        io_out_0_0_valid,
  output        io_out_0_0_bits_head,
  output        io_out_0_0_bits_tail,
  output [63:0] io_out_0_0_bits_payload,
  output [1:0]  io_out_0_0_bits_flow_ingress_node,
  output [1:0]  io_out_0_0_bits_flow_egress_node,
  output [1:0]  io_out_0_0_bits_virt_channel_id,
  input         io_sel_1_0_0_0,
  input         io_sel_0_0_0_0
);
  assign io_out_1_0_valid = io_in_0_0_valid & io_sel_1_0_0_0; // @[Switch.scala 48:67]
  assign io_out_1_0_bits_head = io_in_0_0_bits_flit_head; // @[Switch.scala 36:21 40:18]
  assign io_out_1_0_bits_tail = io_in_0_0_bits_flit_tail; // @[Switch.scala 36:21 40:18]
  assign io_out_1_0_bits_payload = io_in_0_0_bits_flit_payload; // @[Switch.scala 36:21 40:18]
  assign io_out_1_0_bits_flow_ingress_node = io_in_0_0_bits_flit_flow_ingress_node; // @[Switch.scala 36:21 40:18]
  assign io_out_1_0_bits_flow_egress_node = io_in_0_0_bits_flit_flow_egress_node; // @[Switch.scala 36:21 40:18]
  assign io_out_1_0_bits_virt_channel_id = io_in_0_0_bits_out_virt_channel; // @[Switch.scala 36:21 40:18]
  assign io_out_0_0_valid = io_in_0_0_valid & io_sel_0_0_0_0; // @[Switch.scala 48:67]
  assign io_out_0_0_bits_head = io_in_0_0_bits_flit_head; // @[Switch.scala 36:21 40:18]
  assign io_out_0_0_bits_tail = io_in_0_0_bits_flit_tail; // @[Switch.scala 36:21 40:18]
  assign io_out_0_0_bits_payload = io_in_0_0_bits_flit_payload; // @[Switch.scala 36:21 40:18]
  assign io_out_0_0_bits_flow_ingress_node = io_in_0_0_bits_flit_flow_ingress_node; // @[Switch.scala 36:21 40:18]
  assign io_out_0_0_bits_flow_egress_node = io_in_0_0_bits_flit_flow_egress_node; // @[Switch.scala 36:21 40:18]
  assign io_out_0_0_bits_virt_channel_id = io_in_0_0_bits_out_virt_channel; // @[Switch.scala 36:21 40:18]
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(1'h1); // @[Switch.scala 47:13]
    end
    //
    if (~reset) begin
      assert(1'h1); // @[Switch.scala 47:13]
    end
  end
endmodule
module SwitchArbiter(
  input   clock,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input   io_in_0_bits_vc_sel_1_1,
  input   io_in_0_bits_vc_sel_1_2,
  input   io_in_0_bits_vc_sel_1_3,
  input   io_in_0_bits_vc_sel_0_1,
  input   io_in_0_bits_vc_sel_0_2,
  input   io_in_0_bits_vc_sel_0_3,
  input   io_in_0_bits_tail,
  output  io_out_0_valid,
  output  io_out_0_bits_vc_sel_1_1,
  output  io_out_0_bits_vc_sel_1_2,
  output  io_out_0_bits_vc_sel_1_3,
  output  io_out_0_bits_vc_sel_0_1,
  output  io_out_0_bits_vc_sel_0_2,
  output  io_out_0_bits_vc_sel_0_3,
  output  io_chosen_oh_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  lock_0; // @[SwitchAllocator.scala 24:38]
  wire  unassigned = io_in_0_valid & ~lock_0; // @[SwitchAllocator.scala 25:52]
  reg  mask; // @[SwitchAllocator.scala 27:21]
  wire  _sel_T = ~mask; // @[SwitchAllocator.scala 30:60]
  wire  _sel_T_1 = unassigned & ~mask; // @[SwitchAllocator.scala 30:58]
  wire [1:0] _sel_T_2 = {unassigned,_sel_T_1}; // @[Cat.scala 33:92]
  wire [1:0] _sel_T_5 = _sel_T_2[1] ? 2'h2 : 2'h0; // @[Mux.scala 47:70]
  wire [1:0] sel = _sel_T_2[0] ? 2'h1 : _sel_T_5; // @[Mux.scala 47:70]
  wire [1:0] _GEN_3 = {{1'd0}, sel[1]}; // @[SwitchAllocator.scala 32:23]
  wire [1:0] _choices_0_T_1 = sel | _GEN_3; // @[SwitchAllocator.scala 32:23]
  wire  choices_0 = _choices_0_T_1[0]; // @[SwitchAllocator.scala 28:21 32:16]
  wire  chosen = |(io_in_0_valid & lock_0) ? lock_0 : choices_0; // @[SwitchAllocator.scala 42:21]
  wire [1:0] _mask_T_3 = {mask, 1'h0}; // @[SwitchAllocator.scala 60:43]
  wire [1:0] _mask_T_4 = _mask_T_3 | 2'h1; // @[SwitchAllocator.scala 60:49]
  wire [1:0] _mask_T_5 = ~_sel_T ? 2'h0 : _mask_T_4; // @[SwitchAllocator.scala 60:16]
  wire [1:0] _GEN_2 = io_out_0_valid ? {{1'd0}, io_chosen_oh_0} : _mask_T_5; // @[SwitchAllocator.scala 57:27 58:10 60:10]
  wire [1:0] _GEN_4 = reset ? 2'h0 : _GEN_2; // @[SwitchAllocator.scala 27:{21,21}]
  assign io_in_0_ready = |(io_in_0_valid & lock_0) ? lock_0 : choices_0; // @[SwitchAllocator.scala 42:21]
  assign io_out_0_valid = |(io_in_0_valid & chosen); // @[SwitchAllocator.scala 44:45]
  assign io_out_0_bits_vc_sel_1_1 = io_in_0_bits_vc_sel_1_1; // @[SwitchAllocator.scala 45:20]
  assign io_out_0_bits_vc_sel_1_2 = io_in_0_bits_vc_sel_1_2; // @[SwitchAllocator.scala 45:20]
  assign io_out_0_bits_vc_sel_1_3 = io_in_0_bits_vc_sel_1_3; // @[SwitchAllocator.scala 45:20]
  assign io_out_0_bits_vc_sel_0_1 = io_in_0_bits_vc_sel_0_1; // @[SwitchAllocator.scala 45:20]
  assign io_out_0_bits_vc_sel_0_2 = io_in_0_bits_vc_sel_0_2; // @[SwitchAllocator.scala 45:20]
  assign io_out_0_bits_vc_sel_0_3 = io_in_0_bits_vc_sel_0_3; // @[SwitchAllocator.scala 45:20]
  assign io_chosen_oh_0 = |(io_in_0_valid & lock_0) ? lock_0 : choices_0; // @[SwitchAllocator.scala 42:21]
  always @(posedge clock) begin
    if (reset) begin // @[SwitchAllocator.scala 24:38]
      lock_0 <= 1'h0; // @[SwitchAllocator.scala 24:38]
    end else if (io_out_0_valid) begin // @[SwitchAllocator.scala 52:29]
      lock_0 <= chosen & ~io_in_0_bits_tail; // @[SwitchAllocator.scala 53:15]
    end
    mask <= _GEN_4[0]; // @[SwitchAllocator.scala 27:{21,21}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lock_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  mask = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SwitchAllocator(
  input   clock,
  input   reset,
  output  io_req_0_0_ready,
  input   io_req_0_0_valid,
  input   io_req_0_0_bits_vc_sel_1_0,
  input   io_req_0_0_bits_vc_sel_1_1,
  input   io_req_0_0_bits_vc_sel_1_2,
  input   io_req_0_0_bits_vc_sel_1_3,
  input   io_req_0_0_bits_vc_sel_0_0,
  input   io_req_0_0_bits_vc_sel_0_1,
  input   io_req_0_0_bits_vc_sel_0_2,
  input   io_req_0_0_bits_vc_sel_0_3,
  input   io_req_0_0_bits_tail,
  output  io_credit_alloc_1_1_alloc,
  output  io_credit_alloc_1_2_alloc,
  output  io_credit_alloc_1_3_alloc,
  output  io_credit_alloc_0_1_alloc,
  output  io_credit_alloc_0_2_alloc,
  output  io_credit_alloc_0_3_alloc,
  output  io_switch_sel_1_0_0_0,
  output  io_switch_sel_0_0_0_0
);
  wire  arbs_0_clock; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_reset; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_0_ready; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_0_valid; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_0_bits_vc_sel_1_1; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_0_bits_vc_sel_1_2; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_0_bits_vc_sel_1_3; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_0_bits_vc_sel_0_1; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_0_bits_vc_sel_0_2; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_0_bits_vc_sel_0_3; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_0_bits_tail; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_out_0_valid; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_out_0_bits_vc_sel_1_1; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_out_0_bits_vc_sel_1_2; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_out_0_bits_vc_sel_1_3; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_out_0_bits_vc_sel_0_1; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_out_0_bits_vc_sel_0_2; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_out_0_bits_vc_sel_0_3; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_chosen_oh_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_clock; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_reset; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_0_ready; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_0_valid; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_0_bits_vc_sel_1_1; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_0_bits_vc_sel_1_2; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_0_bits_vc_sel_1_3; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_0_bits_vc_sel_0_1; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_0_bits_vc_sel_0_2; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_0_bits_vc_sel_0_3; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_in_0_bits_tail; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_out_0_valid; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_out_0_bits_vc_sel_1_1; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_out_0_bits_vc_sel_1_2; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_out_0_bits_vc_sel_1_3; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_out_0_bits_vc_sel_0_1; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_out_0_bits_vc_sel_0_2; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_out_0_bits_vc_sel_0_3; // @[SwitchAllocator.scala 83:45]
  wire  arbs_1_io_chosen_oh_0; // @[SwitchAllocator.scala 83:45]
  wire  fires_0 = arbs_0_io_in_0_ready & arbs_0_io_in_0_valid; // @[Decoupled.scala 51:35]
  wire  fires_1 = arbs_1_io_in_0_ready & arbs_1_io_in_0_valid; // @[Decoupled.scala 51:35]
  SwitchArbiter arbs_0 ( // @[SwitchAllocator.scala 83:45]
    .clock(arbs_0_clock),
    .reset(arbs_0_reset),
    .io_in_0_ready(arbs_0_io_in_0_ready),
    .io_in_0_valid(arbs_0_io_in_0_valid),
    .io_in_0_bits_vc_sel_1_1(arbs_0_io_in_0_bits_vc_sel_1_1),
    .io_in_0_bits_vc_sel_1_2(arbs_0_io_in_0_bits_vc_sel_1_2),
    .io_in_0_bits_vc_sel_1_3(arbs_0_io_in_0_bits_vc_sel_1_3),
    .io_in_0_bits_vc_sel_0_1(arbs_0_io_in_0_bits_vc_sel_0_1),
    .io_in_0_bits_vc_sel_0_2(arbs_0_io_in_0_bits_vc_sel_0_2),
    .io_in_0_bits_vc_sel_0_3(arbs_0_io_in_0_bits_vc_sel_0_3),
    .io_in_0_bits_tail(arbs_0_io_in_0_bits_tail),
    .io_out_0_valid(arbs_0_io_out_0_valid),
    .io_out_0_bits_vc_sel_1_1(arbs_0_io_out_0_bits_vc_sel_1_1),
    .io_out_0_bits_vc_sel_1_2(arbs_0_io_out_0_bits_vc_sel_1_2),
    .io_out_0_bits_vc_sel_1_3(arbs_0_io_out_0_bits_vc_sel_1_3),
    .io_out_0_bits_vc_sel_0_1(arbs_0_io_out_0_bits_vc_sel_0_1),
    .io_out_0_bits_vc_sel_0_2(arbs_0_io_out_0_bits_vc_sel_0_2),
    .io_out_0_bits_vc_sel_0_3(arbs_0_io_out_0_bits_vc_sel_0_3),
    .io_chosen_oh_0(arbs_0_io_chosen_oh_0)
  );
  SwitchArbiter arbs_1 ( // @[SwitchAllocator.scala 83:45]
    .clock(arbs_1_clock),
    .reset(arbs_1_reset),
    .io_in_0_ready(arbs_1_io_in_0_ready),
    .io_in_0_valid(arbs_1_io_in_0_valid),
    .io_in_0_bits_vc_sel_1_1(arbs_1_io_in_0_bits_vc_sel_1_1),
    .io_in_0_bits_vc_sel_1_2(arbs_1_io_in_0_bits_vc_sel_1_2),
    .io_in_0_bits_vc_sel_1_3(arbs_1_io_in_0_bits_vc_sel_1_3),
    .io_in_0_bits_vc_sel_0_1(arbs_1_io_in_0_bits_vc_sel_0_1),
    .io_in_0_bits_vc_sel_0_2(arbs_1_io_in_0_bits_vc_sel_0_2),
    .io_in_0_bits_vc_sel_0_3(arbs_1_io_in_0_bits_vc_sel_0_3),
    .io_in_0_bits_tail(arbs_1_io_in_0_bits_tail),
    .io_out_0_valid(arbs_1_io_out_0_valid),
    .io_out_0_bits_vc_sel_1_1(arbs_1_io_out_0_bits_vc_sel_1_1),
    .io_out_0_bits_vc_sel_1_2(arbs_1_io_out_0_bits_vc_sel_1_2),
    .io_out_0_bits_vc_sel_1_3(arbs_1_io_out_0_bits_vc_sel_1_3),
    .io_out_0_bits_vc_sel_0_1(arbs_1_io_out_0_bits_vc_sel_0_1),
    .io_out_0_bits_vc_sel_0_2(arbs_1_io_out_0_bits_vc_sel_0_2),
    .io_out_0_bits_vc_sel_0_3(arbs_1_io_out_0_bits_vc_sel_0_3),
    .io_chosen_oh_0(arbs_1_io_chosen_oh_0)
  );
  assign io_req_0_0_ready = fires_0 | fires_1; // @[SwitchAllocator.scala 99:30]
  assign io_credit_alloc_1_1_alloc = arbs_1_io_out_0_valid & arbs_1_io_out_0_bits_vc_sel_1_1; // @[SwitchAllocator.scala 120:33]
  assign io_credit_alloc_1_2_alloc = arbs_1_io_out_0_valid & arbs_1_io_out_0_bits_vc_sel_1_2; // @[SwitchAllocator.scala 120:33]
  assign io_credit_alloc_1_3_alloc = arbs_1_io_out_0_valid & arbs_1_io_out_0_bits_vc_sel_1_3; // @[SwitchAllocator.scala 120:33]
  assign io_credit_alloc_0_1_alloc = arbs_0_io_out_0_valid & arbs_0_io_out_0_bits_vc_sel_0_1; // @[SwitchAllocator.scala 120:33]
  assign io_credit_alloc_0_2_alloc = arbs_0_io_out_0_valid & arbs_0_io_out_0_bits_vc_sel_0_2; // @[SwitchAllocator.scala 120:33]
  assign io_credit_alloc_0_3_alloc = arbs_0_io_out_0_valid & arbs_0_io_out_0_bits_vc_sel_0_3; // @[SwitchAllocator.scala 120:33]
  assign io_switch_sel_1_0_0_0 = arbs_1_io_in_0_valid & arbs_1_io_chosen_oh_0 & arbs_1_io_out_0_valid; // @[SwitchAllocator.scala 108:97]
  assign io_switch_sel_0_0_0_0 = arbs_0_io_in_0_valid & arbs_0_io_chosen_oh_0 & arbs_0_io_out_0_valid; // @[SwitchAllocator.scala 108:97]
  assign arbs_0_clock = clock;
  assign arbs_0_reset = reset;
  assign arbs_0_io_in_0_valid = io_req_0_0_valid & (io_req_0_0_bits_vc_sel_0_0 | io_req_0_0_bits_vc_sel_0_1 |
    io_req_0_0_bits_vc_sel_0_2 | io_req_0_0_bits_vc_sel_0_3); // @[SwitchAllocator.scala 95:37]
  assign arbs_0_io_in_0_bits_vc_sel_1_1 = io_req_0_0_bits_vc_sel_1_1; // @[SwitchAllocator.scala 96:25]
  assign arbs_0_io_in_0_bits_vc_sel_1_2 = io_req_0_0_bits_vc_sel_1_2; // @[SwitchAllocator.scala 96:25]
  assign arbs_0_io_in_0_bits_vc_sel_1_3 = io_req_0_0_bits_vc_sel_1_3; // @[SwitchAllocator.scala 96:25]
  assign arbs_0_io_in_0_bits_vc_sel_0_1 = io_req_0_0_bits_vc_sel_0_1; // @[SwitchAllocator.scala 96:25]
  assign arbs_0_io_in_0_bits_vc_sel_0_2 = io_req_0_0_bits_vc_sel_0_2; // @[SwitchAllocator.scala 96:25]
  assign arbs_0_io_in_0_bits_vc_sel_0_3 = io_req_0_0_bits_vc_sel_0_3; // @[SwitchAllocator.scala 96:25]
  assign arbs_0_io_in_0_bits_tail = io_req_0_0_bits_tail; // @[SwitchAllocator.scala 96:25]
  assign arbs_1_clock = clock;
  assign arbs_1_reset = reset;
  assign arbs_1_io_in_0_valid = io_req_0_0_valid & (io_req_0_0_bits_vc_sel_1_0 | io_req_0_0_bits_vc_sel_1_1 |
    io_req_0_0_bits_vc_sel_1_2 | io_req_0_0_bits_vc_sel_1_3); // @[SwitchAllocator.scala 95:37]
  assign arbs_1_io_in_0_bits_vc_sel_1_1 = io_req_0_0_bits_vc_sel_1_1; // @[SwitchAllocator.scala 96:25]
  assign arbs_1_io_in_0_bits_vc_sel_1_2 = io_req_0_0_bits_vc_sel_1_2; // @[SwitchAllocator.scala 96:25]
  assign arbs_1_io_in_0_bits_vc_sel_1_3 = io_req_0_0_bits_vc_sel_1_3; // @[SwitchAllocator.scala 96:25]
  assign arbs_1_io_in_0_bits_vc_sel_0_1 = io_req_0_0_bits_vc_sel_0_1; // @[SwitchAllocator.scala 96:25]
  assign arbs_1_io_in_0_bits_vc_sel_0_2 = io_req_0_0_bits_vc_sel_0_2; // @[SwitchAllocator.scala 96:25]
  assign arbs_1_io_in_0_bits_vc_sel_0_3 = io_req_0_0_bits_vc_sel_0_3; // @[SwitchAllocator.scala 96:25]
  assign arbs_1_io_in_0_bits_tail = io_req_0_0_bits_tail; // @[SwitchAllocator.scala 96:25]
endmodule
module RotatingSingleVCAllocator(
  input   clock,
  input   reset,
  output  io_req_0_ready,
  input   io_req_0_valid,
  input   io_req_0_bits_vc_sel_1_0,
  input   io_req_0_bits_vc_sel_1_1,
  input   io_req_0_bits_vc_sel_1_2,
  input   io_req_0_bits_vc_sel_1_3,
  input   io_req_0_bits_vc_sel_0_0,
  input   io_req_0_bits_vc_sel_0_1,
  input   io_req_0_bits_vc_sel_0_2,
  input   io_req_0_bits_vc_sel_0_3,
  output  io_resp_0_vc_sel_1_0,
  output  io_resp_0_vc_sel_1_1,
  output  io_resp_0_vc_sel_1_2,
  output  io_resp_0_vc_sel_1_3,
  output  io_resp_0_vc_sel_0_0,
  output  io_resp_0_vc_sel_0_1,
  output  io_resp_0_vc_sel_0_2,
  output  io_resp_0_vc_sel_0_3,
  input   io_channel_status_1_1_occupied,
  input   io_channel_status_1_2_occupied,
  input   io_channel_status_1_3_occupied,
  input   io_channel_status_0_1_occupied,
  input   io_channel_status_0_2_occupied,
  input   io_channel_status_0_3_occupied,
  output  io_out_allocs_1_1_alloc,
  output  io_out_allocs_1_2_alloc,
  output  io_out_allocs_1_3_alloc,
  output  io_out_allocs_0_1_alloc,
  output  io_out_allocs_0_2_alloc,
  output  io_out_allocs_0_3_alloc
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  mask; // @[SingleVCAllocator.scala 16:21]
  wire  in_arb_reqs_0_0_1 = io_req_0_bits_vc_sel_0_1 & ~io_channel_status_0_1_occupied; // @[SingleVCAllocator.scala 28:61]
  wire  in_arb_reqs_0_0_2 = io_req_0_bits_vc_sel_0_2 & ~io_channel_status_0_2_occupied; // @[SingleVCAllocator.scala 28:61]
  wire  in_arb_reqs_0_0_3 = io_req_0_bits_vc_sel_0_3 & ~io_channel_status_0_3_occupied; // @[SingleVCAllocator.scala 28:61]
  wire  in_arb_reqs_0_1_1 = io_req_0_bits_vc_sel_1_1 & ~io_channel_status_1_1_occupied; // @[SingleVCAllocator.scala 28:61]
  wire  in_arb_reqs_0_1_2 = io_req_0_bits_vc_sel_1_2 & ~io_channel_status_1_2_occupied; // @[SingleVCAllocator.scala 28:61]
  wire  in_arb_reqs_0_1_3 = io_req_0_bits_vc_sel_1_3 & ~io_channel_status_1_3_occupied; // @[SingleVCAllocator.scala 28:61]
  wire  _in_arb_vals_0_T_6 = io_req_0_bits_vc_sel_0_0 | in_arb_reqs_0_0_1 | in_arb_reqs_0_0_2 | in_arb_reqs_0_0_3 | (
    io_req_0_bits_vc_sel_1_0 | in_arb_reqs_0_1_1 | in_arb_reqs_0_1_2 | in_arb_reqs_0_1_3); // @[package.scala 73:59]
  wire  in_arb_vals_0 = io_req_0_valid & _in_arb_vals_0_T_6; // @[SingleVCAllocator.scala 32:39]
  wire  _in_arb_filter_T_1 = in_arb_vals_0 & ~mask; // @[SingleVCAllocator.scala 19:84]
  wire [1:0] _in_arb_filter_T_2 = {in_arb_vals_0,_in_arb_filter_T_1}; // @[Cat.scala 33:92]
  wire [1:0] _in_arb_filter_T_5 = _in_arb_filter_T_2[1] ? 2'h2 : 2'h0; // @[Mux.scala 47:70]
  wire [1:0] in_arb_filter = _in_arb_filter_T_2[0] ? 2'h1 : _in_arb_filter_T_5; // @[Mux.scala 47:70]
  wire  _GEN_0 = in_arb_vals_0 | mask; // @[SingleVCAllocator.scala 21:26 22:10 16:21]
  wire  _in_alloc_T = io_req_0_ready & io_req_0_valid; // @[Decoupled.scala 51:35]
  wire [7:0] _in_alloc_T_1 = {in_arb_reqs_0_1_3,in_arb_reqs_0_1_2,in_arb_reqs_0_1_1,io_req_0_bits_vc_sel_1_0,
    in_arb_reqs_0_0_3,in_arb_reqs_0_0_2,in_arb_reqs_0_0_1,io_req_0_bits_vc_sel_0_0}; // @[ISLIP.scala 33:18]
  reg [7:0] in_alloc_mask; // @[ISLIP.scala 17:25]
  wire [7:0] _in_alloc_full_T = ~in_alloc_mask; // @[ISLIP.scala 18:31]
  wire [7:0] _in_alloc_full_T_1 = _in_alloc_T_1 & _in_alloc_full_T; // @[ISLIP.scala 18:29]
  wire [15:0] in_alloc_full = {in_arb_reqs_0_1_3,in_arb_reqs_0_1_2,in_arb_reqs_0_1_1,io_req_0_bits_vc_sel_1_0,
    in_arb_reqs_0_0_3,in_arb_reqs_0_0_2,in_arb_reqs_0_0_1,io_req_0_bits_vc_sel_0_0,_in_alloc_full_T_1}; // @[Cat.scala 33:92]
  wire [15:0] _in_alloc_oh_T_16 = in_alloc_full[15] ? 16'h8000 : 16'h0; // @[Mux.scala 47:70]
  wire [15:0] _in_alloc_oh_T_17 = in_alloc_full[14] ? 16'h4000 : _in_alloc_oh_T_16; // @[Mux.scala 47:70]
  wire [15:0] _in_alloc_oh_T_18 = in_alloc_full[13] ? 16'h2000 : _in_alloc_oh_T_17; // @[Mux.scala 47:70]
  wire [15:0] _in_alloc_oh_T_19 = in_alloc_full[12] ? 16'h1000 : _in_alloc_oh_T_18; // @[Mux.scala 47:70]
  wire [15:0] _in_alloc_oh_T_20 = in_alloc_full[11] ? 16'h800 : _in_alloc_oh_T_19; // @[Mux.scala 47:70]
  wire [15:0] _in_alloc_oh_T_21 = in_alloc_full[10] ? 16'h400 : _in_alloc_oh_T_20; // @[Mux.scala 47:70]
  wire [15:0] _in_alloc_oh_T_22 = in_alloc_full[9] ? 16'h200 : _in_alloc_oh_T_21; // @[Mux.scala 47:70]
  wire [15:0] _in_alloc_oh_T_23 = in_alloc_full[8] ? 16'h100 : _in_alloc_oh_T_22; // @[Mux.scala 47:70]
  wire [15:0] _in_alloc_oh_T_24 = in_alloc_full[7] ? 16'h80 : _in_alloc_oh_T_23; // @[Mux.scala 47:70]
  wire [15:0] _in_alloc_oh_T_25 = in_alloc_full[6] ? 16'h40 : _in_alloc_oh_T_24; // @[Mux.scala 47:70]
  wire [15:0] _in_alloc_oh_T_26 = in_alloc_full[5] ? 16'h20 : _in_alloc_oh_T_25; // @[Mux.scala 47:70]
  wire [15:0] _in_alloc_oh_T_27 = in_alloc_full[4] ? 16'h10 : _in_alloc_oh_T_26; // @[Mux.scala 47:70]
  wire [15:0] _in_alloc_oh_T_28 = in_alloc_full[3] ? 16'h8 : _in_alloc_oh_T_27; // @[Mux.scala 47:70]
  wire [15:0] _in_alloc_oh_T_29 = in_alloc_full[2] ? 16'h4 : _in_alloc_oh_T_28; // @[Mux.scala 47:70]
  wire [15:0] _in_alloc_oh_T_30 = in_alloc_full[1] ? 16'h2 : _in_alloc_oh_T_29; // @[Mux.scala 47:70]
  wire [15:0] in_alloc_oh = in_alloc_full[0] ? 16'h1 : _in_alloc_oh_T_30; // @[Mux.scala 47:70]
  wire [7:0] in_alloc_sel = in_alloc_oh[7:0] | in_alloc_oh[15:8]; // @[ISLIP.scala 20:28]
  wire [7:0] _in_alloc_mask_T_16 = in_alloc_sel[7] ? 8'hff : 8'h0; // @[Mux.scala 101:16]
  wire [7:0] _in_alloc_mask_T_17 = in_alloc_sel[6] ? 8'h7f : _in_alloc_mask_T_16; // @[Mux.scala 101:16]
  wire [7:0] _in_alloc_mask_T_18 = in_alloc_sel[5] ? 8'h3f : _in_alloc_mask_T_17; // @[Mux.scala 101:16]
  wire [7:0] _in_alloc_mask_T_19 = in_alloc_sel[4] ? 8'h1f : _in_alloc_mask_T_18; // @[Mux.scala 101:16]
  wire [7:0] _in_alloc_mask_T_20 = in_alloc_sel[3] ? 8'hf : _in_alloc_mask_T_19; // @[Mux.scala 101:16]
  wire [7:0] _in_alloc_mask_T_21 = in_alloc_sel[2] ? 8'h7 : _in_alloc_mask_T_20; // @[Mux.scala 101:16]
  wire [7:0] _T = {io_resp_0_vc_sel_1_3,io_resp_0_vc_sel_1_2,io_resp_0_vc_sel_1_1,io_resp_0_vc_sel_1_0,
    io_resp_0_vc_sel_0_3,io_resp_0_vc_sel_0_2,io_resp_0_vc_sel_0_1,io_resp_0_vc_sel_0_0}; // @[SingleVCAllocator.scala 53:39]
  wire [1:0] _T_9 = _T[0] + _T[1]; // @[Bitwise.scala 51:90]
  wire [1:0] _T_11 = _T[2] + _T[3]; // @[Bitwise.scala 51:90]
  wire [2:0] _T_13 = _T_9 + _T_11; // @[Bitwise.scala 51:90]
  wire [1:0] _T_15 = _T[4] + _T[5]; // @[Bitwise.scala 51:90]
  wire [1:0] _T_17 = _T[6] + _T[7]; // @[Bitwise.scala 51:90]
  wire [2:0] _T_19 = _T_15 + _T_17; // @[Bitwise.scala 51:90]
  wire [3:0] _T_21 = _T_13 + _T_19; // @[Bitwise.scala 51:90]
  assign io_req_0_ready = in_arb_filter[0] | in_arb_filter[1]; // @[SingleVCAllocator.scala 20:57]
  assign io_resp_0_vc_sel_1_0 = in_arb_vals_0 & in_alloc_sel[4]; // @[SingleVCAllocator.scala 41:18]
  assign io_resp_0_vc_sel_1_1 = in_arb_vals_0 & in_alloc_sel[5]; // @[SingleVCAllocator.scala 41:18]
  assign io_resp_0_vc_sel_1_2 = in_arb_vals_0 & in_alloc_sel[6]; // @[SingleVCAllocator.scala 41:18]
  assign io_resp_0_vc_sel_1_3 = in_arb_vals_0 & in_alloc_sel[7]; // @[SingleVCAllocator.scala 41:18]
  assign io_resp_0_vc_sel_0_0 = in_arb_vals_0 & in_alloc_sel[0]; // @[SingleVCAllocator.scala 41:18]
  assign io_resp_0_vc_sel_0_1 = in_arb_vals_0 & in_alloc_sel[1]; // @[SingleVCAllocator.scala 41:18]
  assign io_resp_0_vc_sel_0_2 = in_arb_vals_0 & in_alloc_sel[2]; // @[SingleVCAllocator.scala 41:18]
  assign io_resp_0_vc_sel_0_3 = in_arb_vals_0 & in_alloc_sel[3]; // @[SingleVCAllocator.scala 41:18]
  assign io_out_allocs_1_1_alloc = in_arb_vals_0 & in_alloc_sel[5]; // @[SingleVCAllocator.scala 41:18]
  assign io_out_allocs_1_2_alloc = in_arb_vals_0 & in_alloc_sel[6]; // @[SingleVCAllocator.scala 41:18]
  assign io_out_allocs_1_3_alloc = in_arb_vals_0 & in_alloc_sel[7]; // @[SingleVCAllocator.scala 41:18]
  assign io_out_allocs_0_1_alloc = in_arb_vals_0 & in_alloc_sel[1]; // @[SingleVCAllocator.scala 41:18]
  assign io_out_allocs_0_2_alloc = in_arb_vals_0 & in_alloc_sel[2]; // @[SingleVCAllocator.scala 41:18]
  assign io_out_allocs_0_3_alloc = in_arb_vals_0 & in_alloc_sel[3]; // @[SingleVCAllocator.scala 41:18]
  always @(posedge clock) begin
    if (reset) begin // @[SingleVCAllocator.scala 16:21]
      mask <= 1'h0; // @[SingleVCAllocator.scala 16:21]
    end else begin
      mask <= _GEN_0;
    end
    if (reset) begin // @[ISLIP.scala 17:25]
      in_alloc_mask <= 8'h0; // @[ISLIP.scala 17:25]
    end else if (_in_alloc_T) begin // @[ISLIP.scala 21:19]
      if (in_alloc_sel[0]) begin // @[Mux.scala 101:16]
        in_alloc_mask <= 8'h1;
      end else if (in_alloc_sel[1]) begin // @[Mux.scala 101:16]
        in_alloc_mask <= 8'h3;
      end else begin
        in_alloc_mask <= _in_alloc_mask_T_21;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(_T_21 <= 4'h1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at SingleVCAllocator.scala:53 assert(PopCount(io.resp(i).vc_sel.asUInt) <= 1.U)\n"); // @[SingleVCAllocator.scala 53:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mask = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  in_alloc_mask = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(_T_21 <= 4'h1); // @[SingleVCAllocator.scala 53:11]
    end
  end
endmodule
module RouteComputer(
  input  [1:0] io_req_0_bits_flow_ingress_node,
  input  [1:0] io_req_0_bits_flow_egress_node,
  output       io_resp_0_vc_sel_1_0,
  output       io_resp_0_vc_sel_1_1,
  output       io_resp_0_vc_sel_1_2,
  output       io_resp_0_vc_sel_1_3,
  output       io_resp_0_vc_sel_0_0,
  output       io_resp_0_vc_sel_0_1,
  output       io_resp_0_vc_sel_0_2,
  output       io_resp_0_vc_sel_0_3
);
  wire [5:0] addr = {2'h0,io_req_0_bits_flow_ingress_node,io_req_0_bits_flow_egress_node}; // @[RouteComputer.scala 74:27]
  wire [5:0] decoded_invInputs = ~addr; // @[pla.scala 78:21]
  wire  decoded_andMatrixInput_0 = decoded_invInputs[1]; // @[pla.scala 91:29]
  wire  decoded_andMatrixInput_1 = decoded_invInputs[2]; // @[pla.scala 91:29]
  wire  decoded_andMatrixInput_2 = decoded_invInputs[3]; // @[pla.scala 91:29]
  wire  decoded_andMatrixInput_3 = decoded_invInputs[4]; // @[pla.scala 91:29]
  wire  decoded_andMatrixInput_4 = decoded_invInputs[5]; // @[pla.scala 91:29]
  wire [4:0] _decoded_T = {decoded_andMatrixInput_0,decoded_andMatrixInput_1,decoded_andMatrixInput_2,
    decoded_andMatrixInput_3,decoded_andMatrixInput_4}; // @[Cat.scala 33:92]
  wire  _decoded_T_1 = &_decoded_T; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_0_1 = addr[1]; // @[pla.scala 90:45]
  wire [4:0] _decoded_T_2 = {decoded_andMatrixInput_0_1,decoded_andMatrixInput_1,decoded_andMatrixInput_2,
    decoded_andMatrixInput_3,decoded_andMatrixInput_4}; // @[Cat.scala 33:92]
  wire  _decoded_T_3 = &_decoded_T_2; // @[pla.scala 98:74]
  wire  _decoded_orMatrixOutputs_T = |_decoded_T_3; // @[pla.scala 114:39]
  wire  _decoded_orMatrixOutputs_T_3 = |_decoded_T_1; // @[pla.scala 114:39]
  wire [7:0] decoded_orMatrixOutputs = {1'h0,_decoded_orMatrixOutputs_T_3,_decoded_orMatrixOutputs_T_3,
    _decoded_orMatrixOutputs_T_3,1'h0,_decoded_orMatrixOutputs_T,_decoded_orMatrixOutputs_T,_decoded_orMatrixOutputs_T}; // @[Cat.scala 33:92]
  wire [7:0] decoded_invMatrixOutputs = {decoded_orMatrixOutputs[7],decoded_orMatrixOutputs[6],decoded_orMatrixOutputs[5
    ],decoded_orMatrixOutputs[4],decoded_orMatrixOutputs[3],decoded_orMatrixOutputs[2],decoded_orMatrixOutputs[1],
    decoded_orMatrixOutputs[0]}; // @[Cat.scala 33:92]
  wire [7:0] _GEN_0 = {{4'd0}, decoded_invMatrixOutputs[7:4]}; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_7 = _GEN_0 & 8'hf; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_9 = {decoded_invMatrixOutputs[3:0], 4'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _decoded_T_11 = _decoded_T_9 & 8'hf0; // @[Bitwise.scala 108:80]
  wire [7:0] _decoded_T_12 = _decoded_T_7 | _decoded_T_11; // @[Bitwise.scala 108:39]
  wire [7:0] _GEN_1 = {{2'd0}, _decoded_T_12[7:2]}; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_17 = _GEN_1 & 8'h33; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_19 = {_decoded_T_12[5:0], 2'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _decoded_T_21 = _decoded_T_19 & 8'hcc; // @[Bitwise.scala 108:80]
  wire [7:0] _decoded_T_22 = _decoded_T_17 | _decoded_T_21; // @[Bitwise.scala 108:39]
  wire [7:0] _GEN_2 = {{1'd0}, _decoded_T_22[7:1]}; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_27 = _GEN_2 & 8'h55; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_29 = {_decoded_T_22[6:0], 1'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _decoded_T_31 = _decoded_T_29 & 8'haa; // @[Bitwise.scala 108:80]
  wire [7:0] decoded = _decoded_T_27 | _decoded_T_31; // @[Bitwise.scala 108:39]
  assign io_resp_0_vc_sel_1_0 = decoded[4]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_1_1 = decoded[5]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_1_2 = decoded[6]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_1_3 = decoded[7]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_0_0 = decoded[0]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_0_1 = decoded[1]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_0_2 = decoded[2]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_0_3 = decoded[3]; // @[RouteComputer.scala 90:46]
endmodule
module Router(
  input         clock,
  input         reset,
  output        auto_ingress_nodes_in_flit_ready,
  input         auto_ingress_nodes_in_flit_valid,
  input         auto_ingress_nodes_in_flit_bits_head,
  input         auto_ingress_nodes_in_flit_bits_tail,
  input  [63:0] auto_ingress_nodes_in_flit_bits_payload,
  input         auto_ingress_nodes_in_flit_bits_egress_id,
  output        auto_source_nodes_out_1_flit_0_valid,
  output        auto_source_nodes_out_1_flit_0_bits_head,
  output        auto_source_nodes_out_1_flit_0_bits_tail,
  output [63:0] auto_source_nodes_out_1_flit_0_bits_payload,
  output [1:0]  auto_source_nodes_out_1_flit_0_bits_flow_ingress_node,
  output [1:0]  auto_source_nodes_out_1_flit_0_bits_flow_egress_node,
  output [1:0]  auto_source_nodes_out_1_flit_0_bits_virt_channel_id,
  input  [3:0]  auto_source_nodes_out_1_credit_return,
  input  [3:0]  auto_source_nodes_out_1_vc_free,
  output        auto_source_nodes_out_0_flit_0_valid,
  output        auto_source_nodes_out_0_flit_0_bits_head,
  output        auto_source_nodes_out_0_flit_0_bits_tail,
  output [63:0] auto_source_nodes_out_0_flit_0_bits_payload,
  output [1:0]  auto_source_nodes_out_0_flit_0_bits_flow_ingress_node,
  output [1:0]  auto_source_nodes_out_0_flit_0_bits_flow_egress_node,
  output [1:0]  auto_source_nodes_out_0_flit_0_bits_virt_channel_id,
  input  [3:0]  auto_source_nodes_out_0_credit_return,
  input  [3:0]  auto_source_nodes_out_0_vc_free
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire  ingress_unit_0_from_0_clock; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_reset; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_router_req_valid; // @[Router.scala 116:13]
  wire [1:0] ingress_unit_0_from_0_io_router_req_bits_flow_ingress_node; // @[Router.scala 116:13]
  wire [1:0] ingress_unit_0_from_0_io_router_req_bits_flow_egress_node; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_router_resp_vc_sel_1_0; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_router_resp_vc_sel_1_1; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_router_resp_vc_sel_1_2; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_router_resp_vc_sel_1_3; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_router_resp_vc_sel_0_0; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_router_resp_vc_sel_0_1; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_router_resp_vc_sel_0_2; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_router_resp_vc_sel_0_3; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_vcalloc_req_ready; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_vcalloc_req_valid; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_vcalloc_req_bits_vc_sel_1_0; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_vcalloc_req_bits_vc_sel_1_1; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_vcalloc_req_bits_vc_sel_1_2; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_vcalloc_req_bits_vc_sel_1_3; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_0; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_1; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_2; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_3; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_vcalloc_resp_vc_sel_1_0; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_vcalloc_resp_vc_sel_1_1; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_vcalloc_resp_vc_sel_1_2; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_vcalloc_resp_vc_sel_1_3; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_vcalloc_resp_vc_sel_0_0; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_vcalloc_resp_vc_sel_0_1; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_vcalloc_resp_vc_sel_0_2; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_vcalloc_resp_vc_sel_0_3; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_out_credit_available_1_1; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_out_credit_available_1_2; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_out_credit_available_1_3; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_out_credit_available_0_1; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_out_credit_available_0_2; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_out_credit_available_0_3; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_salloc_req_0_ready; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_salloc_req_0_valid; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_salloc_req_0_bits_vc_sel_1_0; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_salloc_req_0_bits_vc_sel_1_1; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_salloc_req_0_bits_vc_sel_1_2; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_salloc_req_0_bits_vc_sel_1_3; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_0; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_1; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_2; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_3; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_salloc_req_0_bits_tail; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_out_0_valid; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_out_0_bits_flit_head; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_out_0_bits_flit_tail; // @[Router.scala 116:13]
  wire [63:0] ingress_unit_0_from_0_io_out_0_bits_flit_payload; // @[Router.scala 116:13]
  wire [1:0] ingress_unit_0_from_0_io_out_0_bits_flit_flow_ingress_node; // @[Router.scala 116:13]
  wire [1:0] ingress_unit_0_from_0_io_out_0_bits_flit_flow_egress_node; // @[Router.scala 116:13]
  wire [1:0] ingress_unit_0_from_0_io_out_0_bits_out_virt_channel; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_in_ready; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_in_valid; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_in_bits_head; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_in_bits_tail; // @[Router.scala 116:13]
  wire [63:0] ingress_unit_0_from_0_io_in_bits_payload; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_0_io_in_bits_egress_id; // @[Router.scala 116:13]
  wire  output_unit_0_to_1_clock; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_reset; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_in_0_valid; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_in_0_bits_head; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_in_0_bits_tail; // @[Router.scala 122:13]
  wire [63:0] output_unit_0_to_1_io_in_0_bits_payload; // @[Router.scala 122:13]
  wire [1:0] output_unit_0_to_1_io_in_0_bits_flow_ingress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_0_to_1_io_in_0_bits_flow_egress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_0_to_1_io_in_0_bits_virt_channel_id; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_credit_available_1; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_credit_available_2; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_credit_available_3; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_channel_status_1_occupied; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_channel_status_2_occupied; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_channel_status_3_occupied; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_allocs_1_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_allocs_2_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_allocs_3_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_credit_alloc_1_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_credit_alloc_2_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_credit_alloc_3_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_out_flit_0_valid; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_out_flit_0_bits_head; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_out_flit_0_bits_tail; // @[Router.scala 122:13]
  wire [63:0] output_unit_0_to_1_io_out_flit_0_bits_payload; // @[Router.scala 122:13]
  wire [1:0] output_unit_0_to_1_io_out_flit_0_bits_flow_ingress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_0_to_1_io_out_flit_0_bits_flow_egress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_0_to_1_io_out_flit_0_bits_virt_channel_id; // @[Router.scala 122:13]
  wire [3:0] output_unit_0_to_1_io_out_credit_return; // @[Router.scala 122:13]
  wire [3:0] output_unit_0_to_1_io_out_vc_free; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_clock; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_reset; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_in_0_valid; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_in_0_bits_head; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_in_0_bits_tail; // @[Router.scala 122:13]
  wire [63:0] output_unit_1_to_3_io_in_0_bits_payload; // @[Router.scala 122:13]
  wire [1:0] output_unit_1_to_3_io_in_0_bits_flow_ingress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_1_to_3_io_in_0_bits_flow_egress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_1_to_3_io_in_0_bits_virt_channel_id; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_credit_available_1; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_credit_available_2; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_credit_available_3; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_channel_status_1_occupied; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_channel_status_2_occupied; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_channel_status_3_occupied; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_allocs_1_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_allocs_2_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_allocs_3_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_credit_alloc_1_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_credit_alloc_2_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_credit_alloc_3_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_out_flit_0_valid; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_out_flit_0_bits_head; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_out_flit_0_bits_tail; // @[Router.scala 122:13]
  wire [63:0] output_unit_1_to_3_io_out_flit_0_bits_payload; // @[Router.scala 122:13]
  wire [1:0] output_unit_1_to_3_io_out_flit_0_bits_flow_ingress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_1_to_3_io_out_flit_0_bits_flow_egress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_1_to_3_io_out_flit_0_bits_virt_channel_id; // @[Router.scala 122:13]
  wire [3:0] output_unit_1_to_3_io_out_credit_return; // @[Router.scala 122:13]
  wire [3:0] output_unit_1_to_3_io_out_vc_free; // @[Router.scala 122:13]
  wire  switch_clock; // @[Router.scala 129:24]
  wire  switch_reset; // @[Router.scala 129:24]
  wire  switch_io_in_0_0_valid; // @[Router.scala 129:24]
  wire  switch_io_in_0_0_bits_flit_head; // @[Router.scala 129:24]
  wire  switch_io_in_0_0_bits_flit_tail; // @[Router.scala 129:24]
  wire [63:0] switch_io_in_0_0_bits_flit_payload; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_0_0_bits_flit_flow_ingress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_0_0_bits_flit_flow_egress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_0_0_bits_out_virt_channel; // @[Router.scala 129:24]
  wire  switch_io_out_1_0_valid; // @[Router.scala 129:24]
  wire  switch_io_out_1_0_bits_head; // @[Router.scala 129:24]
  wire  switch_io_out_1_0_bits_tail; // @[Router.scala 129:24]
  wire [63:0] switch_io_out_1_0_bits_payload; // @[Router.scala 129:24]
  wire [1:0] switch_io_out_1_0_bits_flow_ingress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_out_1_0_bits_flow_egress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_out_1_0_bits_virt_channel_id; // @[Router.scala 129:24]
  wire  switch_io_out_0_0_valid; // @[Router.scala 129:24]
  wire  switch_io_out_0_0_bits_head; // @[Router.scala 129:24]
  wire  switch_io_out_0_0_bits_tail; // @[Router.scala 129:24]
  wire [63:0] switch_io_out_0_0_bits_payload; // @[Router.scala 129:24]
  wire [1:0] switch_io_out_0_0_bits_flow_ingress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_out_0_0_bits_flow_egress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_out_0_0_bits_virt_channel_id; // @[Router.scala 129:24]
  wire  switch_io_sel_1_0_0_0; // @[Router.scala 129:24]
  wire  switch_io_sel_0_0_0_0; // @[Router.scala 129:24]
  wire  switch_allocator_clock; // @[Router.scala 130:34]
  wire  switch_allocator_reset; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_ready; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_valid; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_1_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_1_1; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_1_2; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_1_3; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_0_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_0_1; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_0_2; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_0_3; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_tail; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_1_1_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_1_2_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_1_3_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_0_1_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_0_2_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_0_3_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_1_0_0_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_0_0_0_0; // @[Router.scala 130:34]
  wire  vc_allocator_clock; // @[Router.scala 131:30]
  wire  vc_allocator_reset; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_ready; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_valid; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_1_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_1_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_1_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_1_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_0_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_0_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_0_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_0_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_1_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_1_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_1_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_1_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_0_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_0_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_0_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_0_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_1_1_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_1_2_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_1_3_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_0_1_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_0_2_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_0_3_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_1_1_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_1_2_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_1_3_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_0_1_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_0_2_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_0_3_alloc; // @[Router.scala 131:30]
  wire [1:0] route_computer_io_req_0_bits_flow_ingress_node; // @[Router.scala 134:32]
  wire [1:0] route_computer_io_req_0_bits_flow_egress_node; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_1_0; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_1_1; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_1_2; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_1_3; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_0_0; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_0_1; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_0_2; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_0_3; // @[Router.scala 134:32]
  wire [19:0] plusarg_reader_out; // @[PlusArg.scala 80:11]
  reg  switch_io_sel_REG_1_0_0_0; // @[Router.scala 176:14]
  reg  switch_io_sel_REG_0_0_0_0; // @[Router.scala 176:14]
  reg [63:0] debug_tsc; // @[Router.scala 193:28]
  wire [63:0] _debug_tsc_T_1 = debug_tsc + 64'h1; // @[Router.scala 194:28]
  reg [63:0] debug_sample; // @[Router.scala 195:31]
  wire [63:0] _debug_sample_T_1 = debug_sample + 64'h1; // @[Router.scala 196:34]
  wire [19:0] _T_1 = plusarg_reader_out - 20'h1; // @[Router.scala 198:40]
  wire [63:0] _GEN_2 = {{44'd0}, _T_1}; // @[Router.scala 198:24]
  wire  _T_2 = debug_sample == _GEN_2; // @[Router.scala 198:24]
  wire  bundleIn_0_flit_ready = ingress_unit_0_from_0_io_in_ready; // @[Nodes.scala 1215:84 Router.scala 142:68]
  wire  _T_3 = bundleIn_0_flit_ready & auto_ingress_nodes_in_flit_valid; // @[Decoupled.scala 51:35]
  reg [63:0] util_ctr; // @[Router.scala 201:29]
  reg  fired; // @[Router.scala 202:26]
  wire [63:0] _GEN_3 = {{63'd0}, _T_3}; // @[Router.scala 203:28]
  wire [63:0] _util_ctr_T_1 = util_ctr + _GEN_3; // @[Router.scala 203:28]
  wire  _T_9 = plusarg_reader_out != 20'h0 & _T_2 & fired; // @[Router.scala 205:71]
  wire  fires_count = vc_allocator_io_req_0_ready & vc_allocator_io_req_0_valid; // @[Decoupled.scala 51:35]
  IngressUnit ingress_unit_0_from_0 ( // @[Router.scala 116:13]
    .clock(ingress_unit_0_from_0_clock),
    .reset(ingress_unit_0_from_0_reset),
    .io_router_req_valid(ingress_unit_0_from_0_io_router_req_valid),
    .io_router_req_bits_flow_ingress_node(ingress_unit_0_from_0_io_router_req_bits_flow_ingress_node),
    .io_router_req_bits_flow_egress_node(ingress_unit_0_from_0_io_router_req_bits_flow_egress_node),
    .io_router_resp_vc_sel_1_0(ingress_unit_0_from_0_io_router_resp_vc_sel_1_0),
    .io_router_resp_vc_sel_1_1(ingress_unit_0_from_0_io_router_resp_vc_sel_1_1),
    .io_router_resp_vc_sel_1_2(ingress_unit_0_from_0_io_router_resp_vc_sel_1_2),
    .io_router_resp_vc_sel_1_3(ingress_unit_0_from_0_io_router_resp_vc_sel_1_3),
    .io_router_resp_vc_sel_0_0(ingress_unit_0_from_0_io_router_resp_vc_sel_0_0),
    .io_router_resp_vc_sel_0_1(ingress_unit_0_from_0_io_router_resp_vc_sel_0_1),
    .io_router_resp_vc_sel_0_2(ingress_unit_0_from_0_io_router_resp_vc_sel_0_2),
    .io_router_resp_vc_sel_0_3(ingress_unit_0_from_0_io_router_resp_vc_sel_0_3),
    .io_vcalloc_req_ready(ingress_unit_0_from_0_io_vcalloc_req_ready),
    .io_vcalloc_req_valid(ingress_unit_0_from_0_io_vcalloc_req_valid),
    .io_vcalloc_req_bits_vc_sel_1_0(ingress_unit_0_from_0_io_vcalloc_req_bits_vc_sel_1_0),
    .io_vcalloc_req_bits_vc_sel_1_1(ingress_unit_0_from_0_io_vcalloc_req_bits_vc_sel_1_1),
    .io_vcalloc_req_bits_vc_sel_1_2(ingress_unit_0_from_0_io_vcalloc_req_bits_vc_sel_1_2),
    .io_vcalloc_req_bits_vc_sel_1_3(ingress_unit_0_from_0_io_vcalloc_req_bits_vc_sel_1_3),
    .io_vcalloc_req_bits_vc_sel_0_0(ingress_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_0),
    .io_vcalloc_req_bits_vc_sel_0_1(ingress_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_1),
    .io_vcalloc_req_bits_vc_sel_0_2(ingress_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_2),
    .io_vcalloc_req_bits_vc_sel_0_3(ingress_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_3),
    .io_vcalloc_resp_vc_sel_1_0(ingress_unit_0_from_0_io_vcalloc_resp_vc_sel_1_0),
    .io_vcalloc_resp_vc_sel_1_1(ingress_unit_0_from_0_io_vcalloc_resp_vc_sel_1_1),
    .io_vcalloc_resp_vc_sel_1_2(ingress_unit_0_from_0_io_vcalloc_resp_vc_sel_1_2),
    .io_vcalloc_resp_vc_sel_1_3(ingress_unit_0_from_0_io_vcalloc_resp_vc_sel_1_3),
    .io_vcalloc_resp_vc_sel_0_0(ingress_unit_0_from_0_io_vcalloc_resp_vc_sel_0_0),
    .io_vcalloc_resp_vc_sel_0_1(ingress_unit_0_from_0_io_vcalloc_resp_vc_sel_0_1),
    .io_vcalloc_resp_vc_sel_0_2(ingress_unit_0_from_0_io_vcalloc_resp_vc_sel_0_2),
    .io_vcalloc_resp_vc_sel_0_3(ingress_unit_0_from_0_io_vcalloc_resp_vc_sel_0_3),
    .io_out_credit_available_1_1(ingress_unit_0_from_0_io_out_credit_available_1_1),
    .io_out_credit_available_1_2(ingress_unit_0_from_0_io_out_credit_available_1_2),
    .io_out_credit_available_1_3(ingress_unit_0_from_0_io_out_credit_available_1_3),
    .io_out_credit_available_0_1(ingress_unit_0_from_0_io_out_credit_available_0_1),
    .io_out_credit_available_0_2(ingress_unit_0_from_0_io_out_credit_available_0_2),
    .io_out_credit_available_0_3(ingress_unit_0_from_0_io_out_credit_available_0_3),
    .io_salloc_req_0_ready(ingress_unit_0_from_0_io_salloc_req_0_ready),
    .io_salloc_req_0_valid(ingress_unit_0_from_0_io_salloc_req_0_valid),
    .io_salloc_req_0_bits_vc_sel_1_0(ingress_unit_0_from_0_io_salloc_req_0_bits_vc_sel_1_0),
    .io_salloc_req_0_bits_vc_sel_1_1(ingress_unit_0_from_0_io_salloc_req_0_bits_vc_sel_1_1),
    .io_salloc_req_0_bits_vc_sel_1_2(ingress_unit_0_from_0_io_salloc_req_0_bits_vc_sel_1_2),
    .io_salloc_req_0_bits_vc_sel_1_3(ingress_unit_0_from_0_io_salloc_req_0_bits_vc_sel_1_3),
    .io_salloc_req_0_bits_vc_sel_0_0(ingress_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_0),
    .io_salloc_req_0_bits_vc_sel_0_1(ingress_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_1),
    .io_salloc_req_0_bits_vc_sel_0_2(ingress_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_2),
    .io_salloc_req_0_bits_vc_sel_0_3(ingress_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_3),
    .io_salloc_req_0_bits_tail(ingress_unit_0_from_0_io_salloc_req_0_bits_tail),
    .io_out_0_valid(ingress_unit_0_from_0_io_out_0_valid),
    .io_out_0_bits_flit_head(ingress_unit_0_from_0_io_out_0_bits_flit_head),
    .io_out_0_bits_flit_tail(ingress_unit_0_from_0_io_out_0_bits_flit_tail),
    .io_out_0_bits_flit_payload(ingress_unit_0_from_0_io_out_0_bits_flit_payload),
    .io_out_0_bits_flit_flow_ingress_node(ingress_unit_0_from_0_io_out_0_bits_flit_flow_ingress_node),
    .io_out_0_bits_flit_flow_egress_node(ingress_unit_0_from_0_io_out_0_bits_flit_flow_egress_node),
    .io_out_0_bits_out_virt_channel(ingress_unit_0_from_0_io_out_0_bits_out_virt_channel),
    .io_in_ready(ingress_unit_0_from_0_io_in_ready),
    .io_in_valid(ingress_unit_0_from_0_io_in_valid),
    .io_in_bits_head(ingress_unit_0_from_0_io_in_bits_head),
    .io_in_bits_tail(ingress_unit_0_from_0_io_in_bits_tail),
    .io_in_bits_payload(ingress_unit_0_from_0_io_in_bits_payload),
    .io_in_bits_egress_id(ingress_unit_0_from_0_io_in_bits_egress_id)
  );
  OutputUnit output_unit_0_to_1 ( // @[Router.scala 122:13]
    .clock(output_unit_0_to_1_clock),
    .reset(output_unit_0_to_1_reset),
    .io_in_0_valid(output_unit_0_to_1_io_in_0_valid),
    .io_in_0_bits_head(output_unit_0_to_1_io_in_0_bits_head),
    .io_in_0_bits_tail(output_unit_0_to_1_io_in_0_bits_tail),
    .io_in_0_bits_payload(output_unit_0_to_1_io_in_0_bits_payload),
    .io_in_0_bits_flow_ingress_node(output_unit_0_to_1_io_in_0_bits_flow_ingress_node),
    .io_in_0_bits_flow_egress_node(output_unit_0_to_1_io_in_0_bits_flow_egress_node),
    .io_in_0_bits_virt_channel_id(output_unit_0_to_1_io_in_0_bits_virt_channel_id),
    .io_credit_available_1(output_unit_0_to_1_io_credit_available_1),
    .io_credit_available_2(output_unit_0_to_1_io_credit_available_2),
    .io_credit_available_3(output_unit_0_to_1_io_credit_available_3),
    .io_channel_status_1_occupied(output_unit_0_to_1_io_channel_status_1_occupied),
    .io_channel_status_2_occupied(output_unit_0_to_1_io_channel_status_2_occupied),
    .io_channel_status_3_occupied(output_unit_0_to_1_io_channel_status_3_occupied),
    .io_allocs_1_alloc(output_unit_0_to_1_io_allocs_1_alloc),
    .io_allocs_2_alloc(output_unit_0_to_1_io_allocs_2_alloc),
    .io_allocs_3_alloc(output_unit_0_to_1_io_allocs_3_alloc),
    .io_credit_alloc_1_alloc(output_unit_0_to_1_io_credit_alloc_1_alloc),
    .io_credit_alloc_2_alloc(output_unit_0_to_1_io_credit_alloc_2_alloc),
    .io_credit_alloc_3_alloc(output_unit_0_to_1_io_credit_alloc_3_alloc),
    .io_out_flit_0_valid(output_unit_0_to_1_io_out_flit_0_valid),
    .io_out_flit_0_bits_head(output_unit_0_to_1_io_out_flit_0_bits_head),
    .io_out_flit_0_bits_tail(output_unit_0_to_1_io_out_flit_0_bits_tail),
    .io_out_flit_0_bits_payload(output_unit_0_to_1_io_out_flit_0_bits_payload),
    .io_out_flit_0_bits_flow_ingress_node(output_unit_0_to_1_io_out_flit_0_bits_flow_ingress_node),
    .io_out_flit_0_bits_flow_egress_node(output_unit_0_to_1_io_out_flit_0_bits_flow_egress_node),
    .io_out_flit_0_bits_virt_channel_id(output_unit_0_to_1_io_out_flit_0_bits_virt_channel_id),
    .io_out_credit_return(output_unit_0_to_1_io_out_credit_return),
    .io_out_vc_free(output_unit_0_to_1_io_out_vc_free)
  );
  OutputUnit output_unit_1_to_3 ( // @[Router.scala 122:13]
    .clock(output_unit_1_to_3_clock),
    .reset(output_unit_1_to_3_reset),
    .io_in_0_valid(output_unit_1_to_3_io_in_0_valid),
    .io_in_0_bits_head(output_unit_1_to_3_io_in_0_bits_head),
    .io_in_0_bits_tail(output_unit_1_to_3_io_in_0_bits_tail),
    .io_in_0_bits_payload(output_unit_1_to_3_io_in_0_bits_payload),
    .io_in_0_bits_flow_ingress_node(output_unit_1_to_3_io_in_0_bits_flow_ingress_node),
    .io_in_0_bits_flow_egress_node(output_unit_1_to_3_io_in_0_bits_flow_egress_node),
    .io_in_0_bits_virt_channel_id(output_unit_1_to_3_io_in_0_bits_virt_channel_id),
    .io_credit_available_1(output_unit_1_to_3_io_credit_available_1),
    .io_credit_available_2(output_unit_1_to_3_io_credit_available_2),
    .io_credit_available_3(output_unit_1_to_3_io_credit_available_3),
    .io_channel_status_1_occupied(output_unit_1_to_3_io_channel_status_1_occupied),
    .io_channel_status_2_occupied(output_unit_1_to_3_io_channel_status_2_occupied),
    .io_channel_status_3_occupied(output_unit_1_to_3_io_channel_status_3_occupied),
    .io_allocs_1_alloc(output_unit_1_to_3_io_allocs_1_alloc),
    .io_allocs_2_alloc(output_unit_1_to_3_io_allocs_2_alloc),
    .io_allocs_3_alloc(output_unit_1_to_3_io_allocs_3_alloc),
    .io_credit_alloc_1_alloc(output_unit_1_to_3_io_credit_alloc_1_alloc),
    .io_credit_alloc_2_alloc(output_unit_1_to_3_io_credit_alloc_2_alloc),
    .io_credit_alloc_3_alloc(output_unit_1_to_3_io_credit_alloc_3_alloc),
    .io_out_flit_0_valid(output_unit_1_to_3_io_out_flit_0_valid),
    .io_out_flit_0_bits_head(output_unit_1_to_3_io_out_flit_0_bits_head),
    .io_out_flit_0_bits_tail(output_unit_1_to_3_io_out_flit_0_bits_tail),
    .io_out_flit_0_bits_payload(output_unit_1_to_3_io_out_flit_0_bits_payload),
    .io_out_flit_0_bits_flow_ingress_node(output_unit_1_to_3_io_out_flit_0_bits_flow_ingress_node),
    .io_out_flit_0_bits_flow_egress_node(output_unit_1_to_3_io_out_flit_0_bits_flow_egress_node),
    .io_out_flit_0_bits_virt_channel_id(output_unit_1_to_3_io_out_flit_0_bits_virt_channel_id),
    .io_out_credit_return(output_unit_1_to_3_io_out_credit_return),
    .io_out_vc_free(output_unit_1_to_3_io_out_vc_free)
  );
  Switch switch ( // @[Router.scala 129:24]
    .clock(switch_clock),
    .reset(switch_reset),
    .io_in_0_0_valid(switch_io_in_0_0_valid),
    .io_in_0_0_bits_flit_head(switch_io_in_0_0_bits_flit_head),
    .io_in_0_0_bits_flit_tail(switch_io_in_0_0_bits_flit_tail),
    .io_in_0_0_bits_flit_payload(switch_io_in_0_0_bits_flit_payload),
    .io_in_0_0_bits_flit_flow_ingress_node(switch_io_in_0_0_bits_flit_flow_ingress_node),
    .io_in_0_0_bits_flit_flow_egress_node(switch_io_in_0_0_bits_flit_flow_egress_node),
    .io_in_0_0_bits_out_virt_channel(switch_io_in_0_0_bits_out_virt_channel),
    .io_out_1_0_valid(switch_io_out_1_0_valid),
    .io_out_1_0_bits_head(switch_io_out_1_0_bits_head),
    .io_out_1_0_bits_tail(switch_io_out_1_0_bits_tail),
    .io_out_1_0_bits_payload(switch_io_out_1_0_bits_payload),
    .io_out_1_0_bits_flow_ingress_node(switch_io_out_1_0_bits_flow_ingress_node),
    .io_out_1_0_bits_flow_egress_node(switch_io_out_1_0_bits_flow_egress_node),
    .io_out_1_0_bits_virt_channel_id(switch_io_out_1_0_bits_virt_channel_id),
    .io_out_0_0_valid(switch_io_out_0_0_valid),
    .io_out_0_0_bits_head(switch_io_out_0_0_bits_head),
    .io_out_0_0_bits_tail(switch_io_out_0_0_bits_tail),
    .io_out_0_0_bits_payload(switch_io_out_0_0_bits_payload),
    .io_out_0_0_bits_flow_ingress_node(switch_io_out_0_0_bits_flow_ingress_node),
    .io_out_0_0_bits_flow_egress_node(switch_io_out_0_0_bits_flow_egress_node),
    .io_out_0_0_bits_virt_channel_id(switch_io_out_0_0_bits_virt_channel_id),
    .io_sel_1_0_0_0(switch_io_sel_1_0_0_0),
    .io_sel_0_0_0_0(switch_io_sel_0_0_0_0)
  );
  SwitchAllocator switch_allocator ( // @[Router.scala 130:34]
    .clock(switch_allocator_clock),
    .reset(switch_allocator_reset),
    .io_req_0_0_ready(switch_allocator_io_req_0_0_ready),
    .io_req_0_0_valid(switch_allocator_io_req_0_0_valid),
    .io_req_0_0_bits_vc_sel_1_0(switch_allocator_io_req_0_0_bits_vc_sel_1_0),
    .io_req_0_0_bits_vc_sel_1_1(switch_allocator_io_req_0_0_bits_vc_sel_1_1),
    .io_req_0_0_bits_vc_sel_1_2(switch_allocator_io_req_0_0_bits_vc_sel_1_2),
    .io_req_0_0_bits_vc_sel_1_3(switch_allocator_io_req_0_0_bits_vc_sel_1_3),
    .io_req_0_0_bits_vc_sel_0_0(switch_allocator_io_req_0_0_bits_vc_sel_0_0),
    .io_req_0_0_bits_vc_sel_0_1(switch_allocator_io_req_0_0_bits_vc_sel_0_1),
    .io_req_0_0_bits_vc_sel_0_2(switch_allocator_io_req_0_0_bits_vc_sel_0_2),
    .io_req_0_0_bits_vc_sel_0_3(switch_allocator_io_req_0_0_bits_vc_sel_0_3),
    .io_req_0_0_bits_tail(switch_allocator_io_req_0_0_bits_tail),
    .io_credit_alloc_1_1_alloc(switch_allocator_io_credit_alloc_1_1_alloc),
    .io_credit_alloc_1_2_alloc(switch_allocator_io_credit_alloc_1_2_alloc),
    .io_credit_alloc_1_3_alloc(switch_allocator_io_credit_alloc_1_3_alloc),
    .io_credit_alloc_0_1_alloc(switch_allocator_io_credit_alloc_0_1_alloc),
    .io_credit_alloc_0_2_alloc(switch_allocator_io_credit_alloc_0_2_alloc),
    .io_credit_alloc_0_3_alloc(switch_allocator_io_credit_alloc_0_3_alloc),
    .io_switch_sel_1_0_0_0(switch_allocator_io_switch_sel_1_0_0_0),
    .io_switch_sel_0_0_0_0(switch_allocator_io_switch_sel_0_0_0_0)
  );
  RotatingSingleVCAllocator vc_allocator ( // @[Router.scala 131:30]
    .clock(vc_allocator_clock),
    .reset(vc_allocator_reset),
    .io_req_0_ready(vc_allocator_io_req_0_ready),
    .io_req_0_valid(vc_allocator_io_req_0_valid),
    .io_req_0_bits_vc_sel_1_0(vc_allocator_io_req_0_bits_vc_sel_1_0),
    .io_req_0_bits_vc_sel_1_1(vc_allocator_io_req_0_bits_vc_sel_1_1),
    .io_req_0_bits_vc_sel_1_2(vc_allocator_io_req_0_bits_vc_sel_1_2),
    .io_req_0_bits_vc_sel_1_3(vc_allocator_io_req_0_bits_vc_sel_1_3),
    .io_req_0_bits_vc_sel_0_0(vc_allocator_io_req_0_bits_vc_sel_0_0),
    .io_req_0_bits_vc_sel_0_1(vc_allocator_io_req_0_bits_vc_sel_0_1),
    .io_req_0_bits_vc_sel_0_2(vc_allocator_io_req_0_bits_vc_sel_0_2),
    .io_req_0_bits_vc_sel_0_3(vc_allocator_io_req_0_bits_vc_sel_0_3),
    .io_resp_0_vc_sel_1_0(vc_allocator_io_resp_0_vc_sel_1_0),
    .io_resp_0_vc_sel_1_1(vc_allocator_io_resp_0_vc_sel_1_1),
    .io_resp_0_vc_sel_1_2(vc_allocator_io_resp_0_vc_sel_1_2),
    .io_resp_0_vc_sel_1_3(vc_allocator_io_resp_0_vc_sel_1_3),
    .io_resp_0_vc_sel_0_0(vc_allocator_io_resp_0_vc_sel_0_0),
    .io_resp_0_vc_sel_0_1(vc_allocator_io_resp_0_vc_sel_0_1),
    .io_resp_0_vc_sel_0_2(vc_allocator_io_resp_0_vc_sel_0_2),
    .io_resp_0_vc_sel_0_3(vc_allocator_io_resp_0_vc_sel_0_3),
    .io_channel_status_1_1_occupied(vc_allocator_io_channel_status_1_1_occupied),
    .io_channel_status_1_2_occupied(vc_allocator_io_channel_status_1_2_occupied),
    .io_channel_status_1_3_occupied(vc_allocator_io_channel_status_1_3_occupied),
    .io_channel_status_0_1_occupied(vc_allocator_io_channel_status_0_1_occupied),
    .io_channel_status_0_2_occupied(vc_allocator_io_channel_status_0_2_occupied),
    .io_channel_status_0_3_occupied(vc_allocator_io_channel_status_0_3_occupied),
    .io_out_allocs_1_1_alloc(vc_allocator_io_out_allocs_1_1_alloc),
    .io_out_allocs_1_2_alloc(vc_allocator_io_out_allocs_1_2_alloc),
    .io_out_allocs_1_3_alloc(vc_allocator_io_out_allocs_1_3_alloc),
    .io_out_allocs_0_1_alloc(vc_allocator_io_out_allocs_0_1_alloc),
    .io_out_allocs_0_2_alloc(vc_allocator_io_out_allocs_0_2_alloc),
    .io_out_allocs_0_3_alloc(vc_allocator_io_out_allocs_0_3_alloc)
  );
  RouteComputer route_computer ( // @[Router.scala 134:32]
    .io_req_0_bits_flow_ingress_node(route_computer_io_req_0_bits_flow_ingress_node),
    .io_req_0_bits_flow_egress_node(route_computer_io_req_0_bits_flow_egress_node),
    .io_resp_0_vc_sel_1_0(route_computer_io_resp_0_vc_sel_1_0),
    .io_resp_0_vc_sel_1_1(route_computer_io_resp_0_vc_sel_1_1),
    .io_resp_0_vc_sel_1_2(route_computer_io_resp_0_vc_sel_1_2),
    .io_resp_0_vc_sel_1_3(route_computer_io_resp_0_vc_sel_1_3),
    .io_resp_0_vc_sel_0_0(route_computer_io_resp_0_vc_sel_0_0),
    .io_resp_0_vc_sel_0_1(route_computer_io_resp_0_vc_sel_0_1),
    .io_resp_0_vc_sel_0_2(route_computer_io_resp_0_vc_sel_0_2),
    .io_resp_0_vc_sel_0_3(route_computer_io_resp_0_vc_sel_0_3)
  );
  plusarg_reader #(.FORMAT("noc_util_sample_rate=%d"), .DEFAULT(0), .WIDTH(20)) plusarg_reader ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_out)
  );
  assign auto_ingress_nodes_in_flit_ready = ingress_unit_0_from_0_io_in_ready; // @[Nodes.scala 1215:84 Router.scala 142:68]
  assign auto_source_nodes_out_1_flit_0_valid = output_unit_1_to_3_io_out_flit_0_valid; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_1_flit_0_bits_head = output_unit_1_to_3_io_out_flit_0_bits_head; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_1_flit_0_bits_tail = output_unit_1_to_3_io_out_flit_0_bits_tail; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_1_flit_0_bits_payload = output_unit_1_to_3_io_out_flit_0_bits_payload; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_1_flit_0_bits_flow_ingress_node = output_unit_1_to_3_io_out_flit_0_bits_flow_ingress_node
    ; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_1_flit_0_bits_flow_egress_node = output_unit_1_to_3_io_out_flit_0_bits_flow_egress_node; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_1_flit_0_bits_virt_channel_id = output_unit_1_to_3_io_out_flit_0_bits_virt_channel_id; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_0_flit_0_valid = output_unit_0_to_1_io_out_flit_0_valid; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_0_flit_0_bits_head = output_unit_0_to_1_io_out_flit_0_bits_head; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_0_flit_0_bits_tail = output_unit_0_to_1_io_out_flit_0_bits_tail; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_0_flit_0_bits_payload = output_unit_0_to_1_io_out_flit_0_bits_payload; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_0_flit_0_bits_flow_ingress_node = output_unit_0_to_1_io_out_flit_0_bits_flow_ingress_node
    ; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_0_flit_0_bits_flow_egress_node = output_unit_0_to_1_io_out_flit_0_bits_flow_egress_node; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_0_flit_0_bits_virt_channel_id = output_unit_0_to_1_io_out_flit_0_bits_virt_channel_id; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign ingress_unit_0_from_0_clock = clock;
  assign ingress_unit_0_from_0_reset = reset;
  assign ingress_unit_0_from_0_io_router_resp_vc_sel_1_0 = route_computer_io_resp_0_vc_sel_1_0; // @[Router.scala 148:38]
  assign ingress_unit_0_from_0_io_router_resp_vc_sel_1_1 = route_computer_io_resp_0_vc_sel_1_1; // @[Router.scala 148:38]
  assign ingress_unit_0_from_0_io_router_resp_vc_sel_1_2 = route_computer_io_resp_0_vc_sel_1_2; // @[Router.scala 148:38]
  assign ingress_unit_0_from_0_io_router_resp_vc_sel_1_3 = route_computer_io_resp_0_vc_sel_1_3; // @[Router.scala 148:38]
  assign ingress_unit_0_from_0_io_router_resp_vc_sel_0_0 = route_computer_io_resp_0_vc_sel_0_0; // @[Router.scala 148:38]
  assign ingress_unit_0_from_0_io_router_resp_vc_sel_0_1 = route_computer_io_resp_0_vc_sel_0_1; // @[Router.scala 148:38]
  assign ingress_unit_0_from_0_io_router_resp_vc_sel_0_2 = route_computer_io_resp_0_vc_sel_0_2; // @[Router.scala 148:38]
  assign ingress_unit_0_from_0_io_router_resp_vc_sel_0_3 = route_computer_io_resp_0_vc_sel_0_3; // @[Router.scala 148:38]
  assign ingress_unit_0_from_0_io_vcalloc_req_ready = vc_allocator_io_req_0_ready; // @[Router.scala 151:23]
  assign ingress_unit_0_from_0_io_vcalloc_resp_vc_sel_1_0 = vc_allocator_io_resp_0_vc_sel_1_0; // @[Router.scala 153:39]
  assign ingress_unit_0_from_0_io_vcalloc_resp_vc_sel_1_1 = vc_allocator_io_resp_0_vc_sel_1_1; // @[Router.scala 153:39]
  assign ingress_unit_0_from_0_io_vcalloc_resp_vc_sel_1_2 = vc_allocator_io_resp_0_vc_sel_1_2; // @[Router.scala 153:39]
  assign ingress_unit_0_from_0_io_vcalloc_resp_vc_sel_1_3 = vc_allocator_io_resp_0_vc_sel_1_3; // @[Router.scala 153:39]
  assign ingress_unit_0_from_0_io_vcalloc_resp_vc_sel_0_0 = vc_allocator_io_resp_0_vc_sel_0_0; // @[Router.scala 153:39]
  assign ingress_unit_0_from_0_io_vcalloc_resp_vc_sel_0_1 = vc_allocator_io_resp_0_vc_sel_0_1; // @[Router.scala 153:39]
  assign ingress_unit_0_from_0_io_vcalloc_resp_vc_sel_0_2 = vc_allocator_io_resp_0_vc_sel_0_2; // @[Router.scala 153:39]
  assign ingress_unit_0_from_0_io_vcalloc_resp_vc_sel_0_3 = vc_allocator_io_resp_0_vc_sel_0_3; // @[Router.scala 153:39]
  assign ingress_unit_0_from_0_io_out_credit_available_1_1 = output_unit_1_to_3_io_credit_available_1; // @[Router.scala 162:42]
  assign ingress_unit_0_from_0_io_out_credit_available_1_2 = output_unit_1_to_3_io_credit_available_2; // @[Router.scala 162:42]
  assign ingress_unit_0_from_0_io_out_credit_available_1_3 = output_unit_1_to_3_io_credit_available_3; // @[Router.scala 162:42]
  assign ingress_unit_0_from_0_io_out_credit_available_0_1 = output_unit_0_to_1_io_credit_available_1; // @[Router.scala 162:42]
  assign ingress_unit_0_from_0_io_out_credit_available_0_2 = output_unit_0_to_1_io_credit_available_2; // @[Router.scala 162:42]
  assign ingress_unit_0_from_0_io_out_credit_available_0_3 = output_unit_0_to_1_io_credit_available_3; // @[Router.scala 162:42]
  assign ingress_unit_0_from_0_io_salloc_req_0_ready = switch_allocator_io_req_0_0_ready; // @[Router.scala 165:23]
  assign ingress_unit_0_from_0_io_in_valid = auto_ingress_nodes_in_flit_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign ingress_unit_0_from_0_io_in_bits_head = auto_ingress_nodes_in_flit_bits_head; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign ingress_unit_0_from_0_io_in_bits_tail = auto_ingress_nodes_in_flit_bits_tail; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign ingress_unit_0_from_0_io_in_bits_payload = auto_ingress_nodes_in_flit_bits_payload; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign ingress_unit_0_from_0_io_in_bits_egress_id = auto_ingress_nodes_in_flit_bits_egress_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign output_unit_0_to_1_clock = clock;
  assign output_unit_0_to_1_reset = reset;
  assign output_unit_0_to_1_io_in_0_valid = switch_io_out_0_0_valid; // @[Router.scala 172:29]
  assign output_unit_0_to_1_io_in_0_bits_head = switch_io_out_0_0_bits_head; // @[Router.scala 172:29]
  assign output_unit_0_to_1_io_in_0_bits_tail = switch_io_out_0_0_bits_tail; // @[Router.scala 172:29]
  assign output_unit_0_to_1_io_in_0_bits_payload = switch_io_out_0_0_bits_payload; // @[Router.scala 172:29]
  assign output_unit_0_to_1_io_in_0_bits_flow_ingress_node = switch_io_out_0_0_bits_flow_ingress_node; // @[Router.scala 172:29]
  assign output_unit_0_to_1_io_in_0_bits_flow_egress_node = switch_io_out_0_0_bits_flow_egress_node; // @[Router.scala 172:29]
  assign output_unit_0_to_1_io_in_0_bits_virt_channel_id = switch_io_out_0_0_bits_virt_channel_id; // @[Router.scala 172:29]
  assign output_unit_0_to_1_io_allocs_1_alloc = vc_allocator_io_out_allocs_0_1_alloc; // @[Router.scala 157:33]
  assign output_unit_0_to_1_io_allocs_2_alloc = vc_allocator_io_out_allocs_0_2_alloc; // @[Router.scala 157:33]
  assign output_unit_0_to_1_io_allocs_3_alloc = vc_allocator_io_out_allocs_0_3_alloc; // @[Router.scala 157:33]
  assign output_unit_0_to_1_io_credit_alloc_1_alloc = switch_allocator_io_credit_alloc_0_1_alloc; // @[Router.scala 167:39]
  assign output_unit_0_to_1_io_credit_alloc_2_alloc = switch_allocator_io_credit_alloc_0_2_alloc; // @[Router.scala 167:39]
  assign output_unit_0_to_1_io_credit_alloc_3_alloc = switch_allocator_io_credit_alloc_0_3_alloc; // @[Router.scala 167:39]
  assign output_unit_0_to_1_io_out_credit_return = auto_source_nodes_out_0_credit_return; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign output_unit_0_to_1_io_out_vc_free = auto_source_nodes_out_0_vc_free; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign output_unit_1_to_3_clock = clock;
  assign output_unit_1_to_3_reset = reset;
  assign output_unit_1_to_3_io_in_0_valid = switch_io_out_1_0_valid; // @[Router.scala 172:29]
  assign output_unit_1_to_3_io_in_0_bits_head = switch_io_out_1_0_bits_head; // @[Router.scala 172:29]
  assign output_unit_1_to_3_io_in_0_bits_tail = switch_io_out_1_0_bits_tail; // @[Router.scala 172:29]
  assign output_unit_1_to_3_io_in_0_bits_payload = switch_io_out_1_0_bits_payload; // @[Router.scala 172:29]
  assign output_unit_1_to_3_io_in_0_bits_flow_ingress_node = switch_io_out_1_0_bits_flow_ingress_node; // @[Router.scala 172:29]
  assign output_unit_1_to_3_io_in_0_bits_flow_egress_node = switch_io_out_1_0_bits_flow_egress_node; // @[Router.scala 172:29]
  assign output_unit_1_to_3_io_in_0_bits_virt_channel_id = switch_io_out_1_0_bits_virt_channel_id; // @[Router.scala 172:29]
  assign output_unit_1_to_3_io_allocs_1_alloc = vc_allocator_io_out_allocs_1_1_alloc; // @[Router.scala 157:33]
  assign output_unit_1_to_3_io_allocs_2_alloc = vc_allocator_io_out_allocs_1_2_alloc; // @[Router.scala 157:33]
  assign output_unit_1_to_3_io_allocs_3_alloc = vc_allocator_io_out_allocs_1_3_alloc; // @[Router.scala 157:33]
  assign output_unit_1_to_3_io_credit_alloc_1_alloc = switch_allocator_io_credit_alloc_1_1_alloc; // @[Router.scala 167:39]
  assign output_unit_1_to_3_io_credit_alloc_2_alloc = switch_allocator_io_credit_alloc_1_2_alloc; // @[Router.scala 167:39]
  assign output_unit_1_to_3_io_credit_alloc_3_alloc = switch_allocator_io_credit_alloc_1_3_alloc; // @[Router.scala 167:39]
  assign output_unit_1_to_3_io_out_credit_return = auto_source_nodes_out_1_credit_return; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign output_unit_1_to_3_io_out_vc_free = auto_source_nodes_out_1_vc_free; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign switch_clock = clock;
  assign switch_reset = reset;
  assign switch_io_in_0_0_valid = ingress_unit_0_from_0_io_out_0_valid; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_head = ingress_unit_0_from_0_io_out_0_bits_flit_head; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_tail = ingress_unit_0_from_0_io_out_0_bits_flit_tail; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_payload = ingress_unit_0_from_0_io_out_0_bits_flit_payload; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_flow_ingress_node = ingress_unit_0_from_0_io_out_0_bits_flit_flow_ingress_node; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_flow_egress_node = ingress_unit_0_from_0_io_out_0_bits_flit_flow_egress_node; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_out_virt_channel = ingress_unit_0_from_0_io_out_0_bits_out_virt_channel; // @[Router.scala 170:23]
  assign switch_io_sel_1_0_0_0 = switch_io_sel_REG_1_0_0_0; // @[Router.scala 173:19]
  assign switch_io_sel_0_0_0_0 = switch_io_sel_REG_0_0_0_0; // @[Router.scala 173:19]
  assign switch_allocator_clock = clock;
  assign switch_allocator_reset = reset;
  assign switch_allocator_io_req_0_0_valid = ingress_unit_0_from_0_io_salloc_req_0_valid; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_1_0 = ingress_unit_0_from_0_io_salloc_req_0_bits_vc_sel_1_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_1_1 = ingress_unit_0_from_0_io_salloc_req_0_bits_vc_sel_1_1; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_1_2 = ingress_unit_0_from_0_io_salloc_req_0_bits_vc_sel_1_2; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_1_3 = ingress_unit_0_from_0_io_salloc_req_0_bits_vc_sel_1_3; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_0_0 = ingress_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_0_1 = ingress_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_1; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_0_2 = ingress_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_2; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_0_3 = ingress_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_3; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_tail = ingress_unit_0_from_0_io_salloc_req_0_bits_tail; // @[Router.scala 165:23]
  assign vc_allocator_clock = clock;
  assign vc_allocator_reset = reset;
  assign vc_allocator_io_req_0_valid = ingress_unit_0_from_0_io_vcalloc_req_valid; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_1_0 = ingress_unit_0_from_0_io_vcalloc_req_bits_vc_sel_1_0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_1_1 = ingress_unit_0_from_0_io_vcalloc_req_bits_vc_sel_1_1; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_1_2 = ingress_unit_0_from_0_io_vcalloc_req_bits_vc_sel_1_2; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_1_3 = ingress_unit_0_from_0_io_vcalloc_req_bits_vc_sel_1_3; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_0_0 = ingress_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_0_1 = ingress_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_1; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_0_2 = ingress_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_2; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_0_3 = ingress_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_3; // @[Router.scala 151:23]
  assign vc_allocator_io_channel_status_1_1_occupied = output_unit_1_to_3_io_channel_status_1_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_1_2_occupied = output_unit_1_to_3_io_channel_status_2_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_1_3_occupied = output_unit_1_to_3_io_channel_status_3_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_0_1_occupied = output_unit_0_to_1_io_channel_status_1_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_0_2_occupied = output_unit_0_to_1_io_channel_status_2_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_0_3_occupied = output_unit_0_to_1_io_channel_status_3_occupied; // @[Router.scala 159:23]
  assign route_computer_io_req_0_bits_flow_ingress_node = ingress_unit_0_from_0_io_router_req_bits_flow_ingress_node; // @[Router.scala 146:23]
  assign route_computer_io_req_0_bits_flow_egress_node = ingress_unit_0_from_0_io_router_req_bits_flow_egress_node; // @[Router.scala 146:23]
  always @(posedge clock) begin
    switch_io_sel_REG_1_0_0_0 <= switch_allocator_io_switch_sel_1_0_0_0; // @[Router.scala 176:14]
    switch_io_sel_REG_0_0_0_0 <= switch_allocator_io_switch_sel_0_0_0_0; // @[Router.scala 176:14]
    if (reset) begin // @[Router.scala 193:28]
      debug_tsc <= 64'h0; // @[Router.scala 193:28]
    end else begin
      debug_tsc <= _debug_tsc_T_1; // @[Router.scala 194:15]
    end
    if (reset) begin // @[Router.scala 195:31]
      debug_sample <= 64'h0; // @[Router.scala 195:31]
    end else if (debug_sample == _GEN_2) begin // @[Router.scala 198:47]
      debug_sample <= 64'h0; // @[Router.scala 198:62]
    end else begin
      debug_sample <= _debug_sample_T_1; // @[Router.scala 196:18]
    end
    if (reset) begin // @[Router.scala 201:29]
      util_ctr <= 64'h0; // @[Router.scala 201:29]
    end else begin
      util_ctr <= _util_ctr_T_1; // @[Router.scala 203:16]
    end
    if (reset) begin // @[Router.scala 202:26]
      fired <= 1'h0; // @[Router.scala 202:26]
    end else if (plusarg_reader_out != 20'h0 & _T_2 & fired) begin // @[Router.scala 205:81]
      fired <= _T_3; // @[Router.scala 208:15]
    end else begin
      fired <= fired | _T_3; // @[Router.scala 204:13]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9 & ~reset) begin
          $fwrite(32'h80000002,"nocsample %d i0 0 %d\n",debug_tsc,util_ctr); // @[Router.scala 207:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  switch_io_sel_REG_1_0_0_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  switch_io_sel_REG_0_0_0_0 = _RAND_1[0:0];
  _RAND_2 = {2{`RANDOM}};
  debug_tsc = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  debug_sample = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  util_ctr = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  fired = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ClockSinkDomain(
  output        auto_routers_ingress_nodes_in_flit_ready,
  input         auto_routers_ingress_nodes_in_flit_valid,
  input         auto_routers_ingress_nodes_in_flit_bits_head,
  input         auto_routers_ingress_nodes_in_flit_bits_tail,
  input  [63:0] auto_routers_ingress_nodes_in_flit_bits_payload,
  input         auto_routers_ingress_nodes_in_flit_bits_egress_id,
  output        auto_routers_source_nodes_out_1_flit_0_valid,
  output        auto_routers_source_nodes_out_1_flit_0_bits_head,
  output        auto_routers_source_nodes_out_1_flit_0_bits_tail,
  output [63:0] auto_routers_source_nodes_out_1_flit_0_bits_payload,
  output [1:0]  auto_routers_source_nodes_out_1_flit_0_bits_flow_ingress_node,
  output [1:0]  auto_routers_source_nodes_out_1_flit_0_bits_flow_egress_node,
  output [1:0]  auto_routers_source_nodes_out_1_flit_0_bits_virt_channel_id,
  input  [3:0]  auto_routers_source_nodes_out_1_credit_return,
  input  [3:0]  auto_routers_source_nodes_out_1_vc_free,
  output        auto_routers_source_nodes_out_0_flit_0_valid,
  output        auto_routers_source_nodes_out_0_flit_0_bits_head,
  output        auto_routers_source_nodes_out_0_flit_0_bits_tail,
  output [63:0] auto_routers_source_nodes_out_0_flit_0_bits_payload,
  output [1:0]  auto_routers_source_nodes_out_0_flit_0_bits_flow_ingress_node,
  output [1:0]  auto_routers_source_nodes_out_0_flit_0_bits_flow_egress_node,
  output [1:0]  auto_routers_source_nodes_out_0_flit_0_bits_virt_channel_id,
  input  [3:0]  auto_routers_source_nodes_out_0_credit_return,
  input  [3:0]  auto_routers_source_nodes_out_0_vc_free,
  input         auto_clock_in_clock,
  input         auto_clock_in_reset
);
  wire  routers_clock; // @[NoC.scala 64:22]
  wire  routers_reset; // @[NoC.scala 64:22]
  wire  routers_auto_ingress_nodes_in_flit_ready; // @[NoC.scala 64:22]
  wire  routers_auto_ingress_nodes_in_flit_valid; // @[NoC.scala 64:22]
  wire  routers_auto_ingress_nodes_in_flit_bits_head; // @[NoC.scala 64:22]
  wire  routers_auto_ingress_nodes_in_flit_bits_tail; // @[NoC.scala 64:22]
  wire [63:0] routers_auto_ingress_nodes_in_flit_bits_payload; // @[NoC.scala 64:22]
  wire  routers_auto_ingress_nodes_in_flit_bits_egress_id; // @[NoC.scala 64:22]
  wire  routers_auto_source_nodes_out_1_flit_0_valid; // @[NoC.scala 64:22]
  wire  routers_auto_source_nodes_out_1_flit_0_bits_head; // @[NoC.scala 64:22]
  wire  routers_auto_source_nodes_out_1_flit_0_bits_tail; // @[NoC.scala 64:22]
  wire [63:0] routers_auto_source_nodes_out_1_flit_0_bits_payload; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_source_nodes_out_1_flit_0_bits_flow_ingress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_source_nodes_out_1_flit_0_bits_flow_egress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_source_nodes_out_1_flit_0_bits_virt_channel_id; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_source_nodes_out_1_credit_return; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_source_nodes_out_1_vc_free; // @[NoC.scala 64:22]
  wire  routers_auto_source_nodes_out_0_flit_0_valid; // @[NoC.scala 64:22]
  wire  routers_auto_source_nodes_out_0_flit_0_bits_head; // @[NoC.scala 64:22]
  wire  routers_auto_source_nodes_out_0_flit_0_bits_tail; // @[NoC.scala 64:22]
  wire [63:0] routers_auto_source_nodes_out_0_flit_0_bits_payload; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_source_nodes_out_0_flit_0_bits_flow_ingress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_source_nodes_out_0_flit_0_bits_flow_egress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_source_nodes_out_0_flit_0_bits_virt_channel_id; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_source_nodes_out_0_credit_return; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_source_nodes_out_0_vc_free; // @[NoC.scala 64:22]
  Router routers ( // @[NoC.scala 64:22]
    .clock(routers_clock),
    .reset(routers_reset),
    .auto_ingress_nodes_in_flit_ready(routers_auto_ingress_nodes_in_flit_ready),
    .auto_ingress_nodes_in_flit_valid(routers_auto_ingress_nodes_in_flit_valid),
    .auto_ingress_nodes_in_flit_bits_head(routers_auto_ingress_nodes_in_flit_bits_head),
    .auto_ingress_nodes_in_flit_bits_tail(routers_auto_ingress_nodes_in_flit_bits_tail),
    .auto_ingress_nodes_in_flit_bits_payload(routers_auto_ingress_nodes_in_flit_bits_payload),
    .auto_ingress_nodes_in_flit_bits_egress_id(routers_auto_ingress_nodes_in_flit_bits_egress_id),
    .auto_source_nodes_out_1_flit_0_valid(routers_auto_source_nodes_out_1_flit_0_valid),
    .auto_source_nodes_out_1_flit_0_bits_head(routers_auto_source_nodes_out_1_flit_0_bits_head),
    .auto_source_nodes_out_1_flit_0_bits_tail(routers_auto_source_nodes_out_1_flit_0_bits_tail),
    .auto_source_nodes_out_1_flit_0_bits_payload(routers_auto_source_nodes_out_1_flit_0_bits_payload),
    .auto_source_nodes_out_1_flit_0_bits_flow_ingress_node(routers_auto_source_nodes_out_1_flit_0_bits_flow_ingress_node
      ),
    .auto_source_nodes_out_1_flit_0_bits_flow_egress_node(routers_auto_source_nodes_out_1_flit_0_bits_flow_egress_node),
    .auto_source_nodes_out_1_flit_0_bits_virt_channel_id(routers_auto_source_nodes_out_1_flit_0_bits_virt_channel_id),
    .auto_source_nodes_out_1_credit_return(routers_auto_source_nodes_out_1_credit_return),
    .auto_source_nodes_out_1_vc_free(routers_auto_source_nodes_out_1_vc_free),
    .auto_source_nodes_out_0_flit_0_valid(routers_auto_source_nodes_out_0_flit_0_valid),
    .auto_source_nodes_out_0_flit_0_bits_head(routers_auto_source_nodes_out_0_flit_0_bits_head),
    .auto_source_nodes_out_0_flit_0_bits_tail(routers_auto_source_nodes_out_0_flit_0_bits_tail),
    .auto_source_nodes_out_0_flit_0_bits_payload(routers_auto_source_nodes_out_0_flit_0_bits_payload),
    .auto_source_nodes_out_0_flit_0_bits_flow_ingress_node(routers_auto_source_nodes_out_0_flit_0_bits_flow_ingress_node
      ),
    .auto_source_nodes_out_0_flit_0_bits_flow_egress_node(routers_auto_source_nodes_out_0_flit_0_bits_flow_egress_node),
    .auto_source_nodes_out_0_flit_0_bits_virt_channel_id(routers_auto_source_nodes_out_0_flit_0_bits_virt_channel_id),
    .auto_source_nodes_out_0_credit_return(routers_auto_source_nodes_out_0_credit_return),
    .auto_source_nodes_out_0_vc_free(routers_auto_source_nodes_out_0_vc_free)
  );
  assign auto_routers_ingress_nodes_in_flit_ready = routers_auto_ingress_nodes_in_flit_ready; // @[LazyModule.scala 366:16]
  assign auto_routers_source_nodes_out_1_flit_0_valid = routers_auto_source_nodes_out_1_flit_0_valid; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_1_flit_0_bits_head = routers_auto_source_nodes_out_1_flit_0_bits_head; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_1_flit_0_bits_tail = routers_auto_source_nodes_out_1_flit_0_bits_tail; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_1_flit_0_bits_payload = routers_auto_source_nodes_out_1_flit_0_bits_payload; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_1_flit_0_bits_flow_ingress_node =
    routers_auto_source_nodes_out_1_flit_0_bits_flow_ingress_node; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_1_flit_0_bits_flow_egress_node =
    routers_auto_source_nodes_out_1_flit_0_bits_flow_egress_node; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_1_flit_0_bits_virt_channel_id =
    routers_auto_source_nodes_out_1_flit_0_bits_virt_channel_id; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_0_flit_0_valid = routers_auto_source_nodes_out_0_flit_0_valid; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_0_flit_0_bits_head = routers_auto_source_nodes_out_0_flit_0_bits_head; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_0_flit_0_bits_tail = routers_auto_source_nodes_out_0_flit_0_bits_tail; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_0_flit_0_bits_payload = routers_auto_source_nodes_out_0_flit_0_bits_payload; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_0_flit_0_bits_flow_ingress_node =
    routers_auto_source_nodes_out_0_flit_0_bits_flow_ingress_node; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_0_flit_0_bits_flow_egress_node =
    routers_auto_source_nodes_out_0_flit_0_bits_flow_egress_node; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_0_flit_0_bits_virt_channel_id =
    routers_auto_source_nodes_out_0_flit_0_bits_virt_channel_id; // @[LazyModule.scala 368:12]
  assign routers_clock = auto_clock_in_clock; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign routers_reset = auto_clock_in_reset; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign routers_auto_ingress_nodes_in_flit_valid = auto_routers_ingress_nodes_in_flit_valid; // @[LazyModule.scala 366:16]
  assign routers_auto_ingress_nodes_in_flit_bits_head = auto_routers_ingress_nodes_in_flit_bits_head; // @[LazyModule.scala 366:16]
  assign routers_auto_ingress_nodes_in_flit_bits_tail = auto_routers_ingress_nodes_in_flit_bits_tail; // @[LazyModule.scala 366:16]
  assign routers_auto_ingress_nodes_in_flit_bits_payload = auto_routers_ingress_nodes_in_flit_bits_payload; // @[LazyModule.scala 366:16]
  assign routers_auto_ingress_nodes_in_flit_bits_egress_id = auto_routers_ingress_nodes_in_flit_bits_egress_id; // @[LazyModule.scala 366:16]
  assign routers_auto_source_nodes_out_1_credit_return = auto_routers_source_nodes_out_1_credit_return; // @[LazyModule.scala 368:12]
  assign routers_auto_source_nodes_out_1_vc_free = auto_routers_source_nodes_out_1_vc_free; // @[LazyModule.scala 368:12]
  assign routers_auto_source_nodes_out_0_credit_return = auto_routers_source_nodes_out_0_credit_return; // @[LazyModule.scala 368:12]
  assign routers_auto_source_nodes_out_0_vc_free = auto_routers_source_nodes_out_0_vc_free; // @[LazyModule.scala 368:12]
endmodule
module NoCMonitor(
  input        clock,
  input        reset,
  input        io_in_flit_0_valid,
  input        io_in_flit_0_bits_head,
  input        io_in_flit_0_bits_tail,
  input  [1:0] io_in_flit_0_bits_flow_ingress_node,
  input  [1:0] io_in_flit_0_bits_flow_egress_node,
  input  [1:0] io_in_flit_0_bits_virt_channel_id
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg  in_flight_0; // @[Monitor.scala 16:26]
  reg  in_flight_1; // @[Monitor.scala 16:26]
  reg  in_flight_2; // @[Monitor.scala 16:26]
  reg  in_flight_3; // @[Monitor.scala 16:26]
  wire  _GEN_0 = 2'h0 == io_in_flit_0_bits_virt_channel_id | in_flight_0; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_1 = 2'h1 == io_in_flit_0_bits_virt_channel_id | in_flight_1; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_2 = 2'h2 == io_in_flit_0_bits_virt_channel_id | in_flight_2; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_3 = 2'h3 == io_in_flit_0_bits_virt_channel_id | in_flight_3; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_5 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? in_flight_1 : in_flight_0; // @[Monitor.scala 22:{17,17}]
  wire  _GEN_6 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? in_flight_2 : _GEN_5; // @[Monitor.scala 22:{17,17}]
  wire  _GEN_7 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? in_flight_3 : _GEN_6; // @[Monitor.scala 22:{17,17}]
  wire  _T_2 = ~reset; // @[Monitor.scala 22:16]
  wire  _GEN_8 = io_in_flit_0_bits_head ? _GEN_0 : in_flight_0; // @[Monitor.scala 16:26 20:29]
  wire  _GEN_9 = io_in_flit_0_bits_head ? _GEN_1 : in_flight_1; // @[Monitor.scala 16:26 20:29]
  wire  _GEN_10 = io_in_flit_0_bits_head ? _GEN_2 : in_flight_2; // @[Monitor.scala 16:26 20:29]
  wire  _GEN_11 = io_in_flit_0_bits_head ? _GEN_3 : in_flight_3; // @[Monitor.scala 16:26 20:29]
  wire  _T_4 = io_in_flit_0_valid & io_in_flit_0_bits_head; // @[Monitor.scala 29:22]
  wire  _T_12 = io_in_flit_0_bits_flow_egress_node == 2'h1; // @[Types.scala 54:21]
  wire  _T_13 = io_in_flit_0_bits_flow_ingress_node == 2'h0 & _T_12; // @[Types.scala 53:39]
  wire  _GEN_29 = _T_4 & ~reset; // @[Monitor.scala 22:16]
  always @(posedge clock) begin
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_0 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h0 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_0 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_0 <= _GEN_8;
        end
      end else begin
        in_flight_0 <= _GEN_8;
      end
    end
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_1 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h1 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_1 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_1 <= _GEN_9;
        end
      end else begin
        in_flight_1 <= _GEN_9;
      end
    end
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_2 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h2 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_2 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_2 <= _GEN_10;
        end
      end else begin
        in_flight_2 <= _GEN_10;
      end
    end
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_3 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h3 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_3 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_3 <= _GEN_11;
        end
      end else begin
        in_flight_3 <= _GEN_11;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4 & ~reset & ~(~_GEN_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed: Flit head/tail sequencing is broken\n    at Monitor.scala:22 assert (!in_flight(flit.bits.virt_channel_id), \"Flit head/tail sequencing is broken\")\n"
            ); // @[Monitor.scala 22:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h1 | _T_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h2 | _T_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h3 | _T_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  in_flight_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  in_flight_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  in_flight_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  in_flight_3 = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (_T_4 & ~reset) begin
      assert(~_GEN_7); // @[Monitor.scala 22:16]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h0); // @[Monitor.scala 32:17]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h1 | _T_13); // @[Monitor.scala 32:17]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h2 | _T_13); // @[Monitor.scala 32:17]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h3 | _T_13); // @[Monitor.scala 32:17]
    end
  end
endmodule
module NoCMonitor_1(
  input        clock,
  input        reset,
  input        io_in_flit_0_valid,
  input        io_in_flit_0_bits_head,
  input        io_in_flit_0_bits_tail,
  input  [1:0] io_in_flit_0_bits_flow_ingress_node,
  input  [1:0] io_in_flit_0_bits_flow_egress_node,
  input  [1:0] io_in_flit_0_bits_virt_channel_id
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg  in_flight_0; // @[Monitor.scala 16:26]
  reg  in_flight_1; // @[Monitor.scala 16:26]
  reg  in_flight_2; // @[Monitor.scala 16:26]
  reg  in_flight_3; // @[Monitor.scala 16:26]
  wire  _GEN_0 = 2'h0 == io_in_flit_0_bits_virt_channel_id | in_flight_0; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_1 = 2'h1 == io_in_flit_0_bits_virt_channel_id | in_flight_1; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_2 = 2'h2 == io_in_flit_0_bits_virt_channel_id | in_flight_2; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_3 = 2'h3 == io_in_flit_0_bits_virt_channel_id | in_flight_3; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_5 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? in_flight_1 : in_flight_0; // @[Monitor.scala 22:{17,17}]
  wire  _GEN_6 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? in_flight_2 : _GEN_5; // @[Monitor.scala 22:{17,17}]
  wire  _GEN_7 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? in_flight_3 : _GEN_6; // @[Monitor.scala 22:{17,17}]
  wire  _T_2 = ~reset; // @[Monitor.scala 22:16]
  wire  _GEN_8 = io_in_flit_0_bits_head ? _GEN_0 : in_flight_0; // @[Monitor.scala 16:26 20:29]
  wire  _GEN_9 = io_in_flit_0_bits_head ? _GEN_1 : in_flight_1; // @[Monitor.scala 16:26 20:29]
  wire  _GEN_10 = io_in_flit_0_bits_head ? _GEN_2 : in_flight_2; // @[Monitor.scala 16:26 20:29]
  wire  _GEN_11 = io_in_flit_0_bits_head ? _GEN_3 : in_flight_3; // @[Monitor.scala 16:26 20:29]
  wire  _T_4 = io_in_flit_0_valid & io_in_flit_0_bits_head; // @[Monitor.scala 29:22]
  wire  _T_12 = io_in_flit_0_bits_flow_egress_node == 2'h1; // @[Types.scala 54:21]
  wire  _T_13 = io_in_flit_0_bits_flow_ingress_node == 2'h2 & _T_12; // @[Types.scala 53:39]
  wire  _GEN_29 = _T_4 & ~reset; // @[Monitor.scala 22:16]
  always @(posedge clock) begin
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_0 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h0 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_0 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_0 <= _GEN_8;
        end
      end else begin
        in_flight_0 <= _GEN_8;
      end
    end
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_1 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h1 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_1 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_1 <= _GEN_9;
        end
      end else begin
        in_flight_1 <= _GEN_9;
      end
    end
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_2 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h2 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_2 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_2 <= _GEN_10;
        end
      end else begin
        in_flight_2 <= _GEN_10;
      end
    end
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_3 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h3 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_3 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_3 <= _GEN_11;
        end
      end else begin
        in_flight_3 <= _GEN_11;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4 & ~reset & ~(~_GEN_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed: Flit head/tail sequencing is broken\n    at Monitor.scala:22 assert (!in_flight(flit.bits.virt_channel_id), \"Flit head/tail sequencing is broken\")\n"
            ); // @[Monitor.scala 22:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h1 | _T_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h2 | _T_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h3 | _T_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  in_flight_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  in_flight_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  in_flight_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  in_flight_3 = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (_T_4 & ~reset) begin
      assert(~_GEN_7); // @[Monitor.scala 22:16]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h0); // @[Monitor.scala 32:17]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h1 | _T_13); // @[Monitor.scala 32:17]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h2 | _T_13); // @[Monitor.scala 32:17]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h3 | _T_13); // @[Monitor.scala 32:17]
    end
  end
endmodule
module Queue_4(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_head,
  input         io_enq_bits_tail,
  input  [63:0] io_enq_bits_payload,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_head,
  output        io_deq_bits_tail,
  output [63:0] io_deq_bits_payload
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg  ram_head [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_head_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_head_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_head_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_tail [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_tail_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_tail_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_tail_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_en; // @[Decoupled.scala 273:95]
  reg [63:0] ram_payload [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_payload_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_payload_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [63:0] ram_payload_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [63:0] ram_payload_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_payload_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_payload_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_payload_MPORT_en; // @[Decoupled.scala 273:95]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 278:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  assign ram_head_io_deq_bits_MPORT_en = 1'h1;
  assign ram_head_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_head_io_deq_bits_MPORT_data = ram_head[ram_head_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_head_MPORT_data = io_enq_bits_head;
  assign ram_head_MPORT_addr = 1'h0;
  assign ram_head_MPORT_mask = 1'h1;
  assign ram_head_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tail_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tail_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tail_io_deq_bits_MPORT_data = ram_tail[ram_tail_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_tail_MPORT_data = io_enq_bits_tail;
  assign ram_tail_MPORT_addr = 1'h0;
  assign ram_tail_MPORT_mask = 1'h1;
  assign ram_tail_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_payload_io_deq_bits_MPORT_en = 1'h1;
  assign ram_payload_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_payload_io_deq_bits_MPORT_data = ram_payload[ram_payload_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_payload_MPORT_data = io_enq_bits_payload;
  assign ram_payload_MPORT_addr = 1'h0;
  assign ram_payload_MPORT_mask = 1'h1;
  assign ram_payload_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = io_deq_ready | empty; // @[Decoupled.scala 303:16 323:{24,39}]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_head = ram_head_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_tail = ram_tail_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_payload = ram_payload_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  always @(posedge clock) begin
    if (ram_head_MPORT_en & ram_head_MPORT_mask) begin
      ram_head[ram_head_MPORT_addr] <= ram_head_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_tail_MPORT_en & ram_tail_MPORT_mask) begin
      ram_tail[ram_tail_MPORT_addr] <= ram_tail_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_payload_MPORT_en & ram_payload_MPORT_mask) begin
      ram_payload[ram_payload_MPORT_addr] <= ram_payload_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_head[initvar] = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tail[initvar] = _RAND_1[0:0];
  _RAND_2 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload[initvar] = _RAND_2[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module InputBuffer(
  input         clock,
  input         reset,
  input         io_enq_0_valid,
  input         io_enq_0_bits_head,
  input         io_enq_0_bits_tail,
  input  [63:0] io_enq_0_bits_payload,
  input  [1:0]  io_enq_0_bits_virt_channel_id,
  output        io_deq_0_bits_head,
  output        io_deq_0_bits_tail,
  output [63:0] io_deq_0_bits_payload,
  input         io_deq_1_ready,
  output        io_deq_1_valid,
  output        io_deq_1_bits_head,
  output        io_deq_1_bits_tail,
  output [63:0] io_deq_1_bits_payload,
  input         io_deq_2_ready,
  output        io_deq_2_valid,
  output        io_deq_2_bits_head,
  output        io_deq_2_bits_tail,
  output [63:0] io_deq_2_bits_payload,
  input         io_deq_3_ready,
  output        io_deq_3_valid,
  output        io_deq_3_bits_head,
  output        io_deq_3_bits_tail,
  output [63:0] io_deq_3_bits_payload
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_10;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
`endif // RANDOMIZE_REG_INIT
  reg  mem_head [0:14]; // @[InputUnit.scala 85:18]
  wire  mem_head_qs_0_io_enq_bits_MPORT_en; // @[InputUnit.scala 85:18]
  wire [3:0] mem_head_qs_0_io_enq_bits_MPORT_addr; // @[InputUnit.scala 85:18]
  wire  mem_head_qs_0_io_enq_bits_MPORT_data; // @[InputUnit.scala 85:18]
  wire  mem_head_qs_1_io_enq_bits_MPORT_en; // @[InputUnit.scala 85:18]
  wire [3:0] mem_head_qs_1_io_enq_bits_MPORT_addr; // @[InputUnit.scala 85:18]
  wire  mem_head_qs_1_io_enq_bits_MPORT_data; // @[InputUnit.scala 85:18]
  wire  mem_head_qs_2_io_enq_bits_MPORT_en; // @[InputUnit.scala 85:18]
  wire [3:0] mem_head_qs_2_io_enq_bits_MPORT_addr; // @[InputUnit.scala 85:18]
  wire  mem_head_qs_2_io_enq_bits_MPORT_data; // @[InputUnit.scala 85:18]
  wire  mem_head_qs_3_io_enq_bits_MPORT_en; // @[InputUnit.scala 85:18]
  wire [3:0] mem_head_qs_3_io_enq_bits_MPORT_addr; // @[InputUnit.scala 85:18]
  wire  mem_head_qs_3_io_enq_bits_MPORT_data; // @[InputUnit.scala 85:18]
  wire  mem_head_MPORT_data; // @[InputUnit.scala 85:18]
  wire [3:0] mem_head_MPORT_addr; // @[InputUnit.scala 85:18]
  wire  mem_head_MPORT_mask; // @[InputUnit.scala 85:18]
  wire  mem_head_MPORT_en; // @[InputUnit.scala 85:18]
  reg  mem_tail [0:14]; // @[InputUnit.scala 85:18]
  wire  mem_tail_qs_0_io_enq_bits_MPORT_en; // @[InputUnit.scala 85:18]
  wire [3:0] mem_tail_qs_0_io_enq_bits_MPORT_addr; // @[InputUnit.scala 85:18]
  wire  mem_tail_qs_0_io_enq_bits_MPORT_data; // @[InputUnit.scala 85:18]
  wire  mem_tail_qs_1_io_enq_bits_MPORT_en; // @[InputUnit.scala 85:18]
  wire [3:0] mem_tail_qs_1_io_enq_bits_MPORT_addr; // @[InputUnit.scala 85:18]
  wire  mem_tail_qs_1_io_enq_bits_MPORT_data; // @[InputUnit.scala 85:18]
  wire  mem_tail_qs_2_io_enq_bits_MPORT_en; // @[InputUnit.scala 85:18]
  wire [3:0] mem_tail_qs_2_io_enq_bits_MPORT_addr; // @[InputUnit.scala 85:18]
  wire  mem_tail_qs_2_io_enq_bits_MPORT_data; // @[InputUnit.scala 85:18]
  wire  mem_tail_qs_3_io_enq_bits_MPORT_en; // @[InputUnit.scala 85:18]
  wire [3:0] mem_tail_qs_3_io_enq_bits_MPORT_addr; // @[InputUnit.scala 85:18]
  wire  mem_tail_qs_3_io_enq_bits_MPORT_data; // @[InputUnit.scala 85:18]
  wire  mem_tail_MPORT_data; // @[InputUnit.scala 85:18]
  wire [3:0] mem_tail_MPORT_addr; // @[InputUnit.scala 85:18]
  wire  mem_tail_MPORT_mask; // @[InputUnit.scala 85:18]
  wire  mem_tail_MPORT_en; // @[InputUnit.scala 85:18]
  reg [63:0] mem_payload [0:14]; // @[InputUnit.scala 85:18]
  wire  mem_payload_qs_0_io_enq_bits_MPORT_en; // @[InputUnit.scala 85:18]
  wire [3:0] mem_payload_qs_0_io_enq_bits_MPORT_addr; // @[InputUnit.scala 85:18]
  wire [63:0] mem_payload_qs_0_io_enq_bits_MPORT_data; // @[InputUnit.scala 85:18]
  wire  mem_payload_qs_1_io_enq_bits_MPORT_en; // @[InputUnit.scala 85:18]
  wire [3:0] mem_payload_qs_1_io_enq_bits_MPORT_addr; // @[InputUnit.scala 85:18]
  wire [63:0] mem_payload_qs_1_io_enq_bits_MPORT_data; // @[InputUnit.scala 85:18]
  wire  mem_payload_qs_2_io_enq_bits_MPORT_en; // @[InputUnit.scala 85:18]
  wire [3:0] mem_payload_qs_2_io_enq_bits_MPORT_addr; // @[InputUnit.scala 85:18]
  wire [63:0] mem_payload_qs_2_io_enq_bits_MPORT_data; // @[InputUnit.scala 85:18]
  wire  mem_payload_qs_3_io_enq_bits_MPORT_en; // @[InputUnit.scala 85:18]
  wire [3:0] mem_payload_qs_3_io_enq_bits_MPORT_addr; // @[InputUnit.scala 85:18]
  wire [63:0] mem_payload_qs_3_io_enq_bits_MPORT_data; // @[InputUnit.scala 85:18]
  wire [63:0] mem_payload_MPORT_data; // @[InputUnit.scala 85:18]
  wire [3:0] mem_payload_MPORT_addr; // @[InputUnit.scala 85:18]
  wire  mem_payload_MPORT_mask; // @[InputUnit.scala 85:18]
  wire  mem_payload_MPORT_en; // @[InputUnit.scala 85:18]
  wire  qs_0_clock; // @[InputUnit.scala 90:49]
  wire  qs_0_reset; // @[InputUnit.scala 90:49]
  wire  qs_0_io_enq_ready; // @[InputUnit.scala 90:49]
  wire  qs_0_io_enq_valid; // @[InputUnit.scala 90:49]
  wire  qs_0_io_enq_bits_head; // @[InputUnit.scala 90:49]
  wire  qs_0_io_enq_bits_tail; // @[InputUnit.scala 90:49]
  wire [63:0] qs_0_io_enq_bits_payload; // @[InputUnit.scala 90:49]
  wire  qs_0_io_deq_ready; // @[InputUnit.scala 90:49]
  wire  qs_0_io_deq_valid; // @[InputUnit.scala 90:49]
  wire  qs_0_io_deq_bits_head; // @[InputUnit.scala 90:49]
  wire  qs_0_io_deq_bits_tail; // @[InputUnit.scala 90:49]
  wire [63:0] qs_0_io_deq_bits_payload; // @[InputUnit.scala 90:49]
  wire  qs_1_clock; // @[InputUnit.scala 90:49]
  wire  qs_1_reset; // @[InputUnit.scala 90:49]
  wire  qs_1_io_enq_ready; // @[InputUnit.scala 90:49]
  wire  qs_1_io_enq_valid; // @[InputUnit.scala 90:49]
  wire  qs_1_io_enq_bits_head; // @[InputUnit.scala 90:49]
  wire  qs_1_io_enq_bits_tail; // @[InputUnit.scala 90:49]
  wire [63:0] qs_1_io_enq_bits_payload; // @[InputUnit.scala 90:49]
  wire  qs_1_io_deq_ready; // @[InputUnit.scala 90:49]
  wire  qs_1_io_deq_valid; // @[InputUnit.scala 90:49]
  wire  qs_1_io_deq_bits_head; // @[InputUnit.scala 90:49]
  wire  qs_1_io_deq_bits_tail; // @[InputUnit.scala 90:49]
  wire [63:0] qs_1_io_deq_bits_payload; // @[InputUnit.scala 90:49]
  wire  qs_2_clock; // @[InputUnit.scala 90:49]
  wire  qs_2_reset; // @[InputUnit.scala 90:49]
  wire  qs_2_io_enq_ready; // @[InputUnit.scala 90:49]
  wire  qs_2_io_enq_valid; // @[InputUnit.scala 90:49]
  wire  qs_2_io_enq_bits_head; // @[InputUnit.scala 90:49]
  wire  qs_2_io_enq_bits_tail; // @[InputUnit.scala 90:49]
  wire [63:0] qs_2_io_enq_bits_payload; // @[InputUnit.scala 90:49]
  wire  qs_2_io_deq_ready; // @[InputUnit.scala 90:49]
  wire  qs_2_io_deq_valid; // @[InputUnit.scala 90:49]
  wire  qs_2_io_deq_bits_head; // @[InputUnit.scala 90:49]
  wire  qs_2_io_deq_bits_tail; // @[InputUnit.scala 90:49]
  wire [63:0] qs_2_io_deq_bits_payload; // @[InputUnit.scala 90:49]
  wire  qs_3_clock; // @[InputUnit.scala 90:49]
  wire  qs_3_reset; // @[InputUnit.scala 90:49]
  wire  qs_3_io_enq_ready; // @[InputUnit.scala 90:49]
  wire  qs_3_io_enq_valid; // @[InputUnit.scala 90:49]
  wire  qs_3_io_enq_bits_head; // @[InputUnit.scala 90:49]
  wire  qs_3_io_enq_bits_tail; // @[InputUnit.scala 90:49]
  wire [63:0] qs_3_io_enq_bits_payload; // @[InputUnit.scala 90:49]
  wire  qs_3_io_deq_ready; // @[InputUnit.scala 90:49]
  wire  qs_3_io_deq_valid; // @[InputUnit.scala 90:49]
  wire  qs_3_io_deq_bits_head; // @[InputUnit.scala 90:49]
  wire  qs_3_io_deq_bits_tail; // @[InputUnit.scala 90:49]
  wire [63:0] qs_3_io_deq_bits_payload; // @[InputUnit.scala 90:49]
  reg [3:0] heads_0; // @[InputUnit.scala 86:24]
  reg [3:0] heads_1; // @[InputUnit.scala 86:24]
  reg [3:0] heads_2; // @[InputUnit.scala 86:24]
  reg [3:0] heads_3; // @[InputUnit.scala 86:24]
  reg [3:0] tails_0; // @[InputUnit.scala 87:24]
  reg [3:0] tails_1; // @[InputUnit.scala 87:24]
  reg [3:0] tails_2; // @[InputUnit.scala 87:24]
  reg [3:0] tails_3; // @[InputUnit.scala 87:24]
  wire  empty_0 = heads_0 == tails_0; // @[InputUnit.scala 88:49]
  wire  empty_1 = heads_1 == tails_1; // @[InputUnit.scala 88:49]
  wire  empty_2 = heads_2 == tails_2; // @[InputUnit.scala 88:49]
  wire  empty_3 = heads_3 == tails_3; // @[InputUnit.scala 88:49]
  wire [3:0] vc_sel = 4'h1 << io_enq_0_bits_virt_channel_id; // @[OneHot.scala 57:35]
  wire  _direct_to_q_T_10 = vc_sel[0] & qs_0_io_enq_ready | vc_sel[1] & qs_1_io_enq_ready | vc_sel[2] &
    qs_2_io_enq_ready | vc_sel[3] & qs_3_io_enq_ready; // @[Mux.scala 27:73]
  wire  _direct_to_q_T_21 = vc_sel[0] & empty_0 | vc_sel[1] & empty_1 | vc_sel[2] & empty_2 | vc_sel[3] & empty_3; // @[Mux.scala 27:73]
  wire  direct_to_q = _direct_to_q_T_10 & _direct_to_q_T_21; // @[InputUnit.scala 96:62]
  wire  _T = ~direct_to_q; // @[InputUnit.scala 100:30]
  wire [3:0] _GEN_1 = 2'h1 == io_enq_0_bits_virt_channel_id ? tails_1 : tails_0; // @[]
  wire [3:0] _GEN_2 = 2'h2 == io_enq_0_bits_virt_channel_id ? tails_2 : _GEN_1; // @[]
  wire [3:0] _GEN_3 = 2'h3 == io_enq_0_bits_virt_channel_id ? tails_3 : _GEN_2; // @[]
  wire [2:0] _tails_T_5 = vc_sel[1] ? 3'h4 : 3'h0; // @[Mux.scala 27:73]
  wire [3:0] _tails_T_6 = vc_sel[2] ? 4'h9 : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _tails_T_7 = vc_sel[3] ? 4'he : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _GEN_131 = {{1'd0}, _tails_T_5}; // @[Mux.scala 27:73]
  wire [3:0] _tails_T_9 = _GEN_131 | _tails_T_6; // @[Mux.scala 27:73]
  wire [3:0] _tails_T_10 = _tails_T_9 | _tails_T_7; // @[Mux.scala 27:73]
  wire  _tails_T_11 = _GEN_3 == _tails_T_10; // @[InputUnit.scala 104:14]
  wire [2:0] _tails_T_18 = vc_sel[2] ? 3'h5 : 3'h0; // @[Mux.scala 27:73]
  wire [3:0] _tails_T_19 = vc_sel[3] ? 4'ha : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _GEN_132 = {{1'd0}, _tails_T_18}; // @[Mux.scala 27:73]
  wire [3:0] _tails_T_22 = _GEN_132 | _tails_T_19; // @[Mux.scala 27:73]
  wire [3:0] _tails_T_24 = _GEN_3 + 4'h1; // @[InputUnit.scala 106:14]
  wire  _T_3 = io_enq_0_bits_virt_channel_id == 2'h0; // @[InputUnit.scala 109:46]
  wire  _T_4 = io_enq_0_bits_virt_channel_id == 2'h1; // @[InputUnit.scala 109:46]
  wire  _T_5 = io_enq_0_bits_virt_channel_id == 2'h2; // @[InputUnit.scala 109:46]
  wire  _T_6 = io_enq_0_bits_virt_channel_id == 2'h3; // @[InputUnit.scala 109:46]
  wire  _GEN_24 = io_enq_0_valid & direct_to_q & _T_3; // @[InputUnit.scala 107:50 91:31]
  wire  _GEN_28 = io_enq_0_valid & direct_to_q & _T_4; // @[InputUnit.scala 107:50 91:31]
  wire  _GEN_32 = io_enq_0_valid & direct_to_q & _T_5; // @[InputUnit.scala 107:50 91:31]
  wire  _GEN_36 = io_enq_0_valid & direct_to_q & _T_6; // @[InputUnit.scala 107:50 91:31]
  wire  _GEN_51 = io_enq_0_valid & ~direct_to_q ? 1'h0 : _GEN_24; // @[InputUnit.scala 100:44 91:31]
  wire  _GEN_55 = io_enq_0_valid & ~direct_to_q ? 1'h0 : _GEN_28; // @[InputUnit.scala 100:44 91:31]
  wire  _GEN_59 = io_enq_0_valid & ~direct_to_q ? 1'h0 : _GEN_32; // @[InputUnit.scala 100:44 91:31]
  wire  _GEN_63 = io_enq_0_valid & ~direct_to_q ? 1'h0 : _GEN_36; // @[InputUnit.scala 100:44 91:31]
  wire  can_to_q_0 = ~empty_0 & qs_0_io_enq_ready; // @[InputUnit.scala 117:70]
  wire  can_to_q_1 = ~empty_1 & qs_1_io_enq_ready; // @[InputUnit.scala 117:70]
  wire  can_to_q_2 = ~empty_2 & qs_2_io_enq_ready; // @[InputUnit.scala 117:70]
  wire  can_to_q_3 = ~empty_3 & qs_3_io_enq_ready; // @[InputUnit.scala 117:70]
  wire [3:0] _to_q_oh_enc_T = can_to_q_3 ? 4'h8 : 4'h0; // @[Mux.scala 47:70]
  wire [3:0] _to_q_oh_enc_T_1 = can_to_q_2 ? 4'h4 : _to_q_oh_enc_T; // @[Mux.scala 47:70]
  wire [3:0] _to_q_oh_enc_T_2 = can_to_q_1 ? 4'h2 : _to_q_oh_enc_T_1; // @[Mux.scala 47:70]
  wire [3:0] to_q_oh_enc = can_to_q_0 ? 4'h1 : _to_q_oh_enc_T_2; // @[Mux.scala 47:70]
  wire  to_q_oh_0 = to_q_oh_enc[0]; // @[OneHot.scala 82:30]
  wire  to_q_oh_1 = to_q_oh_enc[1]; // @[OneHot.scala 82:30]
  wire  to_q_oh_2 = to_q_oh_enc[2]; // @[OneHot.scala 82:30]
  wire  to_q_oh_3 = to_q_oh_enc[3]; // @[OneHot.scala 82:30]
  wire [3:0] _to_q_T = {to_q_oh_3,to_q_oh_2,to_q_oh_1,to_q_oh_0}; // @[Cat.scala 33:92]
  wire [1:0] to_q_hi_1 = _to_q_T[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] to_q_lo_1 = _to_q_T[1:0]; // @[OneHot.scala 31:18]
  wire  _to_q_T_1 = |to_q_hi_1; // @[OneHot.scala 32:14]
  wire [1:0] _to_q_T_2 = to_q_hi_1 | to_q_lo_1; // @[OneHot.scala 32:28]
  wire [1:0] to_q = {_to_q_T_1,_to_q_T_2[1]}; // @[Cat.scala 33:92]
  wire  _T_9 = can_to_q_0 | can_to_q_1 | can_to_q_2 | can_to_q_3; // @[package.scala 73:59]
  wire [3:0] _head_T = to_q_oh_0 ? heads_0 : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _head_T_1 = to_q_oh_1 ? heads_1 : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _head_T_2 = to_q_oh_2 ? heads_2 : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _head_T_3 = to_q_oh_3 ? heads_3 : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _head_T_4 = _head_T | _head_T_1; // @[Mux.scala 27:73]
  wire [3:0] _head_T_5 = _head_T_4 | _head_T_2; // @[Mux.scala 27:73]
  wire [3:0] head = _head_T_5 | _head_T_3; // @[Mux.scala 27:73]
  wire [2:0] _heads_T_1 = to_q_oh_1 ? 3'h4 : 3'h0; // @[Mux.scala 27:73]
  wire [3:0] _heads_T_2 = to_q_oh_2 ? 4'h9 : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _heads_T_3 = to_q_oh_3 ? 4'he : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _GEN_133 = {{1'd0}, _heads_T_1}; // @[Mux.scala 27:73]
  wire [3:0] _heads_T_5 = _GEN_133 | _heads_T_2; // @[Mux.scala 27:73]
  wire [3:0] _heads_T_6 = _heads_T_5 | _heads_T_3; // @[Mux.scala 27:73]
  wire  _heads_T_7 = head == _heads_T_6; // @[InputUnit.scala 123:16]
  wire [2:0] _heads_T_10 = to_q_oh_2 ? 3'h5 : 3'h0; // @[Mux.scala 27:73]
  wire [3:0] _heads_T_11 = to_q_oh_3 ? 4'ha : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _GEN_134 = {{1'd0}, _heads_T_10}; // @[Mux.scala 27:73]
  wire [3:0] _heads_T_14 = _GEN_134 | _heads_T_11; // @[Mux.scala 27:73]
  wire [3:0] _heads_T_16 = head + 4'h1; // @[InputUnit.scala 125:16]
  wire  _GEN_71 = to_q_oh_0 | _GEN_51; // @[InputUnit.scala 127:29 128:32]
  wire [63:0] _GEN_75 = to_q_oh_0 ? mem_payload_qs_0_io_enq_bits_MPORT_data : io_enq_0_bits_payload; // @[InputUnit.scala 127:29 129:31]
  wire  _GEN_76 = to_q_oh_0 ? mem_tail_qs_0_io_enq_bits_MPORT_data : io_enq_0_bits_tail; // @[InputUnit.scala 127:29 129:31]
  wire  _GEN_77 = to_q_oh_0 ? mem_head_qs_0_io_enq_bits_MPORT_data : io_enq_0_bits_head; // @[InputUnit.scala 127:29 129:31]
  wire  _GEN_78 = to_q_oh_1 | _GEN_55; // @[InputUnit.scala 127:29 128:32]
  wire [63:0] _GEN_82 = to_q_oh_1 ? mem_payload_qs_1_io_enq_bits_MPORT_data : io_enq_0_bits_payload; // @[InputUnit.scala 127:29 129:31]
  wire  _GEN_83 = to_q_oh_1 ? mem_tail_qs_1_io_enq_bits_MPORT_data : io_enq_0_bits_tail; // @[InputUnit.scala 127:29 129:31]
  wire  _GEN_84 = to_q_oh_1 ? mem_head_qs_1_io_enq_bits_MPORT_data : io_enq_0_bits_head; // @[InputUnit.scala 127:29 129:31]
  wire  _GEN_85 = to_q_oh_2 | _GEN_59; // @[InputUnit.scala 127:29 128:32]
  wire [63:0] _GEN_89 = to_q_oh_2 ? mem_payload_qs_2_io_enq_bits_MPORT_data : io_enq_0_bits_payload; // @[InputUnit.scala 127:29 129:31]
  wire  _GEN_90 = to_q_oh_2 ? mem_tail_qs_2_io_enq_bits_MPORT_data : io_enq_0_bits_tail; // @[InputUnit.scala 127:29 129:31]
  wire  _GEN_91 = to_q_oh_2 ? mem_head_qs_2_io_enq_bits_MPORT_data : io_enq_0_bits_head; // @[InputUnit.scala 127:29 129:31]
  wire  _GEN_92 = to_q_oh_3 | _GEN_63; // @[InputUnit.scala 127:29 128:32]
  wire [63:0] _GEN_96 = to_q_oh_3 ? mem_payload_qs_3_io_enq_bits_MPORT_data : io_enq_0_bits_payload; // @[InputUnit.scala 127:29 129:31]
  wire  _GEN_97 = to_q_oh_3 ? mem_tail_qs_3_io_enq_bits_MPORT_data : io_enq_0_bits_tail; // @[InputUnit.scala 127:29 129:31]
  wire  _GEN_98 = to_q_oh_3 ? mem_head_qs_3_io_enq_bits_MPORT_data : io_enq_0_bits_head; // @[InputUnit.scala 127:29 129:31]
  Queue_4 qs_0 ( // @[InputUnit.scala 90:49]
    .clock(qs_0_clock),
    .reset(qs_0_reset),
    .io_enq_ready(qs_0_io_enq_ready),
    .io_enq_valid(qs_0_io_enq_valid),
    .io_enq_bits_head(qs_0_io_enq_bits_head),
    .io_enq_bits_tail(qs_0_io_enq_bits_tail),
    .io_enq_bits_payload(qs_0_io_enq_bits_payload),
    .io_deq_ready(qs_0_io_deq_ready),
    .io_deq_valid(qs_0_io_deq_valid),
    .io_deq_bits_head(qs_0_io_deq_bits_head),
    .io_deq_bits_tail(qs_0_io_deq_bits_tail),
    .io_deq_bits_payload(qs_0_io_deq_bits_payload)
  );
  Queue_4 qs_1 ( // @[InputUnit.scala 90:49]
    .clock(qs_1_clock),
    .reset(qs_1_reset),
    .io_enq_ready(qs_1_io_enq_ready),
    .io_enq_valid(qs_1_io_enq_valid),
    .io_enq_bits_head(qs_1_io_enq_bits_head),
    .io_enq_bits_tail(qs_1_io_enq_bits_tail),
    .io_enq_bits_payload(qs_1_io_enq_bits_payload),
    .io_deq_ready(qs_1_io_deq_ready),
    .io_deq_valid(qs_1_io_deq_valid),
    .io_deq_bits_head(qs_1_io_deq_bits_head),
    .io_deq_bits_tail(qs_1_io_deq_bits_tail),
    .io_deq_bits_payload(qs_1_io_deq_bits_payload)
  );
  Queue_4 qs_2 ( // @[InputUnit.scala 90:49]
    .clock(qs_2_clock),
    .reset(qs_2_reset),
    .io_enq_ready(qs_2_io_enq_ready),
    .io_enq_valid(qs_2_io_enq_valid),
    .io_enq_bits_head(qs_2_io_enq_bits_head),
    .io_enq_bits_tail(qs_2_io_enq_bits_tail),
    .io_enq_bits_payload(qs_2_io_enq_bits_payload),
    .io_deq_ready(qs_2_io_deq_ready),
    .io_deq_valid(qs_2_io_deq_valid),
    .io_deq_bits_head(qs_2_io_deq_bits_head),
    .io_deq_bits_tail(qs_2_io_deq_bits_tail),
    .io_deq_bits_payload(qs_2_io_deq_bits_payload)
  );
  Queue_4 qs_3 ( // @[InputUnit.scala 90:49]
    .clock(qs_3_clock),
    .reset(qs_3_reset),
    .io_enq_ready(qs_3_io_enq_ready),
    .io_enq_valid(qs_3_io_enq_valid),
    .io_enq_bits_head(qs_3_io_enq_bits_head),
    .io_enq_bits_tail(qs_3_io_enq_bits_tail),
    .io_enq_bits_payload(qs_3_io_enq_bits_payload),
    .io_deq_ready(qs_3_io_deq_ready),
    .io_deq_valid(qs_3_io_deq_valid),
    .io_deq_bits_head(qs_3_io_deq_bits_head),
    .io_deq_bits_tail(qs_3_io_deq_bits_tail),
    .io_deq_bits_payload(qs_3_io_deq_bits_payload)
  );
  assign mem_head_qs_0_io_enq_bits_MPORT_en = _T_9 & to_q_oh_0;
  assign mem_head_qs_0_io_enq_bits_MPORT_addr = _head_T_5 | _head_T_3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_head_qs_0_io_enq_bits_MPORT_data = mem_head[mem_head_qs_0_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `else
  assign mem_head_qs_0_io_enq_bits_MPORT_data = mem_head_qs_0_io_enq_bits_MPORT_addr >= 4'hf ? _RAND_1[0:0] :
    mem_head[mem_head_qs_0_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_head_qs_1_io_enq_bits_MPORT_en = _T_9 & to_q_oh_1;
  assign mem_head_qs_1_io_enq_bits_MPORT_addr = _head_T_5 | _head_T_3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_head_qs_1_io_enq_bits_MPORT_data = mem_head[mem_head_qs_1_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `else
  assign mem_head_qs_1_io_enq_bits_MPORT_data = mem_head_qs_1_io_enq_bits_MPORT_addr >= 4'hf ? _RAND_2[0:0] :
    mem_head[mem_head_qs_1_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_head_qs_2_io_enq_bits_MPORT_en = _T_9 & to_q_oh_2;
  assign mem_head_qs_2_io_enq_bits_MPORT_addr = _head_T_5 | _head_T_3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_head_qs_2_io_enq_bits_MPORT_data = mem_head[mem_head_qs_2_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `else
  assign mem_head_qs_2_io_enq_bits_MPORT_data = mem_head_qs_2_io_enq_bits_MPORT_addr >= 4'hf ? _RAND_3[0:0] :
    mem_head[mem_head_qs_2_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_head_qs_3_io_enq_bits_MPORT_en = _T_9 & to_q_oh_3;
  assign mem_head_qs_3_io_enq_bits_MPORT_addr = _head_T_5 | _head_T_3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_head_qs_3_io_enq_bits_MPORT_data = mem_head[mem_head_qs_3_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `else
  assign mem_head_qs_3_io_enq_bits_MPORT_data = mem_head_qs_3_io_enq_bits_MPORT_addr >= 4'hf ? _RAND_4[0:0] :
    mem_head[mem_head_qs_3_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_head_MPORT_data = io_enq_0_bits_head;
  assign mem_head_MPORT_addr = 2'h3 == io_enq_0_bits_virt_channel_id ? tails_3 : _GEN_2;
  assign mem_head_MPORT_mask = 1'h1;
  assign mem_head_MPORT_en = io_enq_0_valid & _T;
  assign mem_tail_qs_0_io_enq_bits_MPORT_en = _T_9 & to_q_oh_0;
  assign mem_tail_qs_0_io_enq_bits_MPORT_addr = _head_T_5 | _head_T_3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_tail_qs_0_io_enq_bits_MPORT_data = mem_tail[mem_tail_qs_0_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `else
  assign mem_tail_qs_0_io_enq_bits_MPORT_data = mem_tail_qs_0_io_enq_bits_MPORT_addr >= 4'hf ? _RAND_6[0:0] :
    mem_tail[mem_tail_qs_0_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_tail_qs_1_io_enq_bits_MPORT_en = _T_9 & to_q_oh_1;
  assign mem_tail_qs_1_io_enq_bits_MPORT_addr = _head_T_5 | _head_T_3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_tail_qs_1_io_enq_bits_MPORT_data = mem_tail[mem_tail_qs_1_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `else
  assign mem_tail_qs_1_io_enq_bits_MPORT_data = mem_tail_qs_1_io_enq_bits_MPORT_addr >= 4'hf ? _RAND_7[0:0] :
    mem_tail[mem_tail_qs_1_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_tail_qs_2_io_enq_bits_MPORT_en = _T_9 & to_q_oh_2;
  assign mem_tail_qs_2_io_enq_bits_MPORT_addr = _head_T_5 | _head_T_3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_tail_qs_2_io_enq_bits_MPORT_data = mem_tail[mem_tail_qs_2_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `else
  assign mem_tail_qs_2_io_enq_bits_MPORT_data = mem_tail_qs_2_io_enq_bits_MPORT_addr >= 4'hf ? _RAND_8[0:0] :
    mem_tail[mem_tail_qs_2_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_tail_qs_3_io_enq_bits_MPORT_en = _T_9 & to_q_oh_3;
  assign mem_tail_qs_3_io_enq_bits_MPORT_addr = _head_T_5 | _head_T_3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_tail_qs_3_io_enq_bits_MPORT_data = mem_tail[mem_tail_qs_3_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `else
  assign mem_tail_qs_3_io_enq_bits_MPORT_data = mem_tail_qs_3_io_enq_bits_MPORT_addr >= 4'hf ? _RAND_9[0:0] :
    mem_tail[mem_tail_qs_3_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_tail_MPORT_data = io_enq_0_bits_tail;
  assign mem_tail_MPORT_addr = 2'h3 == io_enq_0_bits_virt_channel_id ? tails_3 : _GEN_2;
  assign mem_tail_MPORT_mask = 1'h1;
  assign mem_tail_MPORT_en = io_enq_0_valid & _T;
  assign mem_payload_qs_0_io_enq_bits_MPORT_en = _T_9 & to_q_oh_0;
  assign mem_payload_qs_0_io_enq_bits_MPORT_addr = _head_T_5 | _head_T_3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_payload_qs_0_io_enq_bits_MPORT_data = mem_payload[mem_payload_qs_0_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `else
  assign mem_payload_qs_0_io_enq_bits_MPORT_data = mem_payload_qs_0_io_enq_bits_MPORT_addr >= 4'hf ? _RAND_11[63:0] :
    mem_payload[mem_payload_qs_0_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_payload_qs_1_io_enq_bits_MPORT_en = _T_9 & to_q_oh_1;
  assign mem_payload_qs_1_io_enq_bits_MPORT_addr = _head_T_5 | _head_T_3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_payload_qs_1_io_enq_bits_MPORT_data = mem_payload[mem_payload_qs_1_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `else
  assign mem_payload_qs_1_io_enq_bits_MPORT_data = mem_payload_qs_1_io_enq_bits_MPORT_addr >= 4'hf ? _RAND_12[63:0] :
    mem_payload[mem_payload_qs_1_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_payload_qs_2_io_enq_bits_MPORT_en = _T_9 & to_q_oh_2;
  assign mem_payload_qs_2_io_enq_bits_MPORT_addr = _head_T_5 | _head_T_3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_payload_qs_2_io_enq_bits_MPORT_data = mem_payload[mem_payload_qs_2_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `else
  assign mem_payload_qs_2_io_enq_bits_MPORT_data = mem_payload_qs_2_io_enq_bits_MPORT_addr >= 4'hf ? _RAND_13[63:0] :
    mem_payload[mem_payload_qs_2_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_payload_qs_3_io_enq_bits_MPORT_en = _T_9 & to_q_oh_3;
  assign mem_payload_qs_3_io_enq_bits_MPORT_addr = _head_T_5 | _head_T_3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_payload_qs_3_io_enq_bits_MPORT_data = mem_payload[mem_payload_qs_3_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `else
  assign mem_payload_qs_3_io_enq_bits_MPORT_data = mem_payload_qs_3_io_enq_bits_MPORT_addr >= 4'hf ? _RAND_14[63:0] :
    mem_payload[mem_payload_qs_3_io_enq_bits_MPORT_addr]; // @[InputUnit.scala 85:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_payload_MPORT_data = io_enq_0_bits_payload;
  assign mem_payload_MPORT_addr = 2'h3 == io_enq_0_bits_virt_channel_id ? tails_3 : _GEN_2;
  assign mem_payload_MPORT_mask = 1'h1;
  assign mem_payload_MPORT_en = io_enq_0_valid & _T;
  assign io_deq_0_bits_head = qs_0_io_deq_bits_head; // @[InputUnit.scala 134:19]
  assign io_deq_0_bits_tail = qs_0_io_deq_bits_tail; // @[InputUnit.scala 134:19]
  assign io_deq_0_bits_payload = qs_0_io_deq_bits_payload; // @[InputUnit.scala 134:19]
  assign io_deq_1_valid = qs_1_io_deq_valid; // @[InputUnit.scala 134:19]
  assign io_deq_1_bits_head = qs_1_io_deq_bits_head; // @[InputUnit.scala 134:19]
  assign io_deq_1_bits_tail = qs_1_io_deq_bits_tail; // @[InputUnit.scala 134:19]
  assign io_deq_1_bits_payload = qs_1_io_deq_bits_payload; // @[InputUnit.scala 134:19]
  assign io_deq_2_valid = qs_2_io_deq_valid; // @[InputUnit.scala 134:19]
  assign io_deq_2_bits_head = qs_2_io_deq_bits_head; // @[InputUnit.scala 134:19]
  assign io_deq_2_bits_tail = qs_2_io_deq_bits_tail; // @[InputUnit.scala 134:19]
  assign io_deq_2_bits_payload = qs_2_io_deq_bits_payload; // @[InputUnit.scala 134:19]
  assign io_deq_3_valid = qs_3_io_deq_valid; // @[InputUnit.scala 134:19]
  assign io_deq_3_bits_head = qs_3_io_deq_bits_head; // @[InputUnit.scala 134:19]
  assign io_deq_3_bits_tail = qs_3_io_deq_bits_tail; // @[InputUnit.scala 134:19]
  assign io_deq_3_bits_payload = qs_3_io_deq_bits_payload; // @[InputUnit.scala 134:19]
  assign qs_0_clock = clock;
  assign qs_0_reset = reset;
  assign qs_0_io_enq_valid = _T_9 ? _GEN_71 : _GEN_51; // @[InputUnit.scala 120:27]
  assign qs_0_io_enq_bits_head = _T_9 ? _GEN_77 : io_enq_0_bits_head; // @[InputUnit.scala 120:27]
  assign qs_0_io_enq_bits_tail = _T_9 ? _GEN_76 : io_enq_0_bits_tail; // @[InputUnit.scala 120:27]
  assign qs_0_io_enq_bits_payload = _T_9 ? _GEN_75 : io_enq_0_bits_payload; // @[InputUnit.scala 120:27]
  assign qs_0_io_deq_ready = 1'h0; // @[InputUnit.scala 134:19]
  assign qs_1_clock = clock;
  assign qs_1_reset = reset;
  assign qs_1_io_enq_valid = _T_9 ? _GEN_78 : _GEN_55; // @[InputUnit.scala 120:27]
  assign qs_1_io_enq_bits_head = _T_9 ? _GEN_84 : io_enq_0_bits_head; // @[InputUnit.scala 120:27]
  assign qs_1_io_enq_bits_tail = _T_9 ? _GEN_83 : io_enq_0_bits_tail; // @[InputUnit.scala 120:27]
  assign qs_1_io_enq_bits_payload = _T_9 ? _GEN_82 : io_enq_0_bits_payload; // @[InputUnit.scala 120:27]
  assign qs_1_io_deq_ready = io_deq_1_ready; // @[InputUnit.scala 134:19]
  assign qs_2_clock = clock;
  assign qs_2_reset = reset;
  assign qs_2_io_enq_valid = _T_9 ? _GEN_85 : _GEN_59; // @[InputUnit.scala 120:27]
  assign qs_2_io_enq_bits_head = _T_9 ? _GEN_91 : io_enq_0_bits_head; // @[InputUnit.scala 120:27]
  assign qs_2_io_enq_bits_tail = _T_9 ? _GEN_90 : io_enq_0_bits_tail; // @[InputUnit.scala 120:27]
  assign qs_2_io_enq_bits_payload = _T_9 ? _GEN_89 : io_enq_0_bits_payload; // @[InputUnit.scala 120:27]
  assign qs_2_io_deq_ready = io_deq_2_ready; // @[InputUnit.scala 134:19]
  assign qs_3_clock = clock;
  assign qs_3_reset = reset;
  assign qs_3_io_enq_valid = _T_9 ? _GEN_92 : _GEN_63; // @[InputUnit.scala 120:27]
  assign qs_3_io_enq_bits_head = _T_9 ? _GEN_98 : io_enq_0_bits_head; // @[InputUnit.scala 120:27]
  assign qs_3_io_enq_bits_tail = _T_9 ? _GEN_97 : io_enq_0_bits_tail; // @[InputUnit.scala 120:27]
  assign qs_3_io_enq_bits_payload = _T_9 ? _GEN_96 : io_enq_0_bits_payload; // @[InputUnit.scala 120:27]
  assign qs_3_io_deq_ready = io_deq_3_ready; // @[InputUnit.scala 134:19]
  always @(posedge clock) begin
    if (mem_head_MPORT_en & mem_head_MPORT_mask) begin
      mem_head[mem_head_MPORT_addr] <= mem_head_MPORT_data; // @[InputUnit.scala 85:18]
    end
    if (mem_tail_MPORT_en & mem_tail_MPORT_mask) begin
      mem_tail[mem_tail_MPORT_addr] <= mem_tail_MPORT_data; // @[InputUnit.scala 85:18]
    end
    if (mem_payload_MPORT_en & mem_payload_MPORT_mask) begin
      mem_payload[mem_payload_MPORT_addr] <= mem_payload_MPORT_data; // @[InputUnit.scala 85:18]
    end
    if (reset) begin // @[InputUnit.scala 86:24]
      heads_0 <= 4'h0; // @[InputUnit.scala 86:24]
    end else if (_T_9) begin // @[InputUnit.scala 120:27]
      if (2'h0 == to_q) begin // @[InputUnit.scala 122:21]
        if (_heads_T_7) begin // @[InputUnit.scala 122:27]
          heads_0 <= _heads_T_14;
        end else begin
          heads_0 <= _heads_T_16;
        end
      end
    end
    if (reset) begin // @[InputUnit.scala 86:24]
      heads_1 <= 4'h0; // @[InputUnit.scala 86:24]
    end else if (_T_9) begin // @[InputUnit.scala 120:27]
      if (2'h1 == to_q) begin // @[InputUnit.scala 122:21]
        if (_heads_T_7) begin // @[InputUnit.scala 122:27]
          heads_1 <= _heads_T_14;
        end else begin
          heads_1 <= _heads_T_16;
        end
      end
    end
    if (reset) begin // @[InputUnit.scala 86:24]
      heads_2 <= 4'h5; // @[InputUnit.scala 86:24]
    end else if (_T_9) begin // @[InputUnit.scala 120:27]
      if (2'h2 == to_q) begin // @[InputUnit.scala 122:21]
        if (_heads_T_7) begin // @[InputUnit.scala 122:27]
          heads_2 <= _heads_T_14;
        end else begin
          heads_2 <= _heads_T_16;
        end
      end
    end
    if (reset) begin // @[InputUnit.scala 86:24]
      heads_3 <= 4'ha; // @[InputUnit.scala 86:24]
    end else if (_T_9) begin // @[InputUnit.scala 120:27]
      if (2'h3 == to_q) begin // @[InputUnit.scala 122:21]
        if (_heads_T_7) begin // @[InputUnit.scala 122:27]
          heads_3 <= _heads_T_14;
        end else begin
          heads_3 <= _heads_T_16;
        end
      end
    end
    if (reset) begin // @[InputUnit.scala 87:24]
      tails_0 <= 4'h0; // @[InputUnit.scala 87:24]
    end else if (io_enq_0_valid & ~direct_to_q) begin // @[InputUnit.scala 100:44]
      if (2'h0 == io_enq_0_bits_virt_channel_id) begin // @[InputUnit.scala 103:45]
        if (_tails_T_11) begin // @[InputUnit.scala 103:51]
          tails_0 <= _tails_T_22;
        end else begin
          tails_0 <= _tails_T_24;
        end
      end
    end
    if (reset) begin // @[InputUnit.scala 87:24]
      tails_1 <= 4'h0; // @[InputUnit.scala 87:24]
    end else if (io_enq_0_valid & ~direct_to_q) begin // @[InputUnit.scala 100:44]
      if (2'h1 == io_enq_0_bits_virt_channel_id) begin // @[InputUnit.scala 103:45]
        if (_tails_T_11) begin // @[InputUnit.scala 103:51]
          tails_1 <= _tails_T_22;
        end else begin
          tails_1 <= _tails_T_24;
        end
      end
    end
    if (reset) begin // @[InputUnit.scala 87:24]
      tails_2 <= 4'h5; // @[InputUnit.scala 87:24]
    end else if (io_enq_0_valid & ~direct_to_q) begin // @[InputUnit.scala 100:44]
      if (2'h2 == io_enq_0_bits_virt_channel_id) begin // @[InputUnit.scala 103:45]
        if (_tails_T_11) begin // @[InputUnit.scala 103:51]
          tails_2 <= _tails_T_22;
        end else begin
          tails_2 <= _tails_T_24;
        end
      end
    end
    if (reset) begin // @[InputUnit.scala 87:24]
      tails_3 <= 4'ha; // @[InputUnit.scala 87:24]
    end else if (io_enq_0_valid & ~direct_to_q) begin // @[InputUnit.scala 100:44]
      if (2'h3 == io_enq_0_bits_virt_channel_id) begin // @[InputUnit.scala 103:45]
        if (_tails_T_11) begin // @[InputUnit.scala 103:51]
          tails_3 <= _tails_T_22;
        end else begin
          tails_3 <= _tails_T_24;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {1{`RANDOM}};
  _RAND_2 = {1{`RANDOM}};
  _RAND_3 = {1{`RANDOM}};
  _RAND_4 = {1{`RANDOM}};
  _RAND_6 = {1{`RANDOM}};
  _RAND_7 = {1{`RANDOM}};
  _RAND_8 = {1{`RANDOM}};
  _RAND_9 = {1{`RANDOM}};
  _RAND_11 = {2{`RANDOM}};
  _RAND_12 = {2{`RANDOM}};
  _RAND_13 = {2{`RANDOM}};
  _RAND_14 = {2{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 15; initvar = initvar+1)
    mem_head[initvar] = _RAND_0[0:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 15; initvar = initvar+1)
    mem_tail[initvar] = _RAND_5[0:0];
  _RAND_10 = {2{`RANDOM}};
  for (initvar = 0; initvar < 15; initvar = initvar+1)
    mem_payload[initvar] = _RAND_10[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  heads_0 = _RAND_15[3:0];
  _RAND_16 = {1{`RANDOM}};
  heads_1 = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  heads_2 = _RAND_17[3:0];
  _RAND_18 = {1{`RANDOM}};
  heads_3 = _RAND_18[3:0];
  _RAND_19 = {1{`RANDOM}};
  tails_0 = _RAND_19[3:0];
  _RAND_20 = {1{`RANDOM}};
  tails_1 = _RAND_20[3:0];
  _RAND_21 = {1{`RANDOM}};
  tails_2 = _RAND_21[3:0];
  _RAND_22 = {1{`RANDOM}};
  tails_3 = _RAND_22[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Arbiter(
  input        io_in_1_valid,
  output       io_in_2_ready,
  input        io_in_2_valid,
  output       io_in_3_ready,
  input        io_in_3_valid,
  output       io_out_valid,
  output [1:0] io_out_bits_src_virt_id
);
  wire [1:0] _GEN_0 = io_in_2_valid ? 2'h2 : 2'h3; // @[Arbiter.scala 135:13 138:26 139:17]
  wire  grant_3 = ~(io_in_1_valid | io_in_2_valid); // @[Arbiter.scala 45:78]
  assign io_in_2_ready = ~io_in_1_valid; // @[Arbiter.scala 45:78]
  assign io_in_3_ready = ~(io_in_1_valid | io_in_2_valid); // @[Arbiter.scala 45:78]
  assign io_out_valid = ~grant_3 | io_in_3_valid; // @[Arbiter.scala 147:31]
  assign io_out_bits_src_virt_id = io_in_1_valid ? 2'h1 : _GEN_0; // @[Arbiter.scala 138:26 140:19]
endmodule
module SwitchArbiter_2(
  input        clock,
  input        reset,
  output       io_in_0_ready,
  input        io_in_0_valid,
  output       io_in_1_ready,
  input        io_in_1_valid,
  input        io_in_1_bits_vc_sel_0_0,
  input        io_in_1_bits_tail,
  output       io_in_2_ready,
  input        io_in_2_valid,
  input        io_in_2_bits_vc_sel_0_0,
  input        io_in_2_bits_tail,
  output       io_in_3_ready,
  input        io_in_3_valid,
  input        io_in_3_bits_vc_sel_0_0,
  input        io_in_3_bits_tail,
  input        io_out_0_ready,
  output       io_out_0_valid,
  output       io_out_0_bits_vc_sel_0_0,
  output       io_out_0_bits_tail,
  output [3:0] io_chosen_oh_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] lock_0; // @[SwitchAllocator.scala 24:38]
  wire [3:0] _unassigned_T = {io_in_3_valid,io_in_2_valid,io_in_1_valid,1'h0}; // @[Cat.scala 33:92]
  wire [3:0] _unassigned_T_1 = ~lock_0; // @[SwitchAllocator.scala 25:54]
  wire [3:0] unassigned = _unassigned_T & _unassigned_T_1; // @[SwitchAllocator.scala 25:52]
  reg [3:0] mask; // @[SwitchAllocator.scala 27:21]
  wire [3:0] _GEN_6 = {{3'd0}, mask == 4'h0}; // @[SwitchAllocator.scala 30:58]
  wire [3:0] _sel_T_1 = unassigned & _GEN_6; // @[SwitchAllocator.scala 30:58]
  wire [7:0] _sel_T_2 = {unassigned,_sel_T_1}; // @[Cat.scala 33:92]
  wire [7:0] _sel_T_11 = _sel_T_2[7] ? 8'h80 : 8'h0; // @[Mux.scala 47:70]
  wire [7:0] _sel_T_12 = _sel_T_2[6] ? 8'h40 : _sel_T_11; // @[Mux.scala 47:70]
  wire [7:0] _sel_T_13 = _sel_T_2[5] ? 8'h20 : _sel_T_12; // @[Mux.scala 47:70]
  wire [7:0] _sel_T_14 = _sel_T_2[4] ? 8'h10 : _sel_T_13; // @[Mux.scala 47:70]
  wire [7:0] _sel_T_15 = _sel_T_2[3] ? 8'h8 : _sel_T_14; // @[Mux.scala 47:70]
  wire [7:0] _sel_T_16 = _sel_T_2[2] ? 8'h4 : _sel_T_15; // @[Mux.scala 47:70]
  wire [7:0] _sel_T_17 = _sel_T_2[1] ? 8'h2 : _sel_T_16; // @[Mux.scala 47:70]
  wire [7:0] sel = _sel_T_2[0] ? 8'h1 : _sel_T_17; // @[Mux.scala 47:70]
  wire [7:0] _GEN_7 = {{4'd0}, sel[7:4]}; // @[SwitchAllocator.scala 32:23]
  wire [7:0] _choices_0_T_1 = sel | _GEN_7; // @[SwitchAllocator.scala 32:23]
  wire [3:0] choices_0 = _choices_0_T_1[3:0]; // @[SwitchAllocator.scala 28:21 32:16]
  wire [3:0] in_tails = {io_in_3_bits_tail,io_in_2_bits_tail,io_in_1_bits_tail,1'h0}; // @[Cat.scala 33:92]
  wire [3:0] _chosen_T = _unassigned_T & lock_0; // @[SwitchAllocator.scala 42:33]
  wire [3:0] chosen = |_chosen_T ? lock_0 : choices_0; // @[SwitchAllocator.scala 42:21]
  wire [3:0] _io_out_0_valid_T = _unassigned_T & chosen; // @[SwitchAllocator.scala 44:35]
  wire  _T_17 = io_out_0_ready & io_out_0_valid; // @[Decoupled.scala 51:35]
  wire [3:0] _lock_0_T = ~in_tails; // @[SwitchAllocator.scala 53:27]
  wire [3:0] _lock_0_T_1 = chosen & _lock_0_T; // @[SwitchAllocator.scala 53:25]
  wire [3:0] _GEN_8 = {{1'd0}, io_chosen_oh_0[3:1]}; // @[SwitchAllocator.scala 58:71]
  wire [3:0] _mask_T_4 = io_chosen_oh_0 | _GEN_8; // @[SwitchAllocator.scala 58:71]
  wire [3:0] _GEN_9 = {{2'd0}, io_chosen_oh_0[3:2]}; // @[SwitchAllocator.scala 58:71]
  wire [3:0] _mask_T_5 = _mask_T_4 | _GEN_9; // @[SwitchAllocator.scala 58:71]
  wire [3:0] _GEN_10 = {{3'd0}, io_chosen_oh_0[3]}; // @[SwitchAllocator.scala 58:71]
  wire [3:0] _mask_T_6 = _mask_T_5 | _GEN_10; // @[SwitchAllocator.scala 58:71]
  wire [3:0] _mask_T_7 = ~mask; // @[SwitchAllocator.scala 60:17]
  wire [4:0] _mask_T_9 = {mask, 1'h0}; // @[SwitchAllocator.scala 60:43]
  wire [4:0] _mask_T_10 = _mask_T_9 | 5'h1; // @[SwitchAllocator.scala 60:49]
  wire [4:0] _mask_T_11 = _mask_T_7 == 4'h0 ? 5'h0 : _mask_T_10; // @[SwitchAllocator.scala 60:16]
  wire [4:0] _GEN_5 = _T_17 ? {{1'd0}, _mask_T_6} : _mask_T_11; // @[SwitchAllocator.scala 57:27 58:10 60:10]
  wire [4:0] _GEN_11 = reset ? 5'h0 : _GEN_5; // @[SwitchAllocator.scala 27:{21,21}]
  assign io_in_0_ready = chosen[0] & io_out_0_ready; // @[SwitchAllocator.scala 47:23]
  assign io_in_1_ready = chosen[1] & io_out_0_ready; // @[SwitchAllocator.scala 47:23]
  assign io_in_2_ready = chosen[2] & io_out_0_ready; // @[SwitchAllocator.scala 47:23]
  assign io_in_3_ready = chosen[3] & io_out_0_ready; // @[SwitchAllocator.scala 47:23]
  assign io_out_0_valid = |_io_out_0_valid_T; // @[SwitchAllocator.scala 44:45]
  assign io_out_0_bits_vc_sel_0_0 = chosen[1] & io_in_1_bits_vc_sel_0_0 | chosen[2] & io_in_2_bits_vc_sel_0_0 | chosen[3
    ] & io_in_3_bits_vc_sel_0_0; // @[Mux.scala 27:73]
  assign io_out_0_bits_tail = chosen[1] & io_in_1_bits_tail | chosen[2] & io_in_2_bits_tail | chosen[3] &
    io_in_3_bits_tail; // @[Mux.scala 27:73]
  assign io_chosen_oh_0 = |_chosen_T ? lock_0 : choices_0; // @[SwitchAllocator.scala 42:21]
  always @(posedge clock) begin
    if (reset) begin // @[SwitchAllocator.scala 24:38]
      lock_0 <= 4'h0; // @[SwitchAllocator.scala 24:38]
    end else if (_T_17) begin // @[SwitchAllocator.scala 52:29]
      lock_0 <= _lock_0_T_1; // @[SwitchAllocator.scala 53:15]
    end
    mask <= _GEN_11[3:0]; // @[SwitchAllocator.scala 27:{21,21}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lock_0 = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  mask = _RAND_1[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module InputUnit(
  input         clock,
  input         reset,
  output        io_router_req_valid,
  output [1:0]  io_router_req_bits_src_virt_id,
  input         io_vcalloc_req_ready,
  output        io_vcalloc_req_valid,
  output        io_vcalloc_req_bits_vc_sel_0_0,
  input         io_vcalloc_resp_vc_sel_0_0,
  input         io_out_credit_available_0_0,
  input         io_salloc_req_0_ready,
  output        io_salloc_req_0_valid,
  output        io_salloc_req_0_bits_vc_sel_0_0,
  output        io_salloc_req_0_bits_tail,
  output        io_out_0_valid,
  output        io_out_0_bits_flit_head,
  output        io_out_0_bits_flit_tail,
  output [63:0] io_out_0_bits_flit_payload,
  output [1:0]  io_out_0_bits_flit_flow_ingress_node,
  output [1:0]  io_debug_va_stall,
  output [1:0]  io_debug_sa_stall,
  input         io_in_flit_0_valid,
  input         io_in_flit_0_bits_head,
  input         io_in_flit_0_bits_tail,
  input  [63:0] io_in_flit_0_bits_payload,
  input  [1:0]  io_in_flit_0_bits_flow_ingress_node,
  input  [1:0]  io_in_flit_0_bits_flow_egress_node,
  input  [1:0]  io_in_flit_0_bits_virt_channel_id,
  output [3:0]  io_in_credit_return,
  output [3:0]  io_in_vc_free
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
`endif // RANDOMIZE_REG_INIT
  wire  input_buffer_clock; // @[InputUnit.scala 180:28]
  wire  input_buffer_reset; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_enq_0_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_enq_0_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_enq_0_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_enq_0_bits_payload; // @[InputUnit.scala 180:28]
  wire [1:0] input_buffer_io_enq_0_bits_virt_channel_id; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_0_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_0_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_deq_0_bits_payload; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_ready; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_deq_1_bits_payload; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_ready; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_deq_2_bits_payload; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_3_ready; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_3_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_3_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_3_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_deq_3_bits_payload; // @[InputUnit.scala 180:28]
  wire  route_arbiter_io_in_1_valid; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_2_ready; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_2_valid; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_3_ready; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_3_valid; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_out_valid; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_out_bits_src_virt_id; // @[InputUnit.scala 186:29]
  wire  salloc_arb_clock; // @[InputUnit.scala 279:26]
  wire  salloc_arb_reset; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_tail; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_tail; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_tail; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_tail; // @[InputUnit.scala 279:26]
  wire [3:0] salloc_arb_io_chosen_oh_0; // @[InputUnit.scala 279:26]
  reg [2:0] states_1_g; // @[InputUnit.scala 191:19]
  reg  states_1_vc_sel_0_0; // @[InputUnit.scala 191:19]
  reg [1:0] states_1_flow_ingress_node; // @[InputUnit.scala 191:19]
  reg [2:0] states_2_g; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_0_0; // @[InputUnit.scala 191:19]
  reg [1:0] states_2_flow_ingress_node; // @[InputUnit.scala 191:19]
  reg [2:0] states_3_g; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_0_0; // @[InputUnit.scala 191:19]
  reg [1:0] states_3_flow_ingress_node; // @[InputUnit.scala 191:19]
  wire  _T = io_in_flit_0_valid & io_in_flit_0_bits_head; // @[InputUnit.scala 194:32]
  wire  _T_3 = ~reset; // @[InputUnit.scala 196:13]
  wire [2:0] _GEN_1 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? states_1_g : 3'h0; // @[InputUnit.scala 197:{27,27}]
  wire [2:0] _GEN_2 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? states_2_g : _GEN_1; // @[InputUnit.scala 197:{27,27}]
  wire [2:0] _GEN_3 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? states_3_g : _GEN_2; // @[InputUnit.scala 197:{27,27}]
  wire  at_dest = io_in_flit_0_bits_flow_egress_node == 2'h1; // @[InputUnit.scala 198:57]
  wire [2:0] _states_g_T = at_dest ? 3'h2 : 3'h1; // @[InputUnit.scala 199:26]
  wire [2:0] _GEN_5 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? _states_g_T : states_1_g; // @[InputUnit.scala 191:19 199:{20,20}]
  wire [2:0] _GEN_6 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? _states_g_T : states_2_g; // @[InputUnit.scala 191:19 199:{20,20}]
  wire [2:0] _GEN_7 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? _states_g_T : states_3_g; // @[InputUnit.scala 191:19 199:{20,20}]
  wire  _GEN_9 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_1_vc_sel_0_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_10 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_0_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_11 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_0_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_13 = 2'h1 == io_in_flit_0_bits_virt_channel_id | _GEN_9; // @[InputUnit.scala 203:{44,44}]
  wire  _GEN_14 = 2'h2 == io_in_flit_0_bits_virt_channel_id | _GEN_10; // @[InputUnit.scala 203:{44,44}]
  wire  _GEN_15 = 2'h3 == io_in_flit_0_bits_virt_channel_id | _GEN_11; // @[InputUnit.scala 203:{44,44}]
  wire [2:0] _GEN_41 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_5 : states_1_g; // @[InputUnit.scala 191:19 194:60]
  wire [2:0] _GEN_42 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_6 : states_2_g; // @[InputUnit.scala 191:19 194:60]
  wire [2:0] _GEN_43 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_7 : states_3_g; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_45 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_13 : states_1_vc_sel_0_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_46 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_14 : states_2_vc_sel_0_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_47 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_15 : states_3_vc_sel_0_0; // @[InputUnit.scala 191:19 194:60]
  wire  _T_10 = route_arbiter_io_in_1_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_68 = _T_10 ? 3'h2 : _GEN_41; // @[InputUnit.scala 215:{23,29}]
  wire  _T_11 = route_arbiter_io_in_2_ready & route_arbiter_io_in_2_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_69 = _T_11 ? 3'h2 : _GEN_42; // @[InputUnit.scala 215:{23,29}]
  wire  _T_12 = route_arbiter_io_in_3_ready & route_arbiter_io_in_3_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_70 = _T_12 ? 3'h2 : _GEN_43; // @[InputUnit.scala 215:{23,29}]
  wire [2:0] _GEN_72 = 2'h1 == io_router_req_bits_src_virt_id ? states_1_g : 3'h0; // @[InputUnit.scala 224:{25,25}]
  wire [2:0] _GEN_73 = 2'h2 == io_router_req_bits_src_virt_id ? states_2_g : _GEN_72; // @[InputUnit.scala 224:{25,25}]
  wire [2:0] _GEN_74 = 2'h3 == io_router_req_bits_src_virt_id ? states_3_g : _GEN_73; // @[InputUnit.scala 224:{25,25}]
  wire [2:0] _GEN_76 = 2'h1 == io_router_req_bits_src_virt_id ? 3'h2 : _GEN_68; // @[InputUnit.scala 225:{18,18}]
  wire [2:0] _GEN_77 = 2'h2 == io_router_req_bits_src_virt_id ? 3'h2 : _GEN_69; // @[InputUnit.scala 225:{18,18}]
  wire [2:0] _GEN_78 = 2'h3 == io_router_req_bits_src_virt_id ? 3'h2 : _GEN_70; // @[InputUnit.scala 225:{18,18}]
  wire  _GEN_80 = 2'h1 == io_router_req_bits_src_virt_id ? 1'h0 : _GEN_45; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_81 = 2'h2 == io_router_req_bits_src_virt_id ? 1'h0 : _GEN_46; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_82 = 2'h3 == io_router_req_bits_src_virt_id ? 1'h0 : _GEN_47; // @[InputUnit.scala 227:25 228:26]
  wire [2:0] _GEN_84 = io_router_req_valid ? _GEN_76 : _GEN_68; // @[InputUnit.scala 222:31]
  wire [2:0] _GEN_85 = io_router_req_valid ? _GEN_77 : _GEN_69; // @[InputUnit.scala 222:31]
  wire [2:0] _GEN_86 = io_router_req_valid ? _GEN_78 : _GEN_70; // @[InputUnit.scala 222:31]
  wire  _GEN_88 = io_router_req_valid ? _GEN_80 : _GEN_45; // @[InputUnit.scala 222:31]
  wire  _GEN_89 = io_router_req_valid ? _GEN_81 : _GEN_46; // @[InputUnit.scala 222:31]
  wire  _GEN_90 = io_router_req_valid ? _GEN_82 : _GEN_47; // @[InputUnit.scala 222:31]
  reg [3:0] mask; // @[InputUnit.scala 233:21]
  wire  vcalloc_vals_1 = states_1_g == 3'h2; // @[InputUnit.scala 249:32]
  wire  vcalloc_vals_3 = states_3_g == 3'h2; // @[InputUnit.scala 249:32]
  wire  vcalloc_vals_2 = states_2_g == 3'h2; // @[InputUnit.scala 249:32]
  wire [3:0] _vcalloc_filter_T = {vcalloc_vals_3,vcalloc_vals_2,vcalloc_vals_1,1'h0}; // @[InputUnit.scala 236:59]
  wire [3:0] _vcalloc_filter_T_2 = ~mask; // @[InputUnit.scala 236:89]
  wire [3:0] _vcalloc_filter_T_3 = _vcalloc_filter_T & _vcalloc_filter_T_2; // @[InputUnit.scala 236:87]
  wire [7:0] _vcalloc_filter_T_4 = {vcalloc_vals_3,vcalloc_vals_2,vcalloc_vals_1,1'h0,_vcalloc_filter_T_3}; // @[Cat.scala 33:92]
  wire [7:0] _vcalloc_filter_T_13 = _vcalloc_filter_T_4[7] ? 8'h80 : 8'h0; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_14 = _vcalloc_filter_T_4[6] ? 8'h40 : _vcalloc_filter_T_13; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_15 = _vcalloc_filter_T_4[5] ? 8'h20 : _vcalloc_filter_T_14; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_16 = _vcalloc_filter_T_4[4] ? 8'h10 : _vcalloc_filter_T_15; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_17 = _vcalloc_filter_T_4[3] ? 8'h8 : _vcalloc_filter_T_16; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_18 = _vcalloc_filter_T_4[2] ? 8'h4 : _vcalloc_filter_T_17; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_19 = _vcalloc_filter_T_4[1] ? 8'h2 : _vcalloc_filter_T_18; // @[Mux.scala 47:70]
  wire [7:0] vcalloc_filter = _vcalloc_filter_T_4[0] ? 8'h1 : _vcalloc_filter_T_19; // @[Mux.scala 47:70]
  wire [3:0] vcalloc_sel = vcalloc_filter[3:0] | vcalloc_filter[7:4]; // @[InputUnit.scala 237:58]
  wire [3:0] _mask_T = 4'h1 << io_router_req_bits_src_virt_id; // @[InputUnit.scala 240:18]
  wire [3:0] _mask_T_2 = _mask_T - 4'h1; // @[InputUnit.scala 240:53]
  wire  _T_25 = vcalloc_vals_1 | vcalloc_vals_2 | vcalloc_vals_3; // @[package.scala 73:59]
  wire [1:0] _mask_T_12 = vcalloc_sel[1] ? 2'h3 : 2'h0; // @[Mux.scala 27:73]
  wire [2:0] _mask_T_13 = vcalloc_sel[2] ? 3'h7 : 3'h0; // @[Mux.scala 27:73]
  wire [3:0] _mask_T_14 = vcalloc_sel[3] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [1:0] _GEN_23 = {{1'd0}, vcalloc_sel[0]}; // @[Mux.scala 27:73]
  wire [1:0] _mask_T_15 = _GEN_23 | _mask_T_12; // @[Mux.scala 27:73]
  wire [2:0] _GEN_28 = {{1'd0}, _mask_T_15}; // @[Mux.scala 27:73]
  wire [2:0] _mask_T_16 = _GEN_28 | _mask_T_13; // @[Mux.scala 27:73]
  wire [3:0] _GEN_29 = {{1'd0}, _mask_T_16}; // @[Mux.scala 27:73]
  wire [3:0] _mask_T_17 = _GEN_29 | _mask_T_14; // @[Mux.scala 27:73]
  wire [2:0] _GEN_93 = vcalloc_vals_1 & vcalloc_sel[1] & io_vcalloc_req_ready ? 3'h3 : _GEN_84; // @[InputUnit.scala 253:{76,82}]
  wire [2:0] _GEN_94 = vcalloc_vals_2 & vcalloc_sel[2] & io_vcalloc_req_ready ? 3'h3 : _GEN_85; // @[InputUnit.scala 253:{76,82}]
  wire [2:0] _GEN_95 = vcalloc_vals_3 & vcalloc_sel[3] & io_vcalloc_req_ready ? 3'h3 : _GEN_86; // @[InputUnit.scala 253:{76,82}]
  wire [1:0] _io_debug_va_stall_T = {{1'd0}, vcalloc_vals_1}; // @[Bitwise.scala 51:90]
  wire [1:0] _io_debug_va_stall_T_2 = vcalloc_vals_2 + vcalloc_vals_3; // @[Bitwise.scala 51:90]
  wire [2:0] _io_debug_va_stall_T_4 = _io_debug_va_stall_T + _io_debug_va_stall_T_2; // @[Bitwise.scala 51:90]
  wire [2:0] _GEN_30 = {{2'd0}, io_vcalloc_req_ready}; // @[InputUnit.scala 266:47]
  wire [2:0] _io_debug_va_stall_T_7 = _io_debug_va_stall_T_4 - _GEN_30; // @[InputUnit.scala 266:47]
  wire  _T_35 = io_vcalloc_req_ready & io_vcalloc_req_valid; // @[Decoupled.scala 51:35]
  wire  credit_available = states_1_vc_sel_0_0 & io_out_credit_available_0_0; // @[InputUnit.scala 287:47]
  wire  _T_56 = salloc_arb_io_in_1_ready & salloc_arb_io_in_1_valid; // @[Decoupled.scala 51:35]
  wire  credit_available_1 = states_2_vc_sel_0_0 & io_out_credit_available_0_0; // @[InputUnit.scala 287:47]
  wire  _T_58 = salloc_arb_io_in_2_ready & salloc_arb_io_in_2_valid; // @[Decoupled.scala 51:35]
  wire  credit_available_2 = states_3_vc_sel_0_0 & io_out_credit_available_0_0; // @[InputUnit.scala 287:47]
  wire  _T_60 = salloc_arb_io_in_3_ready & salloc_arb_io_in_3_valid; // @[Decoupled.scala 51:35]
  wire  _io_debug_sa_stall_T_1 = salloc_arb_io_in_0_valid & ~salloc_arb_io_in_0_ready; // @[InputUnit.scala 301:67]
  wire  _io_debug_sa_stall_T_3 = salloc_arb_io_in_1_valid & ~salloc_arb_io_in_1_ready; // @[InputUnit.scala 301:67]
  wire  _io_debug_sa_stall_T_5 = salloc_arb_io_in_2_valid & ~salloc_arb_io_in_2_ready; // @[InputUnit.scala 301:67]
  wire  _io_debug_sa_stall_T_7 = salloc_arb_io_in_3_valid & ~salloc_arb_io_in_3_ready; // @[InputUnit.scala 301:67]
  wire [1:0] _io_debug_sa_stall_T_8 = _io_debug_sa_stall_T_1 + _io_debug_sa_stall_T_3; // @[Bitwise.scala 51:90]
  wire [1:0] _io_debug_sa_stall_T_10 = _io_debug_sa_stall_T_5 + _io_debug_sa_stall_T_7; // @[Bitwise.scala 51:90]
  wire [2:0] _io_debug_sa_stall_T_12 = _io_debug_sa_stall_T_8 + _io_debug_sa_stall_T_10; // @[Bitwise.scala 51:90]
  reg  salloc_outs_0_valid; // @[InputUnit.scala 318:8]
  reg  salloc_outs_0_flit_head; // @[InputUnit.scala 318:8]
  reg  salloc_outs_0_flit_tail; // @[InputUnit.scala 318:8]
  reg [63:0] salloc_outs_0_flit_payload; // @[InputUnit.scala 318:8]
  reg [1:0] salloc_outs_0_flit_flow_ingress_node; // @[InputUnit.scala 318:8]
  wire  _io_in_credit_return_T = salloc_arb_io_out_0_ready & salloc_arb_io_out_0_valid; // @[Decoupled.scala 51:35]
  wire  _io_in_vc_free_T_11 = salloc_arb_io_chosen_oh_0[0] & input_buffer_io_deq_0_bits_tail | salloc_arb_io_chosen_oh_0
    [1] & input_buffer_io_deq_1_bits_tail | salloc_arb_io_chosen_oh_0[2] & input_buffer_io_deq_2_bits_tail |
    salloc_arb_io_chosen_oh_0[3] & input_buffer_io_deq_3_bits_tail; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_4 = salloc_arb_io_chosen_oh_0[0] ? input_buffer_io_deq_0_bits_payload : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_5 = salloc_arb_io_chosen_oh_0[1] ? input_buffer_io_deq_1_bits_payload : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_6 = salloc_arb_io_chosen_oh_0[2] ? input_buffer_io_deq_2_bits_payload : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_7 = salloc_arb_io_chosen_oh_0[3] ? input_buffer_io_deq_3_bits_payload : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_8 = _salloc_outs_0_flit_payload_T_4 | _salloc_outs_0_flit_payload_T_5; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_9 = _salloc_outs_0_flit_payload_T_8 | _salloc_outs_0_flit_payload_T_6; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_26 = salloc_arb_io_chosen_oh_0[1] ? states_1_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_27 = salloc_arb_io_chosen_oh_0[2] ? states_2_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_28 = salloc_arb_io_chosen_oh_0[3] ? states_3_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_30 = _salloc_outs_0_flit_flow_T_26 | _salloc_outs_0_flit_flow_T_27; // @[Mux.scala 27:73]
  InputBuffer input_buffer ( // @[InputUnit.scala 180:28]
    .clock(input_buffer_clock),
    .reset(input_buffer_reset),
    .io_enq_0_valid(input_buffer_io_enq_0_valid),
    .io_enq_0_bits_head(input_buffer_io_enq_0_bits_head),
    .io_enq_0_bits_tail(input_buffer_io_enq_0_bits_tail),
    .io_enq_0_bits_payload(input_buffer_io_enq_0_bits_payload),
    .io_enq_0_bits_virt_channel_id(input_buffer_io_enq_0_bits_virt_channel_id),
    .io_deq_0_bits_head(input_buffer_io_deq_0_bits_head),
    .io_deq_0_bits_tail(input_buffer_io_deq_0_bits_tail),
    .io_deq_0_bits_payload(input_buffer_io_deq_0_bits_payload),
    .io_deq_1_ready(input_buffer_io_deq_1_ready),
    .io_deq_1_valid(input_buffer_io_deq_1_valid),
    .io_deq_1_bits_head(input_buffer_io_deq_1_bits_head),
    .io_deq_1_bits_tail(input_buffer_io_deq_1_bits_tail),
    .io_deq_1_bits_payload(input_buffer_io_deq_1_bits_payload),
    .io_deq_2_ready(input_buffer_io_deq_2_ready),
    .io_deq_2_valid(input_buffer_io_deq_2_valid),
    .io_deq_2_bits_head(input_buffer_io_deq_2_bits_head),
    .io_deq_2_bits_tail(input_buffer_io_deq_2_bits_tail),
    .io_deq_2_bits_payload(input_buffer_io_deq_2_bits_payload),
    .io_deq_3_ready(input_buffer_io_deq_3_ready),
    .io_deq_3_valid(input_buffer_io_deq_3_valid),
    .io_deq_3_bits_head(input_buffer_io_deq_3_bits_head),
    .io_deq_3_bits_tail(input_buffer_io_deq_3_bits_tail),
    .io_deq_3_bits_payload(input_buffer_io_deq_3_bits_payload)
  );
  Arbiter route_arbiter ( // @[InputUnit.scala 186:29]
    .io_in_1_valid(route_arbiter_io_in_1_valid),
    .io_in_2_ready(route_arbiter_io_in_2_ready),
    .io_in_2_valid(route_arbiter_io_in_2_valid),
    .io_in_3_ready(route_arbiter_io_in_3_ready),
    .io_in_3_valid(route_arbiter_io_in_3_valid),
    .io_out_valid(route_arbiter_io_out_valid),
    .io_out_bits_src_virt_id(route_arbiter_io_out_bits_src_virt_id)
  );
  SwitchArbiter_2 salloc_arb ( // @[InputUnit.scala 279:26]
    .clock(salloc_arb_clock),
    .reset(salloc_arb_reset),
    .io_in_0_ready(salloc_arb_io_in_0_ready),
    .io_in_0_valid(salloc_arb_io_in_0_valid),
    .io_in_1_ready(salloc_arb_io_in_1_ready),
    .io_in_1_valid(salloc_arb_io_in_1_valid),
    .io_in_1_bits_vc_sel_0_0(salloc_arb_io_in_1_bits_vc_sel_0_0),
    .io_in_1_bits_tail(salloc_arb_io_in_1_bits_tail),
    .io_in_2_ready(salloc_arb_io_in_2_ready),
    .io_in_2_valid(salloc_arb_io_in_2_valid),
    .io_in_2_bits_vc_sel_0_0(salloc_arb_io_in_2_bits_vc_sel_0_0),
    .io_in_2_bits_tail(salloc_arb_io_in_2_bits_tail),
    .io_in_3_ready(salloc_arb_io_in_3_ready),
    .io_in_3_valid(salloc_arb_io_in_3_valid),
    .io_in_3_bits_vc_sel_0_0(salloc_arb_io_in_3_bits_vc_sel_0_0),
    .io_in_3_bits_tail(salloc_arb_io_in_3_bits_tail),
    .io_out_0_ready(salloc_arb_io_out_0_ready),
    .io_out_0_valid(salloc_arb_io_out_0_valid),
    .io_out_0_bits_vc_sel_0_0(salloc_arb_io_out_0_bits_vc_sel_0_0),
    .io_out_0_bits_tail(salloc_arb_io_out_0_bits_tail),
    .io_chosen_oh_0(salloc_arb_io_chosen_oh_0)
  );
  assign io_router_req_valid = route_arbiter_io_out_valid; // @[InputUnit.scala 189:17]
  assign io_router_req_bits_src_virt_id = route_arbiter_io_out_bits_src_virt_id; // @[InputUnit.scala 189:17]
  assign io_vcalloc_req_valid = vcalloc_vals_1 | vcalloc_vals_2 | vcalloc_vals_3; // @[package.scala 73:59]
  assign io_vcalloc_req_bits_vc_sel_0_0 = vcalloc_sel[1] & states_1_vc_sel_0_0 | vcalloc_sel[2] & states_2_vc_sel_0_0 |
    vcalloc_sel[3] & states_3_vc_sel_0_0; // @[Mux.scala 27:73]
  assign io_salloc_req_0_valid = salloc_arb_io_out_0_valid; // @[InputUnit.scala 302:17 303:19 305:35]
  assign io_salloc_req_0_bits_vc_sel_0_0 = salloc_arb_io_out_0_bits_vc_sel_0_0; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_tail = salloc_arb_io_out_0_bits_tail; // @[InputUnit.scala 302:17]
  assign io_out_0_valid = salloc_outs_0_valid; // @[InputUnit.scala 349:21]
  assign io_out_0_bits_flit_head = salloc_outs_0_flit_head; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_flit_tail = salloc_outs_0_flit_tail; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_flit_payload = salloc_outs_0_flit_payload; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_flit_flow_ingress_node = salloc_outs_0_flit_flow_ingress_node; // @[InputUnit.scala 350:25]
  assign io_debug_va_stall = _io_debug_va_stall_T_7[1:0]; // @[InputUnit.scala 266:21]
  assign io_debug_sa_stall = _io_debug_sa_stall_T_12[1:0]; // @[InputUnit.scala 301:21]
  assign io_in_credit_return = _io_in_credit_return_T ? salloc_arb_io_chosen_oh_0 : 4'h0; // @[InputUnit.scala 322:8]
  assign io_in_vc_free = _io_in_credit_return_T & _io_in_vc_free_T_11 ? salloc_arb_io_chosen_oh_0 : 4'h0; // @[InputUnit.scala 325:8]
  assign input_buffer_clock = clock;
  assign input_buffer_reset = reset;
  assign input_buffer_io_enq_0_valid = io_in_flit_0_valid; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_head = io_in_flit_0_bits_head; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_tail = io_in_flit_0_bits_tail; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_payload = io_in_flit_0_bits_payload; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_virt_channel_id = io_in_flit_0_bits_virt_channel_id; // @[InputUnit.scala 182:28]
  assign input_buffer_io_deq_1_ready = salloc_arb_io_in_1_ready; // @[InputUnit.scala 295:36]
  assign input_buffer_io_deq_2_ready = salloc_arb_io_in_2_ready; // @[InputUnit.scala 295:36]
  assign input_buffer_io_deq_3_ready = salloc_arb_io_in_3_ready; // @[InputUnit.scala 295:36]
  assign route_arbiter_io_in_1_valid = states_1_g == 3'h1; // @[InputUnit.scala 212:22]
  assign route_arbiter_io_in_2_valid = states_2_g == 3'h1; // @[InputUnit.scala 212:22]
  assign route_arbiter_io_in_3_valid = states_3_g == 3'h1; // @[InputUnit.scala 212:22]
  assign salloc_arb_clock = clock;
  assign salloc_arb_reset = reset;
  assign salloc_arb_io_in_0_valid = 1'h0; // @[InputUnit.scala 297:15]
  assign salloc_arb_io_in_1_valid = states_1_g == 3'h3 & credit_available & input_buffer_io_deq_1_valid; // @[InputUnit.scala 288:50]
  assign salloc_arb_io_in_1_bits_vc_sel_0_0 = states_1_vc_sel_0_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_1_bits_tail = input_buffer_io_deq_1_bits_tail; // @[InputUnit.scala 291:19]
  assign salloc_arb_io_in_2_valid = states_2_g == 3'h3 & credit_available_1 & input_buffer_io_deq_2_valid; // @[InputUnit.scala 288:50]
  assign salloc_arb_io_in_2_bits_vc_sel_0_0 = states_2_vc_sel_0_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_tail = input_buffer_io_deq_2_bits_tail; // @[InputUnit.scala 291:19]
  assign salloc_arb_io_in_3_valid = states_3_g == 3'h3 & credit_available_2 & input_buffer_io_deq_3_valid; // @[InputUnit.scala 288:50]
  assign salloc_arb_io_in_3_bits_vc_sel_0_0 = states_3_vc_sel_0_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_tail = input_buffer_io_deq_3_bits_tail; // @[InputUnit.scala 291:19]
  assign salloc_arb_io_out_0_ready = io_salloc_req_0_ready; // @[InputUnit.scala 302:17 303:19 304:39]
  always @(posedge clock) begin
    if (reset) begin // @[InputUnit.scala 377:23]
      states_1_g <= 3'h0; // @[InputUnit.scala 378:24]
    end else if (_T_56 & input_buffer_io_deq_1_bits_tail) begin // @[InputUnit.scala 292:35]
      states_1_g <= 3'h0; // @[InputUnit.scala 293:13]
    end else if (_T_35) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_g <= 3'h3; // @[InputUnit.scala 272:21]
      end else begin
        states_1_g <= _GEN_93;
      end
    end else begin
      states_1_g <= _GEN_93;
    end
    if (_T_35) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_vc_sel_0_0 <= io_vcalloc_resp_vc_sel_0_0; // @[InputUnit.scala 271:26]
      end else begin
        states_1_vc_sel_0_0 <= _GEN_88;
      end
    end else begin
      states_1_vc_sel_0_0 <= _GEN_88;
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h1 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_1_flow_ingress_node <= io_in_flit_0_bits_flow_ingress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (reset) begin // @[InputUnit.scala 377:23]
      states_2_g <= 3'h0; // @[InputUnit.scala 378:24]
    end else if (_T_58 & input_buffer_io_deq_2_bits_tail) begin // @[InputUnit.scala 292:35]
      states_2_g <= 3'h0; // @[InputUnit.scala 293:13]
    end else if (_T_35) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_g <= 3'h3; // @[InputUnit.scala 272:21]
      end else begin
        states_2_g <= _GEN_94;
      end
    end else begin
      states_2_g <= _GEN_94;
    end
    if (_T_35) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_0_0 <= io_vcalloc_resp_vc_sel_0_0; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_0_0 <= _GEN_89;
      end
    end else begin
      states_2_vc_sel_0_0 <= _GEN_89;
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h2 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_2_flow_ingress_node <= io_in_flit_0_bits_flow_ingress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (reset) begin // @[InputUnit.scala 377:23]
      states_3_g <= 3'h0; // @[InputUnit.scala 378:24]
    end else if (_T_60 & input_buffer_io_deq_3_bits_tail) begin // @[InputUnit.scala 292:35]
      states_3_g <= 3'h0; // @[InputUnit.scala 293:13]
    end else if (_T_35) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_g <= 3'h3; // @[InputUnit.scala 272:21]
      end else begin
        states_3_g <= _GEN_95;
      end
    end else begin
      states_3_g <= _GEN_95;
    end
    if (_T_35) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_0_0 <= io_vcalloc_resp_vc_sel_0_0; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_0_0 <= _GEN_90;
      end
    end else begin
      states_3_vc_sel_0_0 <= _GEN_90;
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h3 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_3_flow_ingress_node <= io_in_flit_0_bits_flow_ingress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (reset) begin // @[InputUnit.scala 233:21]
      mask <= 4'h0; // @[InputUnit.scala 233:21]
    end else if (io_router_req_valid) begin // @[InputUnit.scala 239:31]
      mask <= _mask_T_2; // @[InputUnit.scala 240:10]
    end else if (_T_25) begin // @[InputUnit.scala 241:34]
      mask <= _mask_T_17; // @[InputUnit.scala 242:10]
    end
    salloc_outs_0_valid <= salloc_arb_io_out_0_ready & salloc_arb_io_out_0_valid; // @[Decoupled.scala 51:35]
    salloc_outs_0_flit_head <= salloc_arb_io_chosen_oh_0[0] & input_buffer_io_deq_0_bits_head |
      salloc_arb_io_chosen_oh_0[1] & input_buffer_io_deq_1_bits_head | salloc_arb_io_chosen_oh_0[2] &
      input_buffer_io_deq_2_bits_head | salloc_arb_io_chosen_oh_0[3] & input_buffer_io_deq_3_bits_head; // @[Mux.scala 27:73]
    salloc_outs_0_flit_tail <= salloc_arb_io_chosen_oh_0[0] & input_buffer_io_deq_0_bits_tail |
      salloc_arb_io_chosen_oh_0[1] & input_buffer_io_deq_1_bits_tail | salloc_arb_io_chosen_oh_0[2] &
      input_buffer_io_deq_2_bits_tail | salloc_arb_io_chosen_oh_0[3] & input_buffer_io_deq_3_bits_tail; // @[Mux.scala 27:73]
    salloc_outs_0_flit_payload <= _salloc_outs_0_flit_payload_T_9 | _salloc_outs_0_flit_payload_T_7; // @[Mux.scala 27:73]
    salloc_outs_0_flit_flow_ingress_node <= _salloc_outs_0_flit_flow_T_30 | _salloc_outs_0_flit_flow_T_28; // @[Mux.scala 27:73]
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T & _T_3 & ~(_GEN_3 == 3'h0)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:197 assert(states(id).g === g_i)\n"); // @[InputUnit.scala 197:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_router_req_valid & _T_3 & ~(_GEN_74 == 3'h1)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:224 assert(states(id).g === g_r)\n"); // @[InputUnit.scala 224:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_35 & vcalloc_sel[0] & _T_3) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:274 assert(states(i).g === g_v)\n"); // @[InputUnit.scala 274:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_35 & vcalloc_sel[1] & _T_3 & ~vcalloc_vals_1) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:274 assert(states(i).g === g_v)\n"); // @[InputUnit.scala 274:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_35 & vcalloc_sel[2] & _T_3 & ~vcalloc_vals_2) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:274 assert(states(i).g === g_v)\n"); // @[InputUnit.scala 274:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_35 & vcalloc_sel[3] & _T_3 & ~vcalloc_vals_3) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:274 assert(states(i).g === g_v)\n"); // @[InputUnit.scala 274:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  states_1_g = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  states_1_vc_sel_0_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  states_1_flow_ingress_node = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  states_2_g = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  states_2_vc_sel_0_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  states_2_flow_ingress_node = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  states_3_g = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  states_3_vc_sel_0_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  states_3_flow_ingress_node = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  mask = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  salloc_outs_0_valid = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  salloc_outs_0_flit_head = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  salloc_outs_0_flit_tail = _RAND_12[0:0];
  _RAND_13 = {2{`RANDOM}};
  salloc_outs_0_flit_payload = _RAND_13[63:0];
  _RAND_14 = {1{`RANDOM}};
  salloc_outs_0_flit_flow_ingress_node = _RAND_14[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (_T & ~reset) begin
      assert(1'h1); // @[InputUnit.scala 196:13]
    end
    //
    if (_T & _T_3) begin
      assert(_GEN_3 == 3'h0); // @[InputUnit.scala 197:13]
    end
    //
    if (io_router_req_valid & _T_3) begin
      assert(_GEN_74 == 3'h1); // @[InputUnit.scala 224:11]
    end
    //
    if (_T_35 & vcalloc_sel[0] & _T_3) begin
      assert(1'h0); // @[InputUnit.scala 274:17]
    end
    //
    if (_T_35 & vcalloc_sel[1] & _T_3) begin
      assert(vcalloc_vals_1); // @[InputUnit.scala 274:17]
    end
    //
    if (_T_35 & vcalloc_sel[2] & _T_3) begin
      assert(vcalloc_vals_2); // @[InputUnit.scala 274:17]
    end
    //
    if (_T_35 & vcalloc_sel[3] & _T_3) begin
      assert(vcalloc_vals_3); // @[InputUnit.scala 274:17]
    end
  end
endmodule
module Queue_12(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_head,
  input         io_enq_bits_tail,
  input  [63:0] io_enq_bits_payload,
  input         io_enq_bits_ingress_id,
  output        io_deq_valid,
  output        io_deq_bits_head,
  output        io_deq_bits_tail,
  output [63:0] io_deq_bits_payload,
  output        io_deq_bits_ingress_id,
  output [1:0]  io_count
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg  ram_head [0:2]; // @[Decoupled.scala 273:95]
  wire  ram_head_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [1:0] ram_head_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_head_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_head_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_tail [0:2]; // @[Decoupled.scala 273:95]
  wire  ram_tail_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [1:0] ram_tail_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_tail_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_tail_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_en; // @[Decoupled.scala 273:95]
  reg [63:0] ram_payload [0:2]; // @[Decoupled.scala 273:95]
  wire  ram_payload_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [1:0] ram_payload_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [63:0] ram_payload_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [63:0] ram_payload_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_payload_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_payload_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_payload_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_ingress_id [0:2]; // @[Decoupled.scala 273:95]
  wire  ram_ingress_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [1:0] ram_ingress_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_ingress_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_ingress_id_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_ingress_id_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_ingress_id_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_ingress_id_MPORT_en; // @[Decoupled.scala 273:95]
  reg [1:0] enq_ptr_value; // @[Counter.scala 61:40]
  reg [1:0] deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  wrap = enq_ptr_value == 2'h2; // @[Counter.scala 73:24]
  wire [1:0] _value_T_1 = enq_ptr_value + 2'h1; // @[Counter.scala 77:24]
  wire  do_enq = empty ? 1'h0 : _do_enq_T; // @[Decoupled.scala 315:17 280:27]
  wire  wrap_1 = deq_ptr_value == 2'h2; // @[Counter.scala 73:24]
  wire [1:0] _value_T_3 = deq_ptr_value + 2'h1; // @[Counter.scala 77:24]
  wire  do_deq = empty ? 1'h0 : io_deq_valid; // @[Decoupled.scala 315:17 317:14 281:27]
  wire [1:0] ptr_diff = enq_ptr_value - deq_ptr_value; // @[Decoupled.scala 326:32]
  wire [1:0] _io_count_T = maybe_full ? 2'h3 : 2'h0; // @[Decoupled.scala 333:10]
  wire [1:0] _io_count_T_3 = 2'h3 + ptr_diff; // @[Decoupled.scala 334:57]
  wire [1:0] _io_count_T_4 = deq_ptr_value > enq_ptr_value ? _io_count_T_3 : ptr_diff; // @[Decoupled.scala 334:10]
  assign ram_head_io_deq_bits_MPORT_en = 1'h1;
  assign ram_head_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_head_io_deq_bits_MPORT_data = ram_head[ram_head_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  `else
  assign ram_head_io_deq_bits_MPORT_data = ram_head_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_1[0:0] :
    ram_head[ram_head_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_head_MPORT_data = io_enq_bits_head;
  assign ram_head_MPORT_addr = enq_ptr_value;
  assign ram_head_MPORT_mask = 1'h1;
  assign ram_head_MPORT_en = empty ? 1'h0 : _do_enq_T;
  assign ram_tail_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tail_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_tail_io_deq_bits_MPORT_data = ram_tail[ram_tail_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  `else
  assign ram_tail_io_deq_bits_MPORT_data = ram_tail_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_3[0:0] :
    ram_tail[ram_tail_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_tail_MPORT_data = io_enq_bits_tail;
  assign ram_tail_MPORT_addr = enq_ptr_value;
  assign ram_tail_MPORT_mask = 1'h1;
  assign ram_tail_MPORT_en = empty ? 1'h0 : _do_enq_T;
  assign ram_payload_io_deq_bits_MPORT_en = 1'h1;
  assign ram_payload_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_payload_io_deq_bits_MPORT_data = ram_payload[ram_payload_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  `else
  assign ram_payload_io_deq_bits_MPORT_data = ram_payload_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_5[63:0] :
    ram_payload[ram_payload_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_payload_MPORT_data = io_enq_bits_payload;
  assign ram_payload_MPORT_addr = enq_ptr_value;
  assign ram_payload_MPORT_mask = 1'h1;
  assign ram_payload_MPORT_en = empty ? 1'h0 : _do_enq_T;
  assign ram_ingress_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_ingress_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_ingress_id_io_deq_bits_MPORT_data = ram_ingress_id[ram_ingress_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  `else
  assign ram_ingress_id_io_deq_bits_MPORT_data = ram_ingress_id_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_7[0:0] :
    ram_ingress_id[ram_ingress_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_ingress_id_MPORT_data = io_enq_bits_ingress_id;
  assign ram_ingress_id_MPORT_addr = enq_ptr_value;
  assign ram_ingress_id_MPORT_mask = 1'h1;
  assign ram_ingress_id_MPORT_en = empty ? 1'h0 : _do_enq_T;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 302:16 314:{24,39}]
  assign io_deq_bits_head = empty ? io_enq_bits_head : ram_head_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_tail = empty ? io_enq_bits_tail : ram_tail_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_payload = empty ? io_enq_bits_payload : ram_payload_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_ingress_id = empty ? io_enq_bits_ingress_id : ram_ingress_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_count = ptr_match ? _io_count_T : _io_count_T_4; // @[Decoupled.scala 331:20]
  always @(posedge clock) begin
    if (ram_head_MPORT_en & ram_head_MPORT_mask) begin
      ram_head[ram_head_MPORT_addr] <= ram_head_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_tail_MPORT_en & ram_tail_MPORT_mask) begin
      ram_tail[ram_tail_MPORT_addr] <= ram_tail_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_payload_MPORT_en & ram_payload_MPORT_mask) begin
      ram_payload[ram_payload_MPORT_addr] <= ram_payload_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_ingress_id_MPORT_en & ram_ingress_id_MPORT_mask) begin
      ram_ingress_id[ram_ingress_id_MPORT_addr] <= ram_ingress_id_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 2'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      if (wrap) begin // @[Counter.scala 87:20]
        enq_ptr_value <= 2'h0; // @[Counter.scala 87:28]
      end else begin
        enq_ptr_value <= _value_T_1; // @[Counter.scala 77:15]
      end
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 2'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      if (wrap_1) begin // @[Counter.scala 87:20]
        deq_ptr_value <= 2'h0; // @[Counter.scala 87:28]
      end else begin
        deq_ptr_value <= _value_T_3; // @[Counter.scala 77:15]
      end
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      if (empty) begin // @[Decoupled.scala 315:17]
        maybe_full <= 1'h0;
      end else begin
        maybe_full <= _do_enq_T; // @[Decoupled.scala 280:27]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {1{`RANDOM}};
  _RAND_3 = {1{`RANDOM}};
  _RAND_5 = {2{`RANDOM}};
  _RAND_7 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_head[initvar] = _RAND_0[0:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_tail[initvar] = _RAND_2[0:0];
  _RAND_4 = {2{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_payload[initvar] = _RAND_4[63:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram_ingress_id[initvar] = _RAND_6[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  enq_ptr_value = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  deq_ptr_value = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  maybe_full = _RAND_10[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module EgressUnit(
  input         clock,
  input         reset,
  input         io_in_0_valid,
  input         io_in_0_bits_head,
  input         io_in_0_bits_tail,
  input  [63:0] io_in_0_bits_payload,
  input  [1:0]  io_in_0_bits_flow_ingress_node,
  output        io_credit_available_0,
  output        io_channel_status_0_occupied,
  input         io_allocs_0_alloc,
  input         io_credit_alloc_0_alloc,
  input         io_credit_alloc_0_tail,
  output        io_out_valid,
  output        io_out_bits_head,
  output        io_out_bits_tail,
  output [63:0] io_out_bits_payload,
  output        io_out_bits_ingress_id
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  q_clock; // @[EgressUnit.scala 22:17]
  wire  q_reset; // @[EgressUnit.scala 22:17]
  wire  q_io_enq_ready; // @[EgressUnit.scala 22:17]
  wire  q_io_enq_valid; // @[EgressUnit.scala 22:17]
  wire  q_io_enq_bits_head; // @[EgressUnit.scala 22:17]
  wire  q_io_enq_bits_tail; // @[EgressUnit.scala 22:17]
  wire [63:0] q_io_enq_bits_payload; // @[EgressUnit.scala 22:17]
  wire  q_io_enq_bits_ingress_id; // @[EgressUnit.scala 22:17]
  wire  q_io_deq_valid; // @[EgressUnit.scala 22:17]
  wire  q_io_deq_bits_head; // @[EgressUnit.scala 22:17]
  wire  q_io_deq_bits_tail; // @[EgressUnit.scala 22:17]
  wire [63:0] q_io_deq_bits_payload; // @[EgressUnit.scala 22:17]
  wire  q_io_deq_bits_ingress_id; // @[EgressUnit.scala 22:17]
  wire [1:0] q_io_count; // @[EgressUnit.scala 22:17]
  reg  channel_empty; // @[EgressUnit.scala 20:30]
  wire  _GEN_0 = io_credit_alloc_0_alloc & io_credit_alloc_0_tail | channel_empty; // @[EgressUnit.scala 44:62 45:19 20:30]
  wire  _GEN_1 = io_allocs_0_alloc ? 1'h0 : _GEN_0; // @[EgressUnit.scala 49:29 50:19]
  Queue_12 q ( // @[EgressUnit.scala 22:17]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_head(q_io_enq_bits_head),
    .io_enq_bits_tail(q_io_enq_bits_tail),
    .io_enq_bits_payload(q_io_enq_bits_payload),
    .io_enq_bits_ingress_id(q_io_enq_bits_ingress_id),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_head(q_io_deq_bits_head),
    .io_deq_bits_tail(q_io_deq_bits_tail),
    .io_deq_bits_payload(q_io_deq_bits_payload),
    .io_deq_bits_ingress_id(q_io_deq_bits_ingress_id),
    .io_count(q_io_count)
  );
  assign io_credit_available_0 = q_io_count == 2'h0; // @[EgressUnit.scala 40:40]
  assign io_channel_status_0_occupied = ~channel_empty; // @[EgressUnit.scala 41:36]
  assign io_out_valid = q_io_deq_valid; // @[EgressUnit.scala 37:10]
  assign io_out_bits_head = q_io_deq_bits_head; // @[EgressUnit.scala 37:10]
  assign io_out_bits_tail = q_io_deq_bits_tail; // @[EgressUnit.scala 37:10]
  assign io_out_bits_payload = q_io_deq_bits_payload; // @[EgressUnit.scala 37:10]
  assign io_out_bits_ingress_id = q_io_deq_bits_ingress_id; // @[EgressUnit.scala 37:10]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_in_0_valid; // @[EgressUnit.scala 23:18]
  assign q_io_enq_bits_head = io_in_0_bits_head; // @[EgressUnit.scala 24:22]
  assign q_io_enq_bits_tail = io_in_0_bits_tail; // @[EgressUnit.scala 25:22]
  assign q_io_enq_bits_payload = io_in_0_bits_payload; // @[EgressUnit.scala 36:25]
  assign q_io_enq_bits_ingress_id = 2'h2 == io_in_0_bits_flow_ingress_node; // @[EgressUnit.scala 31:39]
  always @(posedge clock) begin
    channel_empty <= reset | _GEN_1; // @[EgressUnit.scala 20:{30,30}]
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~(q_io_enq_valid & ~q_io_enq_ready))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at EgressUnit.scala:38 assert(!(q.io.enq.valid && !q.io.enq.ready))\n"); // @[EgressUnit.scala 38:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  channel_empty = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(~(q_io_enq_valid & ~q_io_enq_ready)); // @[EgressUnit.scala 38:9]
    end
  end
endmodule
module Switch_1(
  input         clock,
  input         reset,
  input         io_in_1_0_valid,
  input         io_in_1_0_bits_flit_head,
  input         io_in_1_0_bits_flit_tail,
  input  [63:0] io_in_1_0_bits_flit_payload,
  input  [1:0]  io_in_1_0_bits_flit_flow_ingress_node,
  input         io_in_0_0_valid,
  input         io_in_0_0_bits_flit_head,
  input         io_in_0_0_bits_flit_tail,
  input  [63:0] io_in_0_0_bits_flit_payload,
  input  [1:0]  io_in_0_0_bits_flit_flow_ingress_node,
  output        io_out_0_0_valid,
  output        io_out_0_0_bits_head,
  output        io_out_0_0_bits_tail,
  output [63:0] io_out_0_0_bits_payload,
  output [1:0]  io_out_0_0_bits_flow_ingress_node,
  input         io_sel_0_0_1_0,
  input         io_sel_0_0_0_0
);
  wire [1:0] sel_flat = {io_sel_0_0_1_0,io_sel_0_0_0_0}; // @[Switch.scala 46:35]
  wire [1:0] _T_2 = sel_flat[0] + sel_flat[1]; // @[Bitwise.scala 51:90]
  wire  _io_out_0_0_valid_T_4 = sel_flat[0] & io_in_0_0_valid | sel_flat[1] & io_in_1_0_valid; // @[Mux.scala 27:73]
  wire [1:0] _io_out_0_0_bits_T_14 = sel_flat[0] ? io_in_0_0_bits_flit_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_0_0_bits_T_15 = sel_flat[1] ? io_in_1_0_bits_flit_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_out_0_0_bits_T_20 = sel_flat[0] ? io_in_0_0_bits_flit_payload : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_out_0_0_bits_T_21 = sel_flat[1] ? io_in_1_0_bits_flit_payload : 64'h0; // @[Mux.scala 27:73]
  assign io_out_0_0_valid = _io_out_0_0_valid_T_4 & sel_flat != 2'h0; // @[Switch.scala 48:67]
  assign io_out_0_0_bits_head = sel_flat[0] & io_in_0_0_bits_flit_head | sel_flat[1] & io_in_1_0_bits_flit_head; // @[Mux.scala 27:73]
  assign io_out_0_0_bits_tail = sel_flat[0] & io_in_0_0_bits_flit_tail | sel_flat[1] & io_in_1_0_bits_flit_tail; // @[Mux.scala 27:73]
  assign io_out_0_0_bits_payload = _io_out_0_0_bits_T_20 | _io_out_0_0_bits_T_21; // @[Mux.scala 27:73]
  assign io_out_0_0_bits_flow_ingress_node = _io_out_0_0_bits_T_14 | _io_out_0_0_bits_T_15; // @[Mux.scala 27:73]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(_T_2 <= 2'h1)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Switch.scala:47 assert(PopCount(sel_flat) <= 1.U)\n"); // @[Switch.scala 47:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(_T_2 <= 2'h1); // @[Switch.scala 47:13]
    end
  end
endmodule
module SwitchArbiter_4(
  input        clock,
  input        reset,
  output       io_in_0_ready,
  input        io_in_0_valid,
  input        io_in_0_bits_vc_sel_0_0,
  input        io_in_0_bits_tail,
  output       io_in_1_ready,
  input        io_in_1_valid,
  input        io_in_1_bits_vc_sel_0_0,
  input        io_in_1_bits_tail,
  output       io_out_0_valid,
  output       io_out_0_bits_vc_sel_0_0,
  output       io_out_0_bits_tail,
  output [1:0] io_chosen_oh_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] lock_0; // @[SwitchAllocator.scala 24:38]
  wire [1:0] _unassigned_T = {io_in_1_valid,io_in_0_valid}; // @[Cat.scala 33:92]
  wire [1:0] _unassigned_T_1 = ~lock_0; // @[SwitchAllocator.scala 25:54]
  wire [1:0] unassigned = _unassigned_T & _unassigned_T_1; // @[SwitchAllocator.scala 25:52]
  reg [1:0] mask; // @[SwitchAllocator.scala 27:21]
  wire [1:0] _GEN_4 = {{1'd0}, mask == 2'h0}; // @[SwitchAllocator.scala 30:58]
  wire [1:0] _sel_T_1 = unassigned & _GEN_4; // @[SwitchAllocator.scala 30:58]
  wire [3:0] _sel_T_2 = {unassigned,_sel_T_1}; // @[Cat.scala 33:92]
  wire [3:0] _sel_T_7 = _sel_T_2[3] ? 4'h8 : 4'h0; // @[Mux.scala 47:70]
  wire [3:0] _sel_T_8 = _sel_T_2[2] ? 4'h4 : _sel_T_7; // @[Mux.scala 47:70]
  wire [3:0] _sel_T_9 = _sel_T_2[1] ? 4'h2 : _sel_T_8; // @[Mux.scala 47:70]
  wire [3:0] sel = _sel_T_2[0] ? 4'h1 : _sel_T_9; // @[Mux.scala 47:70]
  wire [3:0] _GEN_5 = {{2'd0}, sel[3:2]}; // @[SwitchAllocator.scala 32:23]
  wire [3:0] _choices_0_T_1 = sel | _GEN_5; // @[SwitchAllocator.scala 32:23]
  wire [1:0] choices_0 = _choices_0_T_1[1:0]; // @[SwitchAllocator.scala 28:21 32:16]
  wire [1:0] in_tails = {io_in_1_bits_tail,io_in_0_bits_tail}; // @[Cat.scala 33:92]
  wire [1:0] _chosen_T = _unassigned_T & lock_0; // @[SwitchAllocator.scala 42:33]
  wire [1:0] chosen = |_chosen_T ? lock_0 : choices_0; // @[SwitchAllocator.scala 42:21]
  wire [1:0] _io_out_0_valid_T = _unassigned_T & chosen; // @[SwitchAllocator.scala 44:35]
  wire [1:0] _lock_0_T = ~in_tails; // @[SwitchAllocator.scala 53:27]
  wire [1:0] _lock_0_T_1 = chosen & _lock_0_T; // @[SwitchAllocator.scala 53:25]
  wire [1:0] _GEN_6 = {{1'd0}, io_chosen_oh_0[1]}; // @[SwitchAllocator.scala 58:71]
  wire [1:0] _mask_T_2 = io_chosen_oh_0 | _GEN_6; // @[SwitchAllocator.scala 58:71]
  wire [1:0] _mask_T_3 = ~mask; // @[SwitchAllocator.scala 60:17]
  wire [2:0] _mask_T_5 = {mask, 1'h0}; // @[SwitchAllocator.scala 60:43]
  wire [2:0] _mask_T_6 = _mask_T_5 | 3'h1; // @[SwitchAllocator.scala 60:49]
  wire [2:0] _mask_T_7 = _mask_T_3 == 2'h0 ? 3'h0 : _mask_T_6; // @[SwitchAllocator.scala 60:16]
  wire [2:0] _GEN_3 = io_out_0_valid ? {{1'd0}, _mask_T_2} : _mask_T_7; // @[SwitchAllocator.scala 57:27 58:10 60:10]
  wire [2:0] _GEN_7 = reset ? 3'h0 : _GEN_3; // @[SwitchAllocator.scala 27:{21,21}]
  assign io_in_0_ready = chosen[0]; // @[SwitchAllocator.scala 47:19]
  assign io_in_1_ready = chosen[1]; // @[SwitchAllocator.scala 47:19]
  assign io_out_0_valid = |_io_out_0_valid_T; // @[SwitchAllocator.scala 44:45]
  assign io_out_0_bits_vc_sel_0_0 = chosen[0] & io_in_0_bits_vc_sel_0_0 | chosen[1] & io_in_1_bits_vc_sel_0_0; // @[Mux.scala 27:73]
  assign io_out_0_bits_tail = chosen[0] & io_in_0_bits_tail | chosen[1] & io_in_1_bits_tail; // @[Mux.scala 27:73]
  assign io_chosen_oh_0 = |_chosen_T ? lock_0 : choices_0; // @[SwitchAllocator.scala 42:21]
  always @(posedge clock) begin
    if (reset) begin // @[SwitchAllocator.scala 24:38]
      lock_0 <= 2'h0; // @[SwitchAllocator.scala 24:38]
    end else if (io_out_0_valid) begin // @[SwitchAllocator.scala 52:29]
      lock_0 <= _lock_0_T_1; // @[SwitchAllocator.scala 53:15]
    end
    mask <= _GEN_7[1:0]; // @[SwitchAllocator.scala 27:{21,21}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lock_0 = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  mask = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SwitchAllocator_1(
  input   clock,
  input   reset,
  output  io_req_1_0_ready,
  input   io_req_1_0_valid,
  input   io_req_1_0_bits_vc_sel_0_0,
  input   io_req_1_0_bits_tail,
  output  io_req_0_0_ready,
  input   io_req_0_0_valid,
  input   io_req_0_0_bits_vc_sel_0_0,
  input   io_req_0_0_bits_tail,
  output  io_credit_alloc_0_0_alloc,
  output  io_credit_alloc_0_0_tail,
  output  io_switch_sel_0_0_1_0,
  output  io_switch_sel_0_0_0_0
);
  wire  arbs_0_clock; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_reset; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_0_ready; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_0_valid; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_0_bits_vc_sel_0_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_0_bits_tail; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_1_ready; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_1_valid; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_1_bits_vc_sel_0_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_in_1_bits_tail; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_out_0_valid; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_out_0_bits_vc_sel_0_0; // @[SwitchAllocator.scala 83:45]
  wire  arbs_0_io_out_0_bits_tail; // @[SwitchAllocator.scala 83:45]
  wire [1:0] arbs_0_io_chosen_oh_0; // @[SwitchAllocator.scala 83:45]
  SwitchArbiter_4 arbs_0 ( // @[SwitchAllocator.scala 83:45]
    .clock(arbs_0_clock),
    .reset(arbs_0_reset),
    .io_in_0_ready(arbs_0_io_in_0_ready),
    .io_in_0_valid(arbs_0_io_in_0_valid),
    .io_in_0_bits_vc_sel_0_0(arbs_0_io_in_0_bits_vc_sel_0_0),
    .io_in_0_bits_tail(arbs_0_io_in_0_bits_tail),
    .io_in_1_ready(arbs_0_io_in_1_ready),
    .io_in_1_valid(arbs_0_io_in_1_valid),
    .io_in_1_bits_vc_sel_0_0(arbs_0_io_in_1_bits_vc_sel_0_0),
    .io_in_1_bits_tail(arbs_0_io_in_1_bits_tail),
    .io_out_0_valid(arbs_0_io_out_0_valid),
    .io_out_0_bits_vc_sel_0_0(arbs_0_io_out_0_bits_vc_sel_0_0),
    .io_out_0_bits_tail(arbs_0_io_out_0_bits_tail),
    .io_chosen_oh_0(arbs_0_io_chosen_oh_0)
  );
  assign io_req_1_0_ready = arbs_0_io_in_1_ready & arbs_0_io_in_1_valid; // @[Decoupled.scala 51:35]
  assign io_req_0_0_ready = arbs_0_io_in_0_ready & arbs_0_io_in_0_valid; // @[Decoupled.scala 51:35]
  assign io_credit_alloc_0_0_alloc = arbs_0_io_out_0_valid & arbs_0_io_out_0_bits_vc_sel_0_0; // @[SwitchAllocator.scala 120:33]
  assign io_credit_alloc_0_0_tail = arbs_0_io_out_0_valid & arbs_0_io_out_0_bits_vc_sel_0_0 & arbs_0_io_out_0_bits_tail; // @[SwitchAllocator.scala 120:67 122:21 116:44]
  assign io_switch_sel_0_0_1_0 = arbs_0_io_in_1_valid & arbs_0_io_chosen_oh_0[1] & arbs_0_io_out_0_valid; // @[SwitchAllocator.scala 108:97]
  assign io_switch_sel_0_0_0_0 = arbs_0_io_in_0_valid & arbs_0_io_chosen_oh_0[0] & arbs_0_io_out_0_valid; // @[SwitchAllocator.scala 108:97]
  assign arbs_0_clock = clock;
  assign arbs_0_reset = reset;
  assign arbs_0_io_in_0_valid = io_req_0_0_valid & io_req_0_0_bits_vc_sel_0_0; // @[SwitchAllocator.scala 95:37]
  assign arbs_0_io_in_0_bits_vc_sel_0_0 = io_req_0_0_bits_vc_sel_0_0; // @[SwitchAllocator.scala 96:25]
  assign arbs_0_io_in_0_bits_tail = io_req_0_0_bits_tail; // @[SwitchAllocator.scala 96:25]
  assign arbs_0_io_in_1_valid = io_req_1_0_valid & io_req_1_0_bits_vc_sel_0_0; // @[SwitchAllocator.scala 95:37]
  assign arbs_0_io_in_1_bits_vc_sel_0_0 = io_req_1_0_bits_vc_sel_0_0; // @[SwitchAllocator.scala 96:25]
  assign arbs_0_io_in_1_bits_tail = io_req_1_0_bits_tail; // @[SwitchAllocator.scala 96:25]
endmodule
module RotatingSingleVCAllocator_1(
  input   clock,
  input   reset,
  output  io_req_1_ready,
  input   io_req_1_valid,
  input   io_req_1_bits_vc_sel_0_0,
  output  io_req_0_ready,
  input   io_req_0_valid,
  input   io_req_0_bits_vc_sel_0_0,
  output  io_resp_1_vc_sel_0_0,
  output  io_resp_0_vc_sel_0_0,
  input   io_channel_status_0_0_occupied,
  output  io_out_allocs_0_0_alloc
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] mask; // @[SingleVCAllocator.scala 16:21]
  wire  in_arb_reqs_1_0_0 = io_req_1_bits_vc_sel_0_0 & ~io_channel_status_0_0_occupied; // @[SingleVCAllocator.scala 28:61]
  wire  in_arb_vals_1 = io_req_1_valid & in_arb_reqs_1_0_0; // @[SingleVCAllocator.scala 32:39]
  wire  in_arb_reqs_0_0_0 = io_req_0_bits_vc_sel_0_0 & ~io_channel_status_0_0_occupied; // @[SingleVCAllocator.scala 28:61]
  wire  in_arb_vals_0 = io_req_0_valid & in_arb_reqs_0_0_0; // @[SingleVCAllocator.scala 32:39]
  wire [1:0] _in_arb_filter_T = {in_arb_vals_1,in_arb_vals_0}; // @[SingleVCAllocator.scala 19:57]
  wire [1:0] _in_arb_filter_T_2 = ~mask; // @[SingleVCAllocator.scala 19:86]
  wire [1:0] _in_arb_filter_T_3 = _in_arb_filter_T & _in_arb_filter_T_2; // @[SingleVCAllocator.scala 19:84]
  wire [3:0] _in_arb_filter_T_4 = {in_arb_vals_1,in_arb_vals_0,_in_arb_filter_T_3}; // @[Cat.scala 33:92]
  wire [3:0] _in_arb_filter_T_9 = _in_arb_filter_T_4[3] ? 4'h8 : 4'h0; // @[Mux.scala 47:70]
  wire [3:0] _in_arb_filter_T_10 = _in_arb_filter_T_4[2] ? 4'h4 : _in_arb_filter_T_9; // @[Mux.scala 47:70]
  wire [3:0] _in_arb_filter_T_11 = _in_arb_filter_T_4[1] ? 4'h2 : _in_arb_filter_T_10; // @[Mux.scala 47:70]
  wire [3:0] in_arb_filter = _in_arb_filter_T_4[0] ? 4'h1 : _in_arb_filter_T_11; // @[Mux.scala 47:70]
  wire [1:0] in_arb_sel = in_arb_filter[1:0] | in_arb_filter[3:2]; // @[SingleVCAllocator.scala 20:57]
  wire  _T = in_arb_vals_0 | in_arb_vals_1; // @[package.scala 73:59]
  wire [1:0] _mask_T_5 = in_arb_sel[1] ? 2'h3 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _GEN_1 = {{1'd0}, in_arb_sel[0]}; // @[Mux.scala 27:73]
  wire [1:0] _mask_T_6 = _GEN_1 | _mask_T_5; // @[Mux.scala 27:73]
  wire  in_vc_sel_0_0 = in_arb_sel[0] & in_arb_reqs_0_0_0 | in_arb_sel[1] & in_arb_reqs_1_0_0; // @[Mux.scala 27:73]
  assign io_req_1_ready = in_arb_sel[1]; // @[SingleVCAllocator.scala 47:34]
  assign io_req_0_ready = in_arb_sel[0]; // @[SingleVCAllocator.scala 47:34]
  assign io_resp_1_vc_sel_0_0 = _T & in_vc_sel_0_0; // @[SingleVCAllocator.scala 41:18]
  assign io_resp_0_vc_sel_0_0 = _T & in_vc_sel_0_0; // @[SingleVCAllocator.scala 41:18]
  assign io_out_allocs_0_0_alloc = _T & in_vc_sel_0_0; // @[SingleVCAllocator.scala 41:18]
  always @(posedge clock) begin
    if (reset) begin // @[SingleVCAllocator.scala 16:21]
      mask <= 2'h0; // @[SingleVCAllocator.scala 16:21]
    end else if (_T) begin // @[SingleVCAllocator.scala 21:26]
      mask <= _mask_T_6; // @[SingleVCAllocator.scala 22:10]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mask = _RAND_0[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(1'h1); // @[SingleVCAllocator.scala 53:11]
    end
    //
    if (~reset) begin
      assert(1'h1); // @[SingleVCAllocator.scala 53:11]
    end
  end
endmodule
module RouteComputer_1(
  input   clock,
  input   reset,
  input   io_req_1_valid,
  input   io_req_0_valid
);
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~io_req_0_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RouteComputer.scala:48 assert(!req.valid)\n"); // @[RouteComputer.scala 48:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~io_req_1_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RouteComputer.scala:48 assert(!req.valid)\n"); // @[RouteComputer.scala 48:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(~io_req_0_valid); // @[RouteComputer.scala 48:13]
    end
    //
    if (~reset) begin
      assert(~io_req_1_valid); // @[RouteComputer.scala 48:13]
    end
  end
endmodule
module Router_1(
  input         clock,
  input         reset,
  output [1:0]  auto_debug_out_va_stall_0,
  output [1:0]  auto_debug_out_va_stall_1,
  output [1:0]  auto_debug_out_sa_stall_0,
  output [1:0]  auto_debug_out_sa_stall_1,
  output        auto_egress_nodes_out_flit_valid,
  output        auto_egress_nodes_out_flit_bits_head,
  output        auto_egress_nodes_out_flit_bits_tail,
  output [63:0] auto_egress_nodes_out_flit_bits_payload,
  output        auto_egress_nodes_out_flit_bits_ingress_id,
  input         auto_dest_nodes_in_1_flit_0_valid,
  input         auto_dest_nodes_in_1_flit_0_bits_head,
  input         auto_dest_nodes_in_1_flit_0_bits_tail,
  input  [63:0] auto_dest_nodes_in_1_flit_0_bits_payload,
  input  [1:0]  auto_dest_nodes_in_1_flit_0_bits_flow_ingress_node,
  input  [1:0]  auto_dest_nodes_in_1_flit_0_bits_flow_egress_node,
  input  [1:0]  auto_dest_nodes_in_1_flit_0_bits_virt_channel_id,
  output [3:0]  auto_dest_nodes_in_1_credit_return,
  output [3:0]  auto_dest_nodes_in_1_vc_free,
  input         auto_dest_nodes_in_0_flit_0_valid,
  input         auto_dest_nodes_in_0_flit_0_bits_head,
  input         auto_dest_nodes_in_0_flit_0_bits_tail,
  input  [63:0] auto_dest_nodes_in_0_flit_0_bits_payload,
  input  [1:0]  auto_dest_nodes_in_0_flit_0_bits_flow_ingress_node,
  input  [1:0]  auto_dest_nodes_in_0_flit_0_bits_flow_egress_node,
  input  [1:0]  auto_dest_nodes_in_0_flit_0_bits_virt_channel_id,
  output [3:0]  auto_dest_nodes_in_0_credit_return,
  output [3:0]  auto_dest_nodes_in_0_vc_free
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  monitor_clock; // @[Nodes.scala 24:25]
  wire  monitor_reset; // @[Nodes.scala 24:25]
  wire  monitor_io_in_flit_0_valid; // @[Nodes.scala 24:25]
  wire  monitor_io_in_flit_0_bits_head; // @[Nodes.scala 24:25]
  wire  monitor_io_in_flit_0_bits_tail; // @[Nodes.scala 24:25]
  wire [1:0] monitor_io_in_flit_0_bits_flow_ingress_node; // @[Nodes.scala 24:25]
  wire [1:0] monitor_io_in_flit_0_bits_flow_egress_node; // @[Nodes.scala 24:25]
  wire [1:0] monitor_io_in_flit_0_bits_virt_channel_id; // @[Nodes.scala 24:25]
  wire  monitor_1_clock; // @[Nodes.scala 24:25]
  wire  monitor_1_reset; // @[Nodes.scala 24:25]
  wire  monitor_1_io_in_flit_0_valid; // @[Nodes.scala 24:25]
  wire  monitor_1_io_in_flit_0_bits_head; // @[Nodes.scala 24:25]
  wire  monitor_1_io_in_flit_0_bits_tail; // @[Nodes.scala 24:25]
  wire [1:0] monitor_1_io_in_flit_0_bits_flow_ingress_node; // @[Nodes.scala 24:25]
  wire [1:0] monitor_1_io_in_flit_0_bits_flow_egress_node; // @[Nodes.scala 24:25]
  wire [1:0] monitor_1_io_in_flit_0_bits_virt_channel_id; // @[Nodes.scala 24:25]
  wire  input_unit_0_from_0_clock; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_reset; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_router_req_valid; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_0_io_router_req_bits_src_virt_id; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_req_ready; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_req_valid; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_resp_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_out_credit_available_0_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_salloc_req_0_ready; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_salloc_req_0_valid; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_salloc_req_0_bits_tail; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_out_0_valid; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_out_0_bits_flit_head; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_out_0_bits_flit_tail; // @[Router.scala 112:13]
  wire [63:0] input_unit_0_from_0_io_out_0_bits_flit_payload; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_0_io_out_0_bits_flit_flow_ingress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_0_io_debug_va_stall; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_0_io_debug_sa_stall; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_in_flit_0_valid; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_in_flit_0_bits_head; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_in_flit_0_bits_tail; // @[Router.scala 112:13]
  wire [63:0] input_unit_0_from_0_io_in_flit_0_bits_payload; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_0_io_in_flit_0_bits_flow_ingress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_0_io_in_flit_0_bits_flow_egress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_0_io_in_flit_0_bits_virt_channel_id; // @[Router.scala 112:13]
  wire [3:0] input_unit_0_from_0_io_in_credit_return; // @[Router.scala 112:13]
  wire [3:0] input_unit_0_from_0_io_in_vc_free; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_clock; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_reset; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_router_req_valid; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_2_io_router_req_bits_src_virt_id; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_req_ready; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_req_valid; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_resp_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_out_credit_available_0_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_salloc_req_0_ready; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_salloc_req_0_valid; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_salloc_req_0_bits_tail; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_out_0_valid; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_out_0_bits_flit_head; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_out_0_bits_flit_tail; // @[Router.scala 112:13]
  wire [63:0] input_unit_1_from_2_io_out_0_bits_flit_payload; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_2_io_out_0_bits_flit_flow_ingress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_2_io_debug_va_stall; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_2_io_debug_sa_stall; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_in_flit_0_valid; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_in_flit_0_bits_head; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_in_flit_0_bits_tail; // @[Router.scala 112:13]
  wire [63:0] input_unit_1_from_2_io_in_flit_0_bits_payload; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_2_io_in_flit_0_bits_flow_ingress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_2_io_in_flit_0_bits_flow_egress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_2_io_in_flit_0_bits_virt_channel_id; // @[Router.scala 112:13]
  wire [3:0] input_unit_1_from_2_io_in_credit_return; // @[Router.scala 112:13]
  wire [3:0] input_unit_1_from_2_io_in_vc_free; // @[Router.scala 112:13]
  wire  egress_unit_0_to_0_clock; // @[Router.scala 125:13]
  wire  egress_unit_0_to_0_reset; // @[Router.scala 125:13]
  wire  egress_unit_0_to_0_io_in_0_valid; // @[Router.scala 125:13]
  wire  egress_unit_0_to_0_io_in_0_bits_head; // @[Router.scala 125:13]
  wire  egress_unit_0_to_0_io_in_0_bits_tail; // @[Router.scala 125:13]
  wire [63:0] egress_unit_0_to_0_io_in_0_bits_payload; // @[Router.scala 125:13]
  wire [1:0] egress_unit_0_to_0_io_in_0_bits_flow_ingress_node; // @[Router.scala 125:13]
  wire  egress_unit_0_to_0_io_credit_available_0; // @[Router.scala 125:13]
  wire  egress_unit_0_to_0_io_channel_status_0_occupied; // @[Router.scala 125:13]
  wire  egress_unit_0_to_0_io_allocs_0_alloc; // @[Router.scala 125:13]
  wire  egress_unit_0_to_0_io_credit_alloc_0_alloc; // @[Router.scala 125:13]
  wire  egress_unit_0_to_0_io_credit_alloc_0_tail; // @[Router.scala 125:13]
  wire  egress_unit_0_to_0_io_out_valid; // @[Router.scala 125:13]
  wire  egress_unit_0_to_0_io_out_bits_head; // @[Router.scala 125:13]
  wire  egress_unit_0_to_0_io_out_bits_tail; // @[Router.scala 125:13]
  wire [63:0] egress_unit_0_to_0_io_out_bits_payload; // @[Router.scala 125:13]
  wire  egress_unit_0_to_0_io_out_bits_ingress_id; // @[Router.scala 125:13]
  wire  switch_clock; // @[Router.scala 129:24]
  wire  switch_reset; // @[Router.scala 129:24]
  wire  switch_io_in_1_0_valid; // @[Router.scala 129:24]
  wire  switch_io_in_1_0_bits_flit_head; // @[Router.scala 129:24]
  wire  switch_io_in_1_0_bits_flit_tail; // @[Router.scala 129:24]
  wire [63:0] switch_io_in_1_0_bits_flit_payload; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_1_0_bits_flit_flow_ingress_node; // @[Router.scala 129:24]
  wire  switch_io_in_0_0_valid; // @[Router.scala 129:24]
  wire  switch_io_in_0_0_bits_flit_head; // @[Router.scala 129:24]
  wire  switch_io_in_0_0_bits_flit_tail; // @[Router.scala 129:24]
  wire [63:0] switch_io_in_0_0_bits_flit_payload; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_0_0_bits_flit_flow_ingress_node; // @[Router.scala 129:24]
  wire  switch_io_out_0_0_valid; // @[Router.scala 129:24]
  wire  switch_io_out_0_0_bits_head; // @[Router.scala 129:24]
  wire  switch_io_out_0_0_bits_tail; // @[Router.scala 129:24]
  wire [63:0] switch_io_out_0_0_bits_payload; // @[Router.scala 129:24]
  wire [1:0] switch_io_out_0_0_bits_flow_ingress_node; // @[Router.scala 129:24]
  wire  switch_io_sel_0_0_1_0; // @[Router.scala 129:24]
  wire  switch_io_sel_0_0_0_0; // @[Router.scala 129:24]
  wire  switch_allocator_clock; // @[Router.scala 130:34]
  wire  switch_allocator_reset; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_ready; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_valid; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_vc_sel_0_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_tail; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_ready; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_valid; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_0_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_tail; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_0_0_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_0_0_tail; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_0_0_1_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_0_0_0_0; // @[Router.scala 130:34]
  wire  vc_allocator_clock; // @[Router.scala 131:30]
  wire  vc_allocator_reset; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_ready; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_valid; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_bits_vc_sel_0_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_ready; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_valid; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_0_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_1_vc_sel_0_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_0_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_0_0_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_0_0_alloc; // @[Router.scala 131:30]
  wire  route_computer_clock; // @[Router.scala 134:32]
  wire  route_computer_reset; // @[Router.scala 134:32]
  wire  route_computer_io_req_1_valid; // @[Router.scala 134:32]
  wire  route_computer_io_req_0_valid; // @[Router.scala 134:32]
  wire [19:0] plusarg_reader_out; // @[PlusArg.scala 80:11]
  wire  _fires_count_T = vc_allocator_io_req_0_ready & vc_allocator_io_req_0_valid; // @[Decoupled.scala 51:35]
  wire  _fires_count_T_1 = vc_allocator_io_req_1_ready & vc_allocator_io_req_1_valid; // @[Decoupled.scala 51:35]
  reg  switch_io_sel_REG_0_0_1_0; // @[Router.scala 176:14]
  reg  switch_io_sel_REG_0_0_0_0; // @[Router.scala 176:14]
  reg [63:0] debug_tsc; // @[Router.scala 193:28]
  wire [63:0] _debug_tsc_T_1 = debug_tsc + 64'h1; // @[Router.scala 194:28]
  reg [63:0] debug_sample; // @[Router.scala 195:31]
  wire [63:0] _debug_sample_T_1 = debug_sample + 64'h1; // @[Router.scala 196:34]
  wire [19:0] _T_1 = plusarg_reader_out - 20'h1; // @[Router.scala 198:40]
  wire [63:0] _GEN_4 = {{44'd0}, _T_1}; // @[Router.scala 198:24]
  wire  _T_2 = debug_sample == _GEN_4; // @[Router.scala 198:24]
  reg [63:0] util_ctr; // @[Router.scala 201:29]
  reg  fired; // @[Router.scala 202:26]
  wire [63:0] _GEN_5 = {{63'd0}, auto_dest_nodes_in_0_flit_0_valid}; // @[Router.scala 203:28]
  wire [63:0] _util_ctr_T_1 = util_ctr + _GEN_5; // @[Router.scala 203:28]
  wire  _T_8 = plusarg_reader_out != 20'h0 & _T_2 & fired; // @[Router.scala 205:71]
  reg [63:0] util_ctr_1; // @[Router.scala 201:29]
  reg  fired_1; // @[Router.scala 202:26]
  wire [63:0] _GEN_7 = {{63'd0}, auto_dest_nodes_in_1_flit_0_valid}; // @[Router.scala 203:28]
  wire [63:0] _util_ctr_T_3 = util_ctr_1 + _GEN_7; // @[Router.scala 203:28]
  wire  _T_16 = plusarg_reader_out != 20'h0 & _T_2 & fired_1; // @[Router.scala 205:71]
  wire  x1_flit_valid = egress_unit_0_to_0_io_out_valid; // @[Nodes.scala 1212:84 Router.scala 144:65]
  reg [63:0] util_ctr_2; // @[Router.scala 201:29]
  reg  fired_2; // @[Router.scala 202:26]
  wire [63:0] _GEN_9 = {{63'd0}, x1_flit_valid}; // @[Router.scala 203:28]
  wire [63:0] _util_ctr_T_5 = util_ctr_2 + _GEN_9; // @[Router.scala 203:28]
  wire  _T_25 = plusarg_reader_out != 20'h0 & _T_2 & fired_2; // @[Router.scala 205:71]
  wire [1:0] fires_count = _fires_count_T + _fires_count_T_1; // @[Bitwise.scala 51:90]
  NoCMonitor monitor ( // @[Nodes.scala 24:25]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_flit_0_valid(monitor_io_in_flit_0_valid),
    .io_in_flit_0_bits_head(monitor_io_in_flit_0_bits_head),
    .io_in_flit_0_bits_tail(monitor_io_in_flit_0_bits_tail),
    .io_in_flit_0_bits_flow_ingress_node(monitor_io_in_flit_0_bits_flow_ingress_node),
    .io_in_flit_0_bits_flow_egress_node(monitor_io_in_flit_0_bits_flow_egress_node),
    .io_in_flit_0_bits_virt_channel_id(monitor_io_in_flit_0_bits_virt_channel_id)
  );
  NoCMonitor_1 monitor_1 ( // @[Nodes.scala 24:25]
    .clock(monitor_1_clock),
    .reset(monitor_1_reset),
    .io_in_flit_0_valid(monitor_1_io_in_flit_0_valid),
    .io_in_flit_0_bits_head(monitor_1_io_in_flit_0_bits_head),
    .io_in_flit_0_bits_tail(monitor_1_io_in_flit_0_bits_tail),
    .io_in_flit_0_bits_flow_ingress_node(monitor_1_io_in_flit_0_bits_flow_ingress_node),
    .io_in_flit_0_bits_flow_egress_node(monitor_1_io_in_flit_0_bits_flow_egress_node),
    .io_in_flit_0_bits_virt_channel_id(monitor_1_io_in_flit_0_bits_virt_channel_id)
  );
  InputUnit input_unit_0_from_0 ( // @[Router.scala 112:13]
    .clock(input_unit_0_from_0_clock),
    .reset(input_unit_0_from_0_reset),
    .io_router_req_valid(input_unit_0_from_0_io_router_req_valid),
    .io_router_req_bits_src_virt_id(input_unit_0_from_0_io_router_req_bits_src_virt_id),
    .io_vcalloc_req_ready(input_unit_0_from_0_io_vcalloc_req_ready),
    .io_vcalloc_req_valid(input_unit_0_from_0_io_vcalloc_req_valid),
    .io_vcalloc_req_bits_vc_sel_0_0(input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_0),
    .io_vcalloc_resp_vc_sel_0_0(input_unit_0_from_0_io_vcalloc_resp_vc_sel_0_0),
    .io_out_credit_available_0_0(input_unit_0_from_0_io_out_credit_available_0_0),
    .io_salloc_req_0_ready(input_unit_0_from_0_io_salloc_req_0_ready),
    .io_salloc_req_0_valid(input_unit_0_from_0_io_salloc_req_0_valid),
    .io_salloc_req_0_bits_vc_sel_0_0(input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_0),
    .io_salloc_req_0_bits_tail(input_unit_0_from_0_io_salloc_req_0_bits_tail),
    .io_out_0_valid(input_unit_0_from_0_io_out_0_valid),
    .io_out_0_bits_flit_head(input_unit_0_from_0_io_out_0_bits_flit_head),
    .io_out_0_bits_flit_tail(input_unit_0_from_0_io_out_0_bits_flit_tail),
    .io_out_0_bits_flit_payload(input_unit_0_from_0_io_out_0_bits_flit_payload),
    .io_out_0_bits_flit_flow_ingress_node(input_unit_0_from_0_io_out_0_bits_flit_flow_ingress_node),
    .io_debug_va_stall(input_unit_0_from_0_io_debug_va_stall),
    .io_debug_sa_stall(input_unit_0_from_0_io_debug_sa_stall),
    .io_in_flit_0_valid(input_unit_0_from_0_io_in_flit_0_valid),
    .io_in_flit_0_bits_head(input_unit_0_from_0_io_in_flit_0_bits_head),
    .io_in_flit_0_bits_tail(input_unit_0_from_0_io_in_flit_0_bits_tail),
    .io_in_flit_0_bits_payload(input_unit_0_from_0_io_in_flit_0_bits_payload),
    .io_in_flit_0_bits_flow_ingress_node(input_unit_0_from_0_io_in_flit_0_bits_flow_ingress_node),
    .io_in_flit_0_bits_flow_egress_node(input_unit_0_from_0_io_in_flit_0_bits_flow_egress_node),
    .io_in_flit_0_bits_virt_channel_id(input_unit_0_from_0_io_in_flit_0_bits_virt_channel_id),
    .io_in_credit_return(input_unit_0_from_0_io_in_credit_return),
    .io_in_vc_free(input_unit_0_from_0_io_in_vc_free)
  );
  InputUnit input_unit_1_from_2 ( // @[Router.scala 112:13]
    .clock(input_unit_1_from_2_clock),
    .reset(input_unit_1_from_2_reset),
    .io_router_req_valid(input_unit_1_from_2_io_router_req_valid),
    .io_router_req_bits_src_virt_id(input_unit_1_from_2_io_router_req_bits_src_virt_id),
    .io_vcalloc_req_ready(input_unit_1_from_2_io_vcalloc_req_ready),
    .io_vcalloc_req_valid(input_unit_1_from_2_io_vcalloc_req_valid),
    .io_vcalloc_req_bits_vc_sel_0_0(input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_0_0),
    .io_vcalloc_resp_vc_sel_0_0(input_unit_1_from_2_io_vcalloc_resp_vc_sel_0_0),
    .io_out_credit_available_0_0(input_unit_1_from_2_io_out_credit_available_0_0),
    .io_salloc_req_0_ready(input_unit_1_from_2_io_salloc_req_0_ready),
    .io_salloc_req_0_valid(input_unit_1_from_2_io_salloc_req_0_valid),
    .io_salloc_req_0_bits_vc_sel_0_0(input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_0_0),
    .io_salloc_req_0_bits_tail(input_unit_1_from_2_io_salloc_req_0_bits_tail),
    .io_out_0_valid(input_unit_1_from_2_io_out_0_valid),
    .io_out_0_bits_flit_head(input_unit_1_from_2_io_out_0_bits_flit_head),
    .io_out_0_bits_flit_tail(input_unit_1_from_2_io_out_0_bits_flit_tail),
    .io_out_0_bits_flit_payload(input_unit_1_from_2_io_out_0_bits_flit_payload),
    .io_out_0_bits_flit_flow_ingress_node(input_unit_1_from_2_io_out_0_bits_flit_flow_ingress_node),
    .io_debug_va_stall(input_unit_1_from_2_io_debug_va_stall),
    .io_debug_sa_stall(input_unit_1_from_2_io_debug_sa_stall),
    .io_in_flit_0_valid(input_unit_1_from_2_io_in_flit_0_valid),
    .io_in_flit_0_bits_head(input_unit_1_from_2_io_in_flit_0_bits_head),
    .io_in_flit_0_bits_tail(input_unit_1_from_2_io_in_flit_0_bits_tail),
    .io_in_flit_0_bits_payload(input_unit_1_from_2_io_in_flit_0_bits_payload),
    .io_in_flit_0_bits_flow_ingress_node(input_unit_1_from_2_io_in_flit_0_bits_flow_ingress_node),
    .io_in_flit_0_bits_flow_egress_node(input_unit_1_from_2_io_in_flit_0_bits_flow_egress_node),
    .io_in_flit_0_bits_virt_channel_id(input_unit_1_from_2_io_in_flit_0_bits_virt_channel_id),
    .io_in_credit_return(input_unit_1_from_2_io_in_credit_return),
    .io_in_vc_free(input_unit_1_from_2_io_in_vc_free)
  );
  EgressUnit egress_unit_0_to_0 ( // @[Router.scala 125:13]
    .clock(egress_unit_0_to_0_clock),
    .reset(egress_unit_0_to_0_reset),
    .io_in_0_valid(egress_unit_0_to_0_io_in_0_valid),
    .io_in_0_bits_head(egress_unit_0_to_0_io_in_0_bits_head),
    .io_in_0_bits_tail(egress_unit_0_to_0_io_in_0_bits_tail),
    .io_in_0_bits_payload(egress_unit_0_to_0_io_in_0_bits_payload),
    .io_in_0_bits_flow_ingress_node(egress_unit_0_to_0_io_in_0_bits_flow_ingress_node),
    .io_credit_available_0(egress_unit_0_to_0_io_credit_available_0),
    .io_channel_status_0_occupied(egress_unit_0_to_0_io_channel_status_0_occupied),
    .io_allocs_0_alloc(egress_unit_0_to_0_io_allocs_0_alloc),
    .io_credit_alloc_0_alloc(egress_unit_0_to_0_io_credit_alloc_0_alloc),
    .io_credit_alloc_0_tail(egress_unit_0_to_0_io_credit_alloc_0_tail),
    .io_out_valid(egress_unit_0_to_0_io_out_valid),
    .io_out_bits_head(egress_unit_0_to_0_io_out_bits_head),
    .io_out_bits_tail(egress_unit_0_to_0_io_out_bits_tail),
    .io_out_bits_payload(egress_unit_0_to_0_io_out_bits_payload),
    .io_out_bits_ingress_id(egress_unit_0_to_0_io_out_bits_ingress_id)
  );
  Switch_1 switch ( // @[Router.scala 129:24]
    .clock(switch_clock),
    .reset(switch_reset),
    .io_in_1_0_valid(switch_io_in_1_0_valid),
    .io_in_1_0_bits_flit_head(switch_io_in_1_0_bits_flit_head),
    .io_in_1_0_bits_flit_tail(switch_io_in_1_0_bits_flit_tail),
    .io_in_1_0_bits_flit_payload(switch_io_in_1_0_bits_flit_payload),
    .io_in_1_0_bits_flit_flow_ingress_node(switch_io_in_1_0_bits_flit_flow_ingress_node),
    .io_in_0_0_valid(switch_io_in_0_0_valid),
    .io_in_0_0_bits_flit_head(switch_io_in_0_0_bits_flit_head),
    .io_in_0_0_bits_flit_tail(switch_io_in_0_0_bits_flit_tail),
    .io_in_0_0_bits_flit_payload(switch_io_in_0_0_bits_flit_payload),
    .io_in_0_0_bits_flit_flow_ingress_node(switch_io_in_0_0_bits_flit_flow_ingress_node),
    .io_out_0_0_valid(switch_io_out_0_0_valid),
    .io_out_0_0_bits_head(switch_io_out_0_0_bits_head),
    .io_out_0_0_bits_tail(switch_io_out_0_0_bits_tail),
    .io_out_0_0_bits_payload(switch_io_out_0_0_bits_payload),
    .io_out_0_0_bits_flow_ingress_node(switch_io_out_0_0_bits_flow_ingress_node),
    .io_sel_0_0_1_0(switch_io_sel_0_0_1_0),
    .io_sel_0_0_0_0(switch_io_sel_0_0_0_0)
  );
  SwitchAllocator_1 switch_allocator ( // @[Router.scala 130:34]
    .clock(switch_allocator_clock),
    .reset(switch_allocator_reset),
    .io_req_1_0_ready(switch_allocator_io_req_1_0_ready),
    .io_req_1_0_valid(switch_allocator_io_req_1_0_valid),
    .io_req_1_0_bits_vc_sel_0_0(switch_allocator_io_req_1_0_bits_vc_sel_0_0),
    .io_req_1_0_bits_tail(switch_allocator_io_req_1_0_bits_tail),
    .io_req_0_0_ready(switch_allocator_io_req_0_0_ready),
    .io_req_0_0_valid(switch_allocator_io_req_0_0_valid),
    .io_req_0_0_bits_vc_sel_0_0(switch_allocator_io_req_0_0_bits_vc_sel_0_0),
    .io_req_0_0_bits_tail(switch_allocator_io_req_0_0_bits_tail),
    .io_credit_alloc_0_0_alloc(switch_allocator_io_credit_alloc_0_0_alloc),
    .io_credit_alloc_0_0_tail(switch_allocator_io_credit_alloc_0_0_tail),
    .io_switch_sel_0_0_1_0(switch_allocator_io_switch_sel_0_0_1_0),
    .io_switch_sel_0_0_0_0(switch_allocator_io_switch_sel_0_0_0_0)
  );
  RotatingSingleVCAllocator_1 vc_allocator ( // @[Router.scala 131:30]
    .clock(vc_allocator_clock),
    .reset(vc_allocator_reset),
    .io_req_1_ready(vc_allocator_io_req_1_ready),
    .io_req_1_valid(vc_allocator_io_req_1_valid),
    .io_req_1_bits_vc_sel_0_0(vc_allocator_io_req_1_bits_vc_sel_0_0),
    .io_req_0_ready(vc_allocator_io_req_0_ready),
    .io_req_0_valid(vc_allocator_io_req_0_valid),
    .io_req_0_bits_vc_sel_0_0(vc_allocator_io_req_0_bits_vc_sel_0_0),
    .io_resp_1_vc_sel_0_0(vc_allocator_io_resp_1_vc_sel_0_0),
    .io_resp_0_vc_sel_0_0(vc_allocator_io_resp_0_vc_sel_0_0),
    .io_channel_status_0_0_occupied(vc_allocator_io_channel_status_0_0_occupied),
    .io_out_allocs_0_0_alloc(vc_allocator_io_out_allocs_0_0_alloc)
  );
  RouteComputer_1 route_computer ( // @[Router.scala 134:32]
    .clock(route_computer_clock),
    .reset(route_computer_reset),
    .io_req_1_valid(route_computer_io_req_1_valid),
    .io_req_0_valid(route_computer_io_req_0_valid)
  );
  plusarg_reader #(.FORMAT("noc_util_sample_rate=%d"), .DEFAULT(0), .WIDTH(20)) plusarg_reader ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_out)
  );
  assign auto_debug_out_va_stall_0 = input_unit_0_from_0_io_debug_va_stall; // @[Nodes.scala 1212:84 Router.scala 190:92]
  assign auto_debug_out_va_stall_1 = input_unit_1_from_2_io_debug_va_stall; // @[Nodes.scala 1212:84 Router.scala 190:92]
  assign auto_debug_out_sa_stall_0 = input_unit_0_from_0_io_debug_sa_stall; // @[Nodes.scala 1212:84 Router.scala 191:92]
  assign auto_debug_out_sa_stall_1 = input_unit_1_from_2_io_debug_sa_stall; // @[Nodes.scala 1212:84 Router.scala 191:92]
  assign auto_egress_nodes_out_flit_valid = egress_unit_0_to_0_io_out_valid; // @[Nodes.scala 1212:84 Router.scala 144:65]
  assign auto_egress_nodes_out_flit_bits_head = egress_unit_0_to_0_io_out_bits_head; // @[Nodes.scala 1212:84 Router.scala 144:65]
  assign auto_egress_nodes_out_flit_bits_tail = egress_unit_0_to_0_io_out_bits_tail; // @[Nodes.scala 1212:84 Router.scala 144:65]
  assign auto_egress_nodes_out_flit_bits_payload = egress_unit_0_to_0_io_out_bits_payload; // @[Nodes.scala 1212:84 Router.scala 144:65]
  assign auto_egress_nodes_out_flit_bits_ingress_id = egress_unit_0_to_0_io_out_bits_ingress_id; // @[Nodes.scala 1212:84 Router.scala 144:65]
  assign auto_dest_nodes_in_1_credit_return = input_unit_1_from_2_io_in_credit_return; // @[Nodes.scala 1215:84 Router.scala 141:68]
  assign auto_dest_nodes_in_1_vc_free = input_unit_1_from_2_io_in_vc_free; // @[Nodes.scala 1215:84 Router.scala 141:68]
  assign auto_dest_nodes_in_0_credit_return = input_unit_0_from_0_io_in_credit_return; // @[Nodes.scala 1215:84 Router.scala 141:68]
  assign auto_dest_nodes_in_0_vc_free = input_unit_0_from_0_io_in_vc_free; // @[Nodes.scala 1215:84 Router.scala 141:68]
  assign monitor_clock = clock;
  assign monitor_reset = reset;
  assign monitor_io_in_flit_0_valid = auto_dest_nodes_in_0_flit_0_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_io_in_flit_0_bits_head = auto_dest_nodes_in_0_flit_0_bits_head; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_io_in_flit_0_bits_tail = auto_dest_nodes_in_0_flit_0_bits_tail; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_io_in_flit_0_bits_flow_ingress_node = auto_dest_nodes_in_0_flit_0_bits_flow_ingress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_io_in_flit_0_bits_flow_egress_node = auto_dest_nodes_in_0_flit_0_bits_flow_egress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_io_in_flit_0_bits_virt_channel_id = auto_dest_nodes_in_0_flit_0_bits_virt_channel_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_1_clock = clock;
  assign monitor_1_reset = reset;
  assign monitor_1_io_in_flit_0_valid = auto_dest_nodes_in_1_flit_0_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_1_io_in_flit_0_bits_head = auto_dest_nodes_in_1_flit_0_bits_head; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_1_io_in_flit_0_bits_tail = auto_dest_nodes_in_1_flit_0_bits_tail; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_1_io_in_flit_0_bits_flow_ingress_node = auto_dest_nodes_in_1_flit_0_bits_flow_ingress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_1_io_in_flit_0_bits_flow_egress_node = auto_dest_nodes_in_1_flit_0_bits_flow_egress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_1_io_in_flit_0_bits_virt_channel_id = auto_dest_nodes_in_1_flit_0_bits_virt_channel_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_0_clock = clock;
  assign input_unit_0_from_0_reset = reset;
  assign input_unit_0_from_0_io_vcalloc_req_ready = vc_allocator_io_req_0_ready; // @[Router.scala 151:23]
  assign input_unit_0_from_0_io_vcalloc_resp_vc_sel_0_0 = vc_allocator_io_resp_0_vc_sel_0_0; // @[Router.scala 153:39]
  assign input_unit_0_from_0_io_out_credit_available_0_0 = egress_unit_0_to_0_io_credit_available_0; // @[Router.scala 162:42]
  assign input_unit_0_from_0_io_salloc_req_0_ready = switch_allocator_io_req_0_0_ready; // @[Router.scala 165:23]
  assign input_unit_0_from_0_io_in_flit_0_valid = auto_dest_nodes_in_0_flit_0_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_0_io_in_flit_0_bits_head = auto_dest_nodes_in_0_flit_0_bits_head; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_0_io_in_flit_0_bits_tail = auto_dest_nodes_in_0_flit_0_bits_tail; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_0_io_in_flit_0_bits_payload = auto_dest_nodes_in_0_flit_0_bits_payload; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_0_io_in_flit_0_bits_flow_ingress_node = auto_dest_nodes_in_0_flit_0_bits_flow_ingress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_0_io_in_flit_0_bits_flow_egress_node = auto_dest_nodes_in_0_flit_0_bits_flow_egress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_0_io_in_flit_0_bits_virt_channel_id = auto_dest_nodes_in_0_flit_0_bits_virt_channel_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_1_from_2_clock = clock;
  assign input_unit_1_from_2_reset = reset;
  assign input_unit_1_from_2_io_vcalloc_req_ready = vc_allocator_io_req_1_ready; // @[Router.scala 151:23]
  assign input_unit_1_from_2_io_vcalloc_resp_vc_sel_0_0 = vc_allocator_io_resp_1_vc_sel_0_0; // @[Router.scala 153:39]
  assign input_unit_1_from_2_io_out_credit_available_0_0 = egress_unit_0_to_0_io_credit_available_0; // @[Router.scala 162:42]
  assign input_unit_1_from_2_io_salloc_req_0_ready = switch_allocator_io_req_1_0_ready; // @[Router.scala 165:23]
  assign input_unit_1_from_2_io_in_flit_0_valid = auto_dest_nodes_in_1_flit_0_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_1_from_2_io_in_flit_0_bits_head = auto_dest_nodes_in_1_flit_0_bits_head; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_1_from_2_io_in_flit_0_bits_tail = auto_dest_nodes_in_1_flit_0_bits_tail; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_1_from_2_io_in_flit_0_bits_payload = auto_dest_nodes_in_1_flit_0_bits_payload; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_1_from_2_io_in_flit_0_bits_flow_ingress_node = auto_dest_nodes_in_1_flit_0_bits_flow_ingress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_1_from_2_io_in_flit_0_bits_flow_egress_node = auto_dest_nodes_in_1_flit_0_bits_flow_egress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_1_from_2_io_in_flit_0_bits_virt_channel_id = auto_dest_nodes_in_1_flit_0_bits_virt_channel_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign egress_unit_0_to_0_clock = clock;
  assign egress_unit_0_to_0_reset = reset;
  assign egress_unit_0_to_0_io_in_0_valid = switch_io_out_0_0_valid; // @[Router.scala 172:29]
  assign egress_unit_0_to_0_io_in_0_bits_head = switch_io_out_0_0_bits_head; // @[Router.scala 172:29]
  assign egress_unit_0_to_0_io_in_0_bits_tail = switch_io_out_0_0_bits_tail; // @[Router.scala 172:29]
  assign egress_unit_0_to_0_io_in_0_bits_payload = switch_io_out_0_0_bits_payload; // @[Router.scala 172:29]
  assign egress_unit_0_to_0_io_in_0_bits_flow_ingress_node = switch_io_out_0_0_bits_flow_ingress_node; // @[Router.scala 172:29]
  assign egress_unit_0_to_0_io_allocs_0_alloc = vc_allocator_io_out_allocs_0_0_alloc; // @[Router.scala 157:33]
  assign egress_unit_0_to_0_io_credit_alloc_0_alloc = switch_allocator_io_credit_alloc_0_0_alloc; // @[Router.scala 167:39]
  assign egress_unit_0_to_0_io_credit_alloc_0_tail = switch_allocator_io_credit_alloc_0_0_tail; // @[Router.scala 167:39]
  assign switch_clock = clock;
  assign switch_reset = reset;
  assign switch_io_in_1_0_valid = input_unit_1_from_2_io_out_0_valid; // @[Router.scala 170:23]
  assign switch_io_in_1_0_bits_flit_head = input_unit_1_from_2_io_out_0_bits_flit_head; // @[Router.scala 170:23]
  assign switch_io_in_1_0_bits_flit_tail = input_unit_1_from_2_io_out_0_bits_flit_tail; // @[Router.scala 170:23]
  assign switch_io_in_1_0_bits_flit_payload = input_unit_1_from_2_io_out_0_bits_flit_payload; // @[Router.scala 170:23]
  assign switch_io_in_1_0_bits_flit_flow_ingress_node = input_unit_1_from_2_io_out_0_bits_flit_flow_ingress_node; // @[Router.scala 170:23]
  assign switch_io_in_0_0_valid = input_unit_0_from_0_io_out_0_valid; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_head = input_unit_0_from_0_io_out_0_bits_flit_head; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_tail = input_unit_0_from_0_io_out_0_bits_flit_tail; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_payload = input_unit_0_from_0_io_out_0_bits_flit_payload; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_flow_ingress_node = input_unit_0_from_0_io_out_0_bits_flit_flow_ingress_node; // @[Router.scala 170:23]
  assign switch_io_sel_0_0_1_0 = switch_io_sel_REG_0_0_1_0; // @[Router.scala 173:19]
  assign switch_io_sel_0_0_0_0 = switch_io_sel_REG_0_0_0_0; // @[Router.scala 173:19]
  assign switch_allocator_clock = clock;
  assign switch_allocator_reset = reset;
  assign switch_allocator_io_req_1_0_valid = input_unit_1_from_2_io_salloc_req_0_valid; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_vc_sel_0_0 = input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_0_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_tail = input_unit_1_from_2_io_salloc_req_0_bits_tail; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_valid = input_unit_0_from_0_io_salloc_req_0_valid; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_0_0 = input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_tail = input_unit_0_from_0_io_salloc_req_0_bits_tail; // @[Router.scala 165:23]
  assign vc_allocator_clock = clock;
  assign vc_allocator_reset = reset;
  assign vc_allocator_io_req_1_valid = input_unit_1_from_2_io_vcalloc_req_valid; // @[Router.scala 151:23]
  assign vc_allocator_io_req_1_bits_vc_sel_0_0 = input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_0_0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_valid = input_unit_0_from_0_io_vcalloc_req_valid; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_0_0 = input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_0; // @[Router.scala 151:23]
  assign vc_allocator_io_channel_status_0_0_occupied = egress_unit_0_to_0_io_channel_status_0_occupied; // @[Router.scala 159:23]
  assign route_computer_clock = clock;
  assign route_computer_reset = reset;
  assign route_computer_io_req_1_valid = input_unit_1_from_2_io_router_req_valid; // @[Router.scala 146:23]
  assign route_computer_io_req_0_valid = input_unit_0_from_0_io_router_req_valid; // @[Router.scala 146:23]
  always @(posedge clock) begin
    switch_io_sel_REG_0_0_1_0 <= switch_allocator_io_switch_sel_0_0_1_0; // @[Router.scala 176:14]
    switch_io_sel_REG_0_0_0_0 <= switch_allocator_io_switch_sel_0_0_0_0; // @[Router.scala 176:14]
    if (reset) begin // @[Router.scala 193:28]
      debug_tsc <= 64'h0; // @[Router.scala 193:28]
    end else begin
      debug_tsc <= _debug_tsc_T_1; // @[Router.scala 194:15]
    end
    if (reset) begin // @[Router.scala 195:31]
      debug_sample <= 64'h0; // @[Router.scala 195:31]
    end else if (debug_sample == _GEN_4) begin // @[Router.scala 198:47]
      debug_sample <= 64'h0; // @[Router.scala 198:62]
    end else begin
      debug_sample <= _debug_sample_T_1; // @[Router.scala 196:18]
    end
    if (reset) begin // @[Router.scala 201:29]
      util_ctr <= 64'h0; // @[Router.scala 201:29]
    end else begin
      util_ctr <= _util_ctr_T_1; // @[Router.scala 203:16]
    end
    if (reset) begin // @[Router.scala 202:26]
      fired <= 1'h0; // @[Router.scala 202:26]
    end else if (plusarg_reader_out != 20'h0 & _T_2 & fired) begin // @[Router.scala 205:81]
      fired <= auto_dest_nodes_in_0_flit_0_valid; // @[Router.scala 208:15]
    end else begin
      fired <= fired | auto_dest_nodes_in_0_flit_0_valid; // @[Router.scala 204:13]
    end
    if (reset) begin // @[Router.scala 201:29]
      util_ctr_1 <= 64'h0; // @[Router.scala 201:29]
    end else begin
      util_ctr_1 <= _util_ctr_T_3; // @[Router.scala 203:16]
    end
    if (reset) begin // @[Router.scala 202:26]
      fired_1 <= 1'h0; // @[Router.scala 202:26]
    end else if (plusarg_reader_out != 20'h0 & _T_2 & fired_1) begin // @[Router.scala 205:81]
      fired_1 <= auto_dest_nodes_in_1_flit_0_valid; // @[Router.scala 208:15]
    end else begin
      fired_1 <= fired_1 | auto_dest_nodes_in_1_flit_0_valid; // @[Router.scala 204:13]
    end
    if (reset) begin // @[Router.scala 201:29]
      util_ctr_2 <= 64'h0; // @[Router.scala 201:29]
    end else begin
      util_ctr_2 <= _util_ctr_T_5; // @[Router.scala 203:16]
    end
    if (reset) begin // @[Router.scala 202:26]
      fired_2 <= 1'h0; // @[Router.scala 202:26]
    end else if (plusarg_reader_out != 20'h0 & _T_2 & fired_2) begin // @[Router.scala 205:81]
      fired_2 <= x1_flit_valid; // @[Router.scala 208:15]
    end else begin
      fired_2 <= fired_2 | x1_flit_valid; // @[Router.scala 204:13]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8 & ~reset) begin
          $fwrite(32'h80000002,"nocsample %d 0 1 %d\n",debug_tsc,util_ctr); // @[Router.scala 207:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_16 & ~reset) begin
          $fwrite(32'h80000002,"nocsample %d 2 1 %d\n",debug_tsc,util_ctr_1); // @[Router.scala 207:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_25 & ~reset) begin
          $fwrite(32'h80000002,"nocsample %d 1 e0 %d\n",debug_tsc,util_ctr_2); // @[Router.scala 207:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  switch_io_sel_REG_0_0_1_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  switch_io_sel_REG_0_0_0_0 = _RAND_1[0:0];
  _RAND_2 = {2{`RANDOM}};
  debug_tsc = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  debug_sample = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  util_ctr = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  fired = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  util_ctr_1 = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  fired_1 = _RAND_7[0:0];
  _RAND_8 = {2{`RANDOM}};
  util_ctr_2 = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  fired_2 = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ClockSinkDomain_1(
  output [1:0]  auto_routers_debug_out_va_stall_0,
  output [1:0]  auto_routers_debug_out_va_stall_1,
  output [1:0]  auto_routers_debug_out_sa_stall_0,
  output [1:0]  auto_routers_debug_out_sa_stall_1,
  output        auto_routers_egress_nodes_out_flit_valid,
  output        auto_routers_egress_nodes_out_flit_bits_head,
  output        auto_routers_egress_nodes_out_flit_bits_tail,
  output [63:0] auto_routers_egress_nodes_out_flit_bits_payload,
  output        auto_routers_egress_nodes_out_flit_bits_ingress_id,
  input         auto_routers_dest_nodes_in_1_flit_0_valid,
  input         auto_routers_dest_nodes_in_1_flit_0_bits_head,
  input         auto_routers_dest_nodes_in_1_flit_0_bits_tail,
  input  [63:0] auto_routers_dest_nodes_in_1_flit_0_bits_payload,
  input  [1:0]  auto_routers_dest_nodes_in_1_flit_0_bits_flow_ingress_node,
  input  [1:0]  auto_routers_dest_nodes_in_1_flit_0_bits_flow_egress_node,
  input  [1:0]  auto_routers_dest_nodes_in_1_flit_0_bits_virt_channel_id,
  output [3:0]  auto_routers_dest_nodes_in_1_credit_return,
  output [3:0]  auto_routers_dest_nodes_in_1_vc_free,
  input         auto_routers_dest_nodes_in_0_flit_0_valid,
  input         auto_routers_dest_nodes_in_0_flit_0_bits_head,
  input         auto_routers_dest_nodes_in_0_flit_0_bits_tail,
  input  [63:0] auto_routers_dest_nodes_in_0_flit_0_bits_payload,
  input  [1:0]  auto_routers_dest_nodes_in_0_flit_0_bits_flow_ingress_node,
  input  [1:0]  auto_routers_dest_nodes_in_0_flit_0_bits_flow_egress_node,
  input  [1:0]  auto_routers_dest_nodes_in_0_flit_0_bits_virt_channel_id,
  output [3:0]  auto_routers_dest_nodes_in_0_credit_return,
  output [3:0]  auto_routers_dest_nodes_in_0_vc_free,
  input         auto_clock_in_clock,
  input         auto_clock_in_reset
);
  wire  routers_clock; // @[NoC.scala 64:22]
  wire  routers_reset; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_debug_out_va_stall_0; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_debug_out_va_stall_1; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_debug_out_sa_stall_0; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_debug_out_sa_stall_1; // @[NoC.scala 64:22]
  wire  routers_auto_egress_nodes_out_flit_valid; // @[NoC.scala 64:22]
  wire  routers_auto_egress_nodes_out_flit_bits_head; // @[NoC.scala 64:22]
  wire  routers_auto_egress_nodes_out_flit_bits_tail; // @[NoC.scala 64:22]
  wire [63:0] routers_auto_egress_nodes_out_flit_bits_payload; // @[NoC.scala 64:22]
  wire  routers_auto_egress_nodes_out_flit_bits_ingress_id; // @[NoC.scala 64:22]
  wire  routers_auto_dest_nodes_in_1_flit_0_valid; // @[NoC.scala 64:22]
  wire  routers_auto_dest_nodes_in_1_flit_0_bits_head; // @[NoC.scala 64:22]
  wire  routers_auto_dest_nodes_in_1_flit_0_bits_tail; // @[NoC.scala 64:22]
  wire [63:0] routers_auto_dest_nodes_in_1_flit_0_bits_payload; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_dest_nodes_in_1_flit_0_bits_flow_ingress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_dest_nodes_in_1_flit_0_bits_flow_egress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_dest_nodes_in_1_flit_0_bits_virt_channel_id; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_dest_nodes_in_1_credit_return; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_dest_nodes_in_1_vc_free; // @[NoC.scala 64:22]
  wire  routers_auto_dest_nodes_in_0_flit_0_valid; // @[NoC.scala 64:22]
  wire  routers_auto_dest_nodes_in_0_flit_0_bits_head; // @[NoC.scala 64:22]
  wire  routers_auto_dest_nodes_in_0_flit_0_bits_tail; // @[NoC.scala 64:22]
  wire [63:0] routers_auto_dest_nodes_in_0_flit_0_bits_payload; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_dest_nodes_in_0_flit_0_bits_flow_ingress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_dest_nodes_in_0_flit_0_bits_flow_egress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_dest_nodes_in_0_flit_0_bits_virt_channel_id; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_dest_nodes_in_0_credit_return; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_dest_nodes_in_0_vc_free; // @[NoC.scala 64:22]
  Router_1 routers ( // @[NoC.scala 64:22]
    .clock(routers_clock),
    .reset(routers_reset),
    .auto_debug_out_va_stall_0(routers_auto_debug_out_va_stall_0),
    .auto_debug_out_va_stall_1(routers_auto_debug_out_va_stall_1),
    .auto_debug_out_sa_stall_0(routers_auto_debug_out_sa_stall_0),
    .auto_debug_out_sa_stall_1(routers_auto_debug_out_sa_stall_1),
    .auto_egress_nodes_out_flit_valid(routers_auto_egress_nodes_out_flit_valid),
    .auto_egress_nodes_out_flit_bits_head(routers_auto_egress_nodes_out_flit_bits_head),
    .auto_egress_nodes_out_flit_bits_tail(routers_auto_egress_nodes_out_flit_bits_tail),
    .auto_egress_nodes_out_flit_bits_payload(routers_auto_egress_nodes_out_flit_bits_payload),
    .auto_egress_nodes_out_flit_bits_ingress_id(routers_auto_egress_nodes_out_flit_bits_ingress_id),
    .auto_dest_nodes_in_1_flit_0_valid(routers_auto_dest_nodes_in_1_flit_0_valid),
    .auto_dest_nodes_in_1_flit_0_bits_head(routers_auto_dest_nodes_in_1_flit_0_bits_head),
    .auto_dest_nodes_in_1_flit_0_bits_tail(routers_auto_dest_nodes_in_1_flit_0_bits_tail),
    .auto_dest_nodes_in_1_flit_0_bits_payload(routers_auto_dest_nodes_in_1_flit_0_bits_payload),
    .auto_dest_nodes_in_1_flit_0_bits_flow_ingress_node(routers_auto_dest_nodes_in_1_flit_0_bits_flow_ingress_node),
    .auto_dest_nodes_in_1_flit_0_bits_flow_egress_node(routers_auto_dest_nodes_in_1_flit_0_bits_flow_egress_node),
    .auto_dest_nodes_in_1_flit_0_bits_virt_channel_id(routers_auto_dest_nodes_in_1_flit_0_bits_virt_channel_id),
    .auto_dest_nodes_in_1_credit_return(routers_auto_dest_nodes_in_1_credit_return),
    .auto_dest_nodes_in_1_vc_free(routers_auto_dest_nodes_in_1_vc_free),
    .auto_dest_nodes_in_0_flit_0_valid(routers_auto_dest_nodes_in_0_flit_0_valid),
    .auto_dest_nodes_in_0_flit_0_bits_head(routers_auto_dest_nodes_in_0_flit_0_bits_head),
    .auto_dest_nodes_in_0_flit_0_bits_tail(routers_auto_dest_nodes_in_0_flit_0_bits_tail),
    .auto_dest_nodes_in_0_flit_0_bits_payload(routers_auto_dest_nodes_in_0_flit_0_bits_payload),
    .auto_dest_nodes_in_0_flit_0_bits_flow_ingress_node(routers_auto_dest_nodes_in_0_flit_0_bits_flow_ingress_node),
    .auto_dest_nodes_in_0_flit_0_bits_flow_egress_node(routers_auto_dest_nodes_in_0_flit_0_bits_flow_egress_node),
    .auto_dest_nodes_in_0_flit_0_bits_virt_channel_id(routers_auto_dest_nodes_in_0_flit_0_bits_virt_channel_id),
    .auto_dest_nodes_in_0_credit_return(routers_auto_dest_nodes_in_0_credit_return),
    .auto_dest_nodes_in_0_vc_free(routers_auto_dest_nodes_in_0_vc_free)
  );
  assign auto_routers_debug_out_va_stall_0 = routers_auto_debug_out_va_stall_0; // @[LazyModule.scala 368:12]
  assign auto_routers_debug_out_va_stall_1 = routers_auto_debug_out_va_stall_1; // @[LazyModule.scala 368:12]
  assign auto_routers_debug_out_sa_stall_0 = routers_auto_debug_out_sa_stall_0; // @[LazyModule.scala 368:12]
  assign auto_routers_debug_out_sa_stall_1 = routers_auto_debug_out_sa_stall_1; // @[LazyModule.scala 368:12]
  assign auto_routers_egress_nodes_out_flit_valid = routers_auto_egress_nodes_out_flit_valid; // @[LazyModule.scala 368:12]
  assign auto_routers_egress_nodes_out_flit_bits_head = routers_auto_egress_nodes_out_flit_bits_head; // @[LazyModule.scala 368:12]
  assign auto_routers_egress_nodes_out_flit_bits_tail = routers_auto_egress_nodes_out_flit_bits_tail; // @[LazyModule.scala 368:12]
  assign auto_routers_egress_nodes_out_flit_bits_payload = routers_auto_egress_nodes_out_flit_bits_payload; // @[LazyModule.scala 368:12]
  assign auto_routers_egress_nodes_out_flit_bits_ingress_id = routers_auto_egress_nodes_out_flit_bits_ingress_id; // @[LazyModule.scala 368:12]
  assign auto_routers_dest_nodes_in_1_credit_return = routers_auto_dest_nodes_in_1_credit_return; // @[LazyModule.scala 366:16]
  assign auto_routers_dest_nodes_in_1_vc_free = routers_auto_dest_nodes_in_1_vc_free; // @[LazyModule.scala 366:16]
  assign auto_routers_dest_nodes_in_0_credit_return = routers_auto_dest_nodes_in_0_credit_return; // @[LazyModule.scala 366:16]
  assign auto_routers_dest_nodes_in_0_vc_free = routers_auto_dest_nodes_in_0_vc_free; // @[LazyModule.scala 366:16]
  assign routers_clock = auto_clock_in_clock; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign routers_reset = auto_clock_in_reset; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_1_flit_0_valid = auto_routers_dest_nodes_in_1_flit_0_valid; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_1_flit_0_bits_head = auto_routers_dest_nodes_in_1_flit_0_bits_head; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_1_flit_0_bits_tail = auto_routers_dest_nodes_in_1_flit_0_bits_tail; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_1_flit_0_bits_payload = auto_routers_dest_nodes_in_1_flit_0_bits_payload; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_1_flit_0_bits_flow_ingress_node =
    auto_routers_dest_nodes_in_1_flit_0_bits_flow_ingress_node; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_1_flit_0_bits_flow_egress_node =
    auto_routers_dest_nodes_in_1_flit_0_bits_flow_egress_node; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_1_flit_0_bits_virt_channel_id =
    auto_routers_dest_nodes_in_1_flit_0_bits_virt_channel_id; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_0_flit_0_valid = auto_routers_dest_nodes_in_0_flit_0_valid; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_0_flit_0_bits_head = auto_routers_dest_nodes_in_0_flit_0_bits_head; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_0_flit_0_bits_tail = auto_routers_dest_nodes_in_0_flit_0_bits_tail; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_0_flit_0_bits_payload = auto_routers_dest_nodes_in_0_flit_0_bits_payload; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_0_flit_0_bits_flow_ingress_node =
    auto_routers_dest_nodes_in_0_flit_0_bits_flow_ingress_node; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_0_flit_0_bits_flow_egress_node =
    auto_routers_dest_nodes_in_0_flit_0_bits_flow_egress_node; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_0_flit_0_bits_virt_channel_id =
    auto_routers_dest_nodes_in_0_flit_0_bits_virt_channel_id; // @[LazyModule.scala 366:16]
endmodule
module IngressUnit_1(
  input         clock,
  input         reset,
  output        io_router_req_valid,
  output [1:0]  io_router_req_bits_flow_ingress_node,
  output [1:0]  io_router_req_bits_flow_egress_node,
  input         io_router_resp_vc_sel_1_0,
  input         io_router_resp_vc_sel_1_1,
  input         io_router_resp_vc_sel_1_2,
  input         io_router_resp_vc_sel_1_3,
  input         io_router_resp_vc_sel_0_0,
  input         io_router_resp_vc_sel_0_1,
  input         io_router_resp_vc_sel_0_2,
  input         io_router_resp_vc_sel_0_3,
  input         io_vcalloc_req_ready,
  output        io_vcalloc_req_valid,
  output        io_vcalloc_req_bits_vc_sel_1_0,
  output        io_vcalloc_req_bits_vc_sel_1_1,
  output        io_vcalloc_req_bits_vc_sel_1_2,
  output        io_vcalloc_req_bits_vc_sel_1_3,
  output        io_vcalloc_req_bits_vc_sel_0_0,
  output        io_vcalloc_req_bits_vc_sel_0_1,
  output        io_vcalloc_req_bits_vc_sel_0_2,
  output        io_vcalloc_req_bits_vc_sel_0_3,
  input         io_vcalloc_resp_vc_sel_1_0,
  input         io_vcalloc_resp_vc_sel_1_1,
  input         io_vcalloc_resp_vc_sel_1_2,
  input         io_vcalloc_resp_vc_sel_1_3,
  input         io_vcalloc_resp_vc_sel_0_0,
  input         io_vcalloc_resp_vc_sel_0_1,
  input         io_vcalloc_resp_vc_sel_0_2,
  input         io_vcalloc_resp_vc_sel_0_3,
  input         io_out_credit_available_1_1,
  input         io_out_credit_available_1_2,
  input         io_out_credit_available_1_3,
  input         io_out_credit_available_0_1,
  input         io_out_credit_available_0_2,
  input         io_out_credit_available_0_3,
  input         io_salloc_req_0_ready,
  output        io_salloc_req_0_valid,
  output        io_salloc_req_0_bits_vc_sel_1_0,
  output        io_salloc_req_0_bits_vc_sel_1_1,
  output        io_salloc_req_0_bits_vc_sel_1_2,
  output        io_salloc_req_0_bits_vc_sel_1_3,
  output        io_salloc_req_0_bits_vc_sel_0_0,
  output        io_salloc_req_0_bits_vc_sel_0_1,
  output        io_salloc_req_0_bits_vc_sel_0_2,
  output        io_salloc_req_0_bits_vc_sel_0_3,
  output        io_salloc_req_0_bits_tail,
  output        io_out_0_valid,
  output        io_out_0_bits_flit_head,
  output        io_out_0_bits_flit_tail,
  output [63:0] io_out_0_bits_flit_payload,
  output [1:0]  io_out_0_bits_flit_flow_ingress_node,
  output [1:0]  io_out_0_bits_flit_flow_egress_node,
  output [1:0]  io_out_0_bits_out_virt_channel,
  output        io_in_ready,
  input         io_in_valid,
  input         io_in_bits_head,
  input         io_in_bits_tail,
  input  [63:0] io_in_bits_payload,
  input         io_in_bits_egress_id
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  route_buffer_clock; // @[IngressUnit.scala 26:28]
  wire  route_buffer_reset; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_enq_ready; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_enq_valid; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_enq_bits_head; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_enq_bits_tail; // @[IngressUnit.scala 26:28]
  wire [63:0] route_buffer_io_enq_bits_payload; // @[IngressUnit.scala 26:28]
  wire [1:0] route_buffer_io_enq_bits_flow_ingress_node; // @[IngressUnit.scala 26:28]
  wire [1:0] route_buffer_io_enq_bits_flow_egress_node; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_deq_ready; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_deq_valid; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_deq_bits_head; // @[IngressUnit.scala 26:28]
  wire  route_buffer_io_deq_bits_tail; // @[IngressUnit.scala 26:28]
  wire [63:0] route_buffer_io_deq_bits_payload; // @[IngressUnit.scala 26:28]
  wire [1:0] route_buffer_io_deq_bits_flow_ingress_node; // @[IngressUnit.scala 26:28]
  wire [1:0] route_buffer_io_deq_bits_flow_egress_node; // @[IngressUnit.scala 26:28]
  wire  route_q_clock; // @[IngressUnit.scala 27:23]
  wire  route_q_reset; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_ready; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_valid; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_1_0; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_1_1; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_1_2; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_1_3; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_0_0; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_0_1; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_0_2; // @[IngressUnit.scala 27:23]
  wire  route_q_io_enq_bits_vc_sel_0_3; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_ready; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_valid; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_1_0; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_1_1; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_1_2; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_1_3; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_0_0; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_0_1; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_0_2; // @[IngressUnit.scala 27:23]
  wire  route_q_io_deq_bits_vc_sel_0_3; // @[IngressUnit.scala 27:23]
  wire  vcalloc_buffer_clock; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_reset; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_enq_ready; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_enq_valid; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_enq_bits_head; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_enq_bits_tail; // @[IngressUnit.scala 75:30]
  wire [63:0] vcalloc_buffer_io_enq_bits_payload; // @[IngressUnit.scala 75:30]
  wire [1:0] vcalloc_buffer_io_enq_bits_flow_ingress_node; // @[IngressUnit.scala 75:30]
  wire [1:0] vcalloc_buffer_io_enq_bits_flow_egress_node; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_deq_ready; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_deq_valid; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_deq_bits_head; // @[IngressUnit.scala 75:30]
  wire  vcalloc_buffer_io_deq_bits_tail; // @[IngressUnit.scala 75:30]
  wire [63:0] vcalloc_buffer_io_deq_bits_payload; // @[IngressUnit.scala 75:30]
  wire [1:0] vcalloc_buffer_io_deq_bits_flow_ingress_node; // @[IngressUnit.scala 75:30]
  wire [1:0] vcalloc_buffer_io_deq_bits_flow_egress_node; // @[IngressUnit.scala 75:30]
  wire  vcalloc_q_clock; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_reset; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_ready; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_valid; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_1_0; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_1_1; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_1_2; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_1_3; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_0_0; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_0_1; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_0_2; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_enq_bits_vc_sel_0_3; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_ready; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_valid; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_1_0; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_1_1; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_1_2; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_1_3; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_0_0; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_0_1; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_0_2; // @[IngressUnit.scala 76:25]
  wire  vcalloc_q_io_deq_bits_vc_sel_0_3; // @[IngressUnit.scala 76:25]
  wire  _T = ~io_in_bits_egress_id; // @[IngressUnit.scala 30:72]
  wire  _T_2 = _T | io_in_bits_egress_id; // @[package.scala 73:59]
  wire  _T_7 = ~reset; // @[IngressUnit.scala 30:9]
  wire [1:0] _route_buffer_io_enq_bits_flow_egress_node_T_3 = io_in_bits_egress_id ? 2'h3 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _GEN_9 = {{1'd0}, _T}; // @[Mux.scala 27:73]
  wire  at_dest = route_buffer_io_enq_bits_flow_egress_node == 2'h2; // @[IngressUnit.scala 55:59]
  wire  _T_9 = io_in_ready & io_in_valid; // @[Decoupled.scala 51:35]
  wire  _vcalloc_buffer_io_enq_valid_T = ~route_buffer_io_deq_bits_head; // @[IngressUnit.scala 88:30]
  wire  _vcalloc_buffer_io_enq_valid_T_1 = route_q_io_deq_valid | ~route_buffer_io_deq_bits_head; // @[IngressUnit.scala 88:27]
  wire  _vcalloc_buffer_io_enq_valid_T_2 = route_buffer_io_deq_valid & _vcalloc_buffer_io_enq_valid_T_1; // @[IngressUnit.scala 87:61]
  wire  _vcalloc_buffer_io_enq_valid_T_4 = io_vcalloc_req_ready | _vcalloc_buffer_io_enq_valid_T; // @[IngressUnit.scala 89:27]
  wire  _io_vcalloc_req_valid_T_1 = route_buffer_io_deq_valid & route_q_io_deq_valid & route_buffer_io_deq_bits_head; // @[IngressUnit.scala 91:78]
  wire  _route_buffer_io_deq_ready_T_2 = vcalloc_buffer_io_enq_ready & _vcalloc_buffer_io_enq_valid_T_1; // @[IngressUnit.scala 93:61]
  wire  _route_buffer_io_deq_ready_T_5 = _route_buffer_io_deq_ready_T_2 & _vcalloc_buffer_io_enq_valid_T_4; // @[IngressUnit.scala 94:37]
  wire  _route_buffer_io_deq_ready_T_7 = vcalloc_q_io_enq_ready | _vcalloc_buffer_io_enq_valid_T; // @[IngressUnit.scala 96:29]
  wire  _route_q_io_deq_ready_T = route_buffer_io_deq_ready & route_buffer_io_deq_valid; // @[Decoupled.scala 51:35]
  wire [3:0] c_lo = {vcalloc_q_io_deq_bits_vc_sel_0_3,vcalloc_q_io_deq_bits_vc_sel_0_2,vcalloc_q_io_deq_bits_vc_sel_0_1,
    vcalloc_q_io_deq_bits_vc_sel_0_0}; // @[IngressUnit.scala 107:41]
  wire [3:0] c_hi = {vcalloc_q_io_deq_bits_vc_sel_1_3,vcalloc_q_io_deq_bits_vc_sel_1_2,vcalloc_q_io_deq_bits_vc_sel_1_1,
    vcalloc_q_io_deq_bits_vc_sel_1_0}; // @[IngressUnit.scala 107:41]
  wire [7:0] _c_T = {vcalloc_q_io_deq_bits_vc_sel_1_3,vcalloc_q_io_deq_bits_vc_sel_1_2,vcalloc_q_io_deq_bits_vc_sel_1_1,
    vcalloc_q_io_deq_bits_vc_sel_1_0,vcalloc_q_io_deq_bits_vc_sel_0_3,vcalloc_q_io_deq_bits_vc_sel_0_2,
    vcalloc_q_io_deq_bits_vc_sel_0_1,vcalloc_q_io_deq_bits_vc_sel_0_0}; // @[IngressUnit.scala 107:41]
  wire [7:0] _c_T_1 = {io_out_credit_available_1_3,io_out_credit_available_1_2,io_out_credit_available_1_1,1'h1,
    io_out_credit_available_0_3,io_out_credit_available_0_2,io_out_credit_available_0_1,1'h1}; // @[IngressUnit.scala 107:74]
  wire [7:0] _c_T_2 = _c_T & _c_T_1; // @[IngressUnit.scala 107:48]
  wire  c = _c_T_2 != 8'h0; // @[IngressUnit.scala 107:82]
  wire  _vcalloc_q_io_deq_ready_T = vcalloc_buffer_io_deq_ready & vcalloc_buffer_io_deq_valid; // @[Decoupled.scala 51:35]
  reg  out_bundle_valid; // @[IngressUnit.scala 116:8]
  reg  out_bundle_bits_flit_head; // @[IngressUnit.scala 116:8]
  reg  out_bundle_bits_flit_tail; // @[IngressUnit.scala 116:8]
  reg [63:0] out_bundle_bits_flit_payload; // @[IngressUnit.scala 116:8]
  reg [1:0] out_bundle_bits_flit_flow_ingress_node; // @[IngressUnit.scala 116:8]
  reg [1:0] out_bundle_bits_flit_flow_egress_node; // @[IngressUnit.scala 116:8]
  reg [1:0] out_bundle_bits_out_virt_channel; // @[IngressUnit.scala 116:8]
  wire  out_channel_oh_0 = vcalloc_q_io_deq_bits_vc_sel_0_0 | vcalloc_q_io_deq_bits_vc_sel_0_1 |
    vcalloc_q_io_deq_bits_vc_sel_0_2 | vcalloc_q_io_deq_bits_vc_sel_0_3; // @[IngressUnit.scala 123:67]
  wire  out_channel_oh_1 = vcalloc_q_io_deq_bits_vc_sel_1_0 | vcalloc_q_io_deq_bits_vc_sel_1_1 |
    vcalloc_q_io_deq_bits_vc_sel_1_2 | vcalloc_q_io_deq_bits_vc_sel_1_3; // @[IngressUnit.scala 123:67]
  wire [1:0] out_bundle_bits_out_virt_channel_hi_1 = c_lo[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] out_bundle_bits_out_virt_channel_lo_1 = c_lo[1:0]; // @[OneHot.scala 31:18]
  wire  _out_bundle_bits_out_virt_channel_T_1 = |out_bundle_bits_out_virt_channel_hi_1; // @[OneHot.scala 32:14]
  wire [1:0] _out_bundle_bits_out_virt_channel_T_2 = out_bundle_bits_out_virt_channel_hi_1 |
    out_bundle_bits_out_virt_channel_lo_1; // @[OneHot.scala 32:28]
  wire [1:0] _out_bundle_bits_out_virt_channel_T_4 = {_out_bundle_bits_out_virt_channel_T_1,
    _out_bundle_bits_out_virt_channel_T_2[1]}; // @[Cat.scala 33:92]
  wire [1:0] out_bundle_bits_out_virt_channel_hi_3 = c_hi[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] out_bundle_bits_out_virt_channel_lo_3 = c_hi[1:0]; // @[OneHot.scala 31:18]
  wire  _out_bundle_bits_out_virt_channel_T_6 = |out_bundle_bits_out_virt_channel_hi_3; // @[OneHot.scala 32:14]
  wire [1:0] _out_bundle_bits_out_virt_channel_T_7 = out_bundle_bits_out_virt_channel_hi_3 |
    out_bundle_bits_out_virt_channel_lo_3; // @[OneHot.scala 32:28]
  wire [1:0] _out_bundle_bits_out_virt_channel_T_9 = {_out_bundle_bits_out_virt_channel_T_6,
    _out_bundle_bits_out_virt_channel_T_7[1]}; // @[Cat.scala 33:92]
  wire [1:0] _out_bundle_bits_out_virt_channel_T_10 = out_channel_oh_0 ? _out_bundle_bits_out_virt_channel_T_4 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _out_bundle_bits_out_virt_channel_T_11 = out_channel_oh_1 ? _out_bundle_bits_out_virt_channel_T_9 : 2'h0; // @[Mux.scala 27:73]
  Queue route_buffer ( // @[IngressUnit.scala 26:28]
    .clock(route_buffer_clock),
    .reset(route_buffer_reset),
    .io_enq_ready(route_buffer_io_enq_ready),
    .io_enq_valid(route_buffer_io_enq_valid),
    .io_enq_bits_head(route_buffer_io_enq_bits_head),
    .io_enq_bits_tail(route_buffer_io_enq_bits_tail),
    .io_enq_bits_payload(route_buffer_io_enq_bits_payload),
    .io_enq_bits_flow_ingress_node(route_buffer_io_enq_bits_flow_ingress_node),
    .io_enq_bits_flow_egress_node(route_buffer_io_enq_bits_flow_egress_node),
    .io_deq_ready(route_buffer_io_deq_ready),
    .io_deq_valid(route_buffer_io_deq_valid),
    .io_deq_bits_head(route_buffer_io_deq_bits_head),
    .io_deq_bits_tail(route_buffer_io_deq_bits_tail),
    .io_deq_bits_payload(route_buffer_io_deq_bits_payload),
    .io_deq_bits_flow_ingress_node(route_buffer_io_deq_bits_flow_ingress_node),
    .io_deq_bits_flow_egress_node(route_buffer_io_deq_bits_flow_egress_node)
  );
  Queue_1 route_q ( // @[IngressUnit.scala 27:23]
    .clock(route_q_clock),
    .reset(route_q_reset),
    .io_enq_ready(route_q_io_enq_ready),
    .io_enq_valid(route_q_io_enq_valid),
    .io_enq_bits_vc_sel_1_0(route_q_io_enq_bits_vc_sel_1_0),
    .io_enq_bits_vc_sel_1_1(route_q_io_enq_bits_vc_sel_1_1),
    .io_enq_bits_vc_sel_1_2(route_q_io_enq_bits_vc_sel_1_2),
    .io_enq_bits_vc_sel_1_3(route_q_io_enq_bits_vc_sel_1_3),
    .io_enq_bits_vc_sel_0_0(route_q_io_enq_bits_vc_sel_0_0),
    .io_enq_bits_vc_sel_0_1(route_q_io_enq_bits_vc_sel_0_1),
    .io_enq_bits_vc_sel_0_2(route_q_io_enq_bits_vc_sel_0_2),
    .io_enq_bits_vc_sel_0_3(route_q_io_enq_bits_vc_sel_0_3),
    .io_deq_ready(route_q_io_deq_ready),
    .io_deq_valid(route_q_io_deq_valid),
    .io_deq_bits_vc_sel_1_0(route_q_io_deq_bits_vc_sel_1_0),
    .io_deq_bits_vc_sel_1_1(route_q_io_deq_bits_vc_sel_1_1),
    .io_deq_bits_vc_sel_1_2(route_q_io_deq_bits_vc_sel_1_2),
    .io_deq_bits_vc_sel_1_3(route_q_io_deq_bits_vc_sel_1_3),
    .io_deq_bits_vc_sel_0_0(route_q_io_deq_bits_vc_sel_0_0),
    .io_deq_bits_vc_sel_0_1(route_q_io_deq_bits_vc_sel_0_1),
    .io_deq_bits_vc_sel_0_2(route_q_io_deq_bits_vc_sel_0_2),
    .io_deq_bits_vc_sel_0_3(route_q_io_deq_bits_vc_sel_0_3)
  );
  Queue vcalloc_buffer ( // @[IngressUnit.scala 75:30]
    .clock(vcalloc_buffer_clock),
    .reset(vcalloc_buffer_reset),
    .io_enq_ready(vcalloc_buffer_io_enq_ready),
    .io_enq_valid(vcalloc_buffer_io_enq_valid),
    .io_enq_bits_head(vcalloc_buffer_io_enq_bits_head),
    .io_enq_bits_tail(vcalloc_buffer_io_enq_bits_tail),
    .io_enq_bits_payload(vcalloc_buffer_io_enq_bits_payload),
    .io_enq_bits_flow_ingress_node(vcalloc_buffer_io_enq_bits_flow_ingress_node),
    .io_enq_bits_flow_egress_node(vcalloc_buffer_io_enq_bits_flow_egress_node),
    .io_deq_ready(vcalloc_buffer_io_deq_ready),
    .io_deq_valid(vcalloc_buffer_io_deq_valid),
    .io_deq_bits_head(vcalloc_buffer_io_deq_bits_head),
    .io_deq_bits_tail(vcalloc_buffer_io_deq_bits_tail),
    .io_deq_bits_payload(vcalloc_buffer_io_deq_bits_payload),
    .io_deq_bits_flow_ingress_node(vcalloc_buffer_io_deq_bits_flow_ingress_node),
    .io_deq_bits_flow_egress_node(vcalloc_buffer_io_deq_bits_flow_egress_node)
  );
  Queue_3 vcalloc_q ( // @[IngressUnit.scala 76:25]
    .clock(vcalloc_q_clock),
    .reset(vcalloc_q_reset),
    .io_enq_ready(vcalloc_q_io_enq_ready),
    .io_enq_valid(vcalloc_q_io_enq_valid),
    .io_enq_bits_vc_sel_1_0(vcalloc_q_io_enq_bits_vc_sel_1_0),
    .io_enq_bits_vc_sel_1_1(vcalloc_q_io_enq_bits_vc_sel_1_1),
    .io_enq_bits_vc_sel_1_2(vcalloc_q_io_enq_bits_vc_sel_1_2),
    .io_enq_bits_vc_sel_1_3(vcalloc_q_io_enq_bits_vc_sel_1_3),
    .io_enq_bits_vc_sel_0_0(vcalloc_q_io_enq_bits_vc_sel_0_0),
    .io_enq_bits_vc_sel_0_1(vcalloc_q_io_enq_bits_vc_sel_0_1),
    .io_enq_bits_vc_sel_0_2(vcalloc_q_io_enq_bits_vc_sel_0_2),
    .io_enq_bits_vc_sel_0_3(vcalloc_q_io_enq_bits_vc_sel_0_3),
    .io_deq_ready(vcalloc_q_io_deq_ready),
    .io_deq_valid(vcalloc_q_io_deq_valid),
    .io_deq_bits_vc_sel_1_0(vcalloc_q_io_deq_bits_vc_sel_1_0),
    .io_deq_bits_vc_sel_1_1(vcalloc_q_io_deq_bits_vc_sel_1_1),
    .io_deq_bits_vc_sel_1_2(vcalloc_q_io_deq_bits_vc_sel_1_2),
    .io_deq_bits_vc_sel_1_3(vcalloc_q_io_deq_bits_vc_sel_1_3),
    .io_deq_bits_vc_sel_0_0(vcalloc_q_io_deq_bits_vc_sel_0_0),
    .io_deq_bits_vc_sel_0_1(vcalloc_q_io_deq_bits_vc_sel_0_1),
    .io_deq_bits_vc_sel_0_2(vcalloc_q_io_deq_bits_vc_sel_0_2),
    .io_deq_bits_vc_sel_0_3(vcalloc_q_io_deq_bits_vc_sel_0_3)
  );
  assign io_router_req_valid = io_in_valid & route_buffer_io_enq_ready & io_in_bits_head & ~at_dest; // @[IngressUnit.scala 58:86]
  assign io_router_req_bits_flow_ingress_node = route_buffer_io_enq_bits_flow_ingress_node; // @[IngressUnit.scala 53:27]
  assign io_router_req_bits_flow_egress_node = route_buffer_io_enq_bits_flow_egress_node; // @[IngressUnit.scala 53:27]
  assign io_vcalloc_req_valid = _io_vcalloc_req_valid_T_1 & vcalloc_buffer_io_enq_ready & vcalloc_q_io_enq_ready; // @[IngressUnit.scala 92:41]
  assign io_vcalloc_req_bits_vc_sel_1_0 = route_q_io_deq_bits_vc_sel_1_0; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_1_1 = route_q_io_deq_bits_vc_sel_1_1; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_1_2 = route_q_io_deq_bits_vc_sel_1_2; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_1_3 = route_q_io_deq_bits_vc_sel_1_3; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_0_0 = route_q_io_deq_bits_vc_sel_0_0; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_0_1 = route_q_io_deq_bits_vc_sel_0_1; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_0_2 = route_q_io_deq_bits_vc_sel_0_2; // @[IngressUnit.scala 81:30]
  assign io_vcalloc_req_bits_vc_sel_0_3 = route_q_io_deq_bits_vc_sel_0_3; // @[IngressUnit.scala 81:30]
  assign io_salloc_req_0_valid = vcalloc_buffer_io_deq_valid & vcalloc_q_io_deq_valid & c; // @[IngressUnit.scala 109:83]
  assign io_salloc_req_0_bits_vc_sel_1_0 = vcalloc_q_io_deq_bits_vc_sel_1_0; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_1_1 = vcalloc_q_io_deq_bits_vc_sel_1_1; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_1_2 = vcalloc_q_io_deq_bits_vc_sel_1_2; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_1_3 = vcalloc_q_io_deq_bits_vc_sel_1_3; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_0_0 = vcalloc_q_io_deq_bits_vc_sel_0_0; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_0_1 = vcalloc_q_io_deq_bits_vc_sel_0_1; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_0_2 = vcalloc_q_io_deq_bits_vc_sel_0_2; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_vc_sel_0_3 = vcalloc_q_io_deq_bits_vc_sel_0_3; // @[IngressUnit.scala 104:32]
  assign io_salloc_req_0_bits_tail = vcalloc_buffer_io_deq_bits_tail; // @[IngressUnit.scala 105:30]
  assign io_out_0_valid = out_bundle_valid; // @[IngressUnit.scala 118:13]
  assign io_out_0_bits_flit_head = out_bundle_bits_flit_head; // @[IngressUnit.scala 118:13]
  assign io_out_0_bits_flit_tail = out_bundle_bits_flit_tail; // @[IngressUnit.scala 118:13]
  assign io_out_0_bits_flit_payload = out_bundle_bits_flit_payload; // @[IngressUnit.scala 118:13]
  assign io_out_0_bits_flit_flow_ingress_node = out_bundle_bits_flit_flow_ingress_node; // @[IngressUnit.scala 118:13]
  assign io_out_0_bits_flit_flow_egress_node = out_bundle_bits_flit_flow_egress_node; // @[IngressUnit.scala 118:13]
  assign io_out_0_bits_out_virt_channel = out_bundle_bits_out_virt_channel; // @[IngressUnit.scala 118:13]
  assign io_in_ready = route_buffer_io_enq_ready; // @[IngressUnit.scala 59:44]
  assign route_buffer_clock = clock;
  assign route_buffer_reset = reset;
  assign route_buffer_io_enq_valid = io_in_valid; // @[IngressUnit.scala 56:44]
  assign route_buffer_io_enq_bits_head = io_in_bits_head; // @[IngressUnit.scala 32:33]
  assign route_buffer_io_enq_bits_tail = io_in_bits_tail; // @[IngressUnit.scala 33:33]
  assign route_buffer_io_enq_bits_payload = io_in_bits_payload; // @[IngressUnit.scala 50:36]
  assign route_buffer_io_enq_bits_flow_ingress_node = 2'h2; // @[IngressUnit.scala 38:51]
  assign route_buffer_io_enq_bits_flow_egress_node = _GEN_9 | _route_buffer_io_enq_bits_flow_egress_node_T_3; // @[Mux.scala 27:73]
  assign route_buffer_io_deq_ready = _route_buffer_io_deq_ready_T_5 & _route_buffer_io_deq_ready_T_7; // @[IngressUnit.scala 95:37]
  assign route_q_clock = clock;
  assign route_q_reset = reset;
  assign route_q_io_enq_valid = _T_9 & io_in_bits_head & at_dest | io_router_req_valid; // @[IngressUnit.scala 62:24 64:53 65:26]
  assign route_q_io_enq_bits_vc_sel_1_0 = _T_9 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_1_0; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_1_1 = _T_9 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_1_1; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_1_2 = _T_9 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_1_2; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_1_3 = _T_9 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_1_3; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_0_0 = _T_9 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_0_0; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_0_1 = _T_9 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_0_1; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_0_2 = _T_9 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_0_2; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_enq_bits_vc_sel_0_3 = _T_9 & io_in_bits_head & at_dest ? 1'h0 : io_router_resp_vc_sel_0_3; // @[IngressUnit.scala 63:23 64:53 66:52]
  assign route_q_io_deq_ready = _route_q_io_deq_ready_T & route_buffer_io_deq_bits_tail; // @[IngressUnit.scala 97:55]
  assign vcalloc_buffer_clock = clock;
  assign vcalloc_buffer_reset = reset;
  assign vcalloc_buffer_io_enq_valid = _vcalloc_buffer_io_enq_valid_T_2 & _vcalloc_buffer_io_enq_valid_T_4; // @[IngressUnit.scala 88:37]
  assign vcalloc_buffer_io_enq_bits_head = route_buffer_io_deq_bits_head; // @[IngressUnit.scala 79:30]
  assign vcalloc_buffer_io_enq_bits_tail = route_buffer_io_deq_bits_tail; // @[IngressUnit.scala 79:30]
  assign vcalloc_buffer_io_enq_bits_payload = route_buffer_io_deq_bits_payload; // @[IngressUnit.scala 79:30]
  assign vcalloc_buffer_io_enq_bits_flow_ingress_node = route_buffer_io_deq_bits_flow_ingress_node; // @[IngressUnit.scala 79:30]
  assign vcalloc_buffer_io_enq_bits_flow_egress_node = route_buffer_io_deq_bits_flow_egress_node; // @[IngressUnit.scala 79:30]
  assign vcalloc_buffer_io_deq_ready = io_salloc_req_0_ready & vcalloc_q_io_deq_valid & c; // @[IngressUnit.scala 110:83]
  assign vcalloc_q_clock = clock;
  assign vcalloc_q_reset = reset;
  assign vcalloc_q_io_enq_valid = io_vcalloc_req_ready & io_vcalloc_req_valid; // @[Decoupled.scala 51:35]
  assign vcalloc_q_io_enq_bits_vc_sel_1_0 = io_vcalloc_resp_vc_sel_1_0; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_1_1 = io_vcalloc_resp_vc_sel_1_1; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_1_2 = io_vcalloc_resp_vc_sel_1_2; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_1_3 = io_vcalloc_resp_vc_sel_1_3; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_0_0 = io_vcalloc_resp_vc_sel_0_0; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_0_1 = io_vcalloc_resp_vc_sel_0_1; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_0_2 = io_vcalloc_resp_vc_sel_0_2; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_enq_bits_vc_sel_0_3 = io_vcalloc_resp_vc_sel_0_3; // @[IngressUnit.scala 101:25]
  assign vcalloc_q_io_deq_ready = vcalloc_buffer_io_deq_bits_tail & _vcalloc_q_io_deq_ready_T; // @[IngressUnit.scala 111:42]
  always @(posedge clock) begin
    out_bundle_valid <= vcalloc_buffer_io_deq_ready & vcalloc_buffer_io_deq_valid; // @[Decoupled.scala 51:35]
    out_bundle_bits_flit_head <= vcalloc_buffer_io_deq_bits_head; // @[IngressUnit.scala 121:24]
    out_bundle_bits_flit_tail <= vcalloc_buffer_io_deq_bits_tail; // @[IngressUnit.scala 121:24]
    out_bundle_bits_flit_payload <= vcalloc_buffer_io_deq_bits_payload; // @[IngressUnit.scala 121:24]
    out_bundle_bits_flit_flow_ingress_node <= vcalloc_buffer_io_deq_bits_flow_ingress_node; // @[IngressUnit.scala 121:24]
    out_bundle_bits_flit_flow_egress_node <= vcalloc_buffer_io_deq_bits_flow_egress_node; // @[IngressUnit.scala 121:24]
    out_bundle_bits_out_virt_channel <= _out_bundle_bits_out_virt_channel_T_10 | _out_bundle_bits_out_virt_channel_T_11; // @[Mux.scala 27:73]
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~(io_in_valid & ~_T_2))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at IngressUnit.scala:30 assert(!(io.in.valid && !cParam.possibleFlows.toSeq.map(_.egressId.U === io.in.bits.egress_id).orR))\n"
            ); // @[IngressUnit.scala 30:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7 & ~(~(route_q_io_enq_valid & ~route_q_io_enq_ready))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at IngressUnit.scala:73 assert(!(route_q.io.enq.valid && !route_q.io.enq.ready))\n"); // @[IngressUnit.scala 73:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7 & ~(~(vcalloc_q_io_enq_valid & ~vcalloc_q_io_enq_ready))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at IngressUnit.scala:102 assert(!(vcalloc_q.io.enq.valid && !vcalloc_q.io.enq.ready))\n"
            ); // @[IngressUnit.scala 102:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  out_bundle_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  out_bundle_bits_flit_head = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  out_bundle_bits_flit_tail = _RAND_2[0:0];
  _RAND_3 = {2{`RANDOM}};
  out_bundle_bits_flit_payload = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  out_bundle_bits_flit_flow_ingress_node = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  out_bundle_bits_flit_flow_egress_node = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  out_bundle_bits_out_virt_channel = _RAND_6[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(~(io_in_valid & ~_T_2)); // @[IngressUnit.scala 30:9]
    end
    //
    if (_T_7) begin
      assert(~(route_q_io_enq_valid & ~route_q_io_enq_ready)); // @[IngressUnit.scala 73:9]
    end
    //
    if (_T_7) begin
      assert(~(vcalloc_q_io_enq_valid & ~vcalloc_q_io_enq_ready)); // @[IngressUnit.scala 102:9]
    end
  end
endmodule
module RouteComputer_2(
  input  [1:0] io_req_0_bits_flow_ingress_node,
  input  [1:0] io_req_0_bits_flow_egress_node,
  output       io_resp_0_vc_sel_1_0,
  output       io_resp_0_vc_sel_1_1,
  output       io_resp_0_vc_sel_1_2,
  output       io_resp_0_vc_sel_1_3,
  output       io_resp_0_vc_sel_0_0,
  output       io_resp_0_vc_sel_0_1,
  output       io_resp_0_vc_sel_0_2,
  output       io_resp_0_vc_sel_0_3
);
  wire [5:0] addr = {2'h0,io_req_0_bits_flow_ingress_node,io_req_0_bits_flow_egress_node}; // @[RouteComputer.scala 74:27]
  wire [5:0] decoded_invInputs = ~addr; // @[pla.scala 78:21]
  wire  decoded_andMatrixInput_0 = decoded_invInputs[1]; // @[pla.scala 91:29]
  wire  decoded_andMatrixInput_1 = decoded_invInputs[2]; // @[pla.scala 91:29]
  wire  decoded_andMatrixInput_2 = addr[3]; // @[pla.scala 90:45]
  wire  decoded_andMatrixInput_3 = decoded_invInputs[4]; // @[pla.scala 91:29]
  wire  decoded_andMatrixInput_4 = decoded_invInputs[5]; // @[pla.scala 91:29]
  wire [4:0] _decoded_T = {decoded_andMatrixInput_0,decoded_andMatrixInput_1,decoded_andMatrixInput_2,
    decoded_andMatrixInput_3,decoded_andMatrixInput_4}; // @[Cat.scala 33:92]
  wire  _decoded_T_1 = &_decoded_T; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_0_1 = addr[1]; // @[pla.scala 90:45]
  wire [4:0] _decoded_T_2 = {decoded_andMatrixInput_0_1,decoded_andMatrixInput_1,decoded_andMatrixInput_2,
    decoded_andMatrixInput_3,decoded_andMatrixInput_4}; // @[Cat.scala 33:92]
  wire  _decoded_T_3 = &_decoded_T_2; // @[pla.scala 98:74]
  wire  _decoded_orMatrixOutputs_T = |_decoded_T_3; // @[pla.scala 114:39]
  wire  _decoded_orMatrixOutputs_T_3 = |_decoded_T_1; // @[pla.scala 114:39]
  wire [7:0] decoded_orMatrixOutputs = {1'h0,_decoded_orMatrixOutputs_T_3,_decoded_orMatrixOutputs_T_3,
    _decoded_orMatrixOutputs_T_3,1'h0,_decoded_orMatrixOutputs_T,_decoded_orMatrixOutputs_T,_decoded_orMatrixOutputs_T}; // @[Cat.scala 33:92]
  wire [7:0] decoded_invMatrixOutputs = {decoded_orMatrixOutputs[7],decoded_orMatrixOutputs[6],decoded_orMatrixOutputs[5
    ],decoded_orMatrixOutputs[4],decoded_orMatrixOutputs[3],decoded_orMatrixOutputs[2],decoded_orMatrixOutputs[1],
    decoded_orMatrixOutputs[0]}; // @[Cat.scala 33:92]
  wire [7:0] _GEN_0 = {{4'd0}, decoded_invMatrixOutputs[7:4]}; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_7 = _GEN_0 & 8'hf; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_9 = {decoded_invMatrixOutputs[3:0], 4'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _decoded_T_11 = _decoded_T_9 & 8'hf0; // @[Bitwise.scala 108:80]
  wire [7:0] _decoded_T_12 = _decoded_T_7 | _decoded_T_11; // @[Bitwise.scala 108:39]
  wire [7:0] _GEN_1 = {{2'd0}, _decoded_T_12[7:2]}; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_17 = _GEN_1 & 8'h33; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_19 = {_decoded_T_12[5:0], 2'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _decoded_T_21 = _decoded_T_19 & 8'hcc; // @[Bitwise.scala 108:80]
  wire [7:0] _decoded_T_22 = _decoded_T_17 | _decoded_T_21; // @[Bitwise.scala 108:39]
  wire [7:0] _GEN_2 = {{1'd0}, _decoded_T_22[7:1]}; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_27 = _GEN_2 & 8'h55; // @[Bitwise.scala 108:31]
  wire [7:0] _decoded_T_29 = {_decoded_T_22[6:0], 1'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _decoded_T_31 = _decoded_T_29 & 8'haa; // @[Bitwise.scala 108:80]
  wire [7:0] decoded = _decoded_T_27 | _decoded_T_31; // @[Bitwise.scala 108:39]
  assign io_resp_0_vc_sel_1_0 = decoded[4]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_1_1 = decoded[5]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_1_2 = decoded[6]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_1_3 = decoded[7]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_0_0 = decoded[0]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_0_1 = decoded[1]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_0_2 = decoded[2]; // @[RouteComputer.scala 90:46]
  assign io_resp_0_vc_sel_0_3 = decoded[3]; // @[RouteComputer.scala 90:46]
endmodule
module Router_2(
  input         clock,
  input         reset,
  output        auto_ingress_nodes_in_flit_ready,
  input         auto_ingress_nodes_in_flit_valid,
  input         auto_ingress_nodes_in_flit_bits_head,
  input         auto_ingress_nodes_in_flit_bits_tail,
  input  [63:0] auto_ingress_nodes_in_flit_bits_payload,
  input         auto_ingress_nodes_in_flit_bits_egress_id,
  output        auto_source_nodes_out_1_flit_0_valid,
  output        auto_source_nodes_out_1_flit_0_bits_head,
  output        auto_source_nodes_out_1_flit_0_bits_tail,
  output [63:0] auto_source_nodes_out_1_flit_0_bits_payload,
  output [1:0]  auto_source_nodes_out_1_flit_0_bits_flow_ingress_node,
  output [1:0]  auto_source_nodes_out_1_flit_0_bits_flow_egress_node,
  output [1:0]  auto_source_nodes_out_1_flit_0_bits_virt_channel_id,
  input  [3:0]  auto_source_nodes_out_1_credit_return,
  input  [3:0]  auto_source_nodes_out_1_vc_free,
  output        auto_source_nodes_out_0_flit_0_valid,
  output        auto_source_nodes_out_0_flit_0_bits_head,
  output        auto_source_nodes_out_0_flit_0_bits_tail,
  output [63:0] auto_source_nodes_out_0_flit_0_bits_payload,
  output [1:0]  auto_source_nodes_out_0_flit_0_bits_flow_ingress_node,
  output [1:0]  auto_source_nodes_out_0_flit_0_bits_flow_egress_node,
  output [1:0]  auto_source_nodes_out_0_flit_0_bits_virt_channel_id,
  input  [3:0]  auto_source_nodes_out_0_credit_return,
  input  [3:0]  auto_source_nodes_out_0_vc_free
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire  ingress_unit_0_from_1_clock; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_reset; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_router_req_valid; // @[Router.scala 116:13]
  wire [1:0] ingress_unit_0_from_1_io_router_req_bits_flow_ingress_node; // @[Router.scala 116:13]
  wire [1:0] ingress_unit_0_from_1_io_router_req_bits_flow_egress_node; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_router_resp_vc_sel_1_0; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_router_resp_vc_sel_1_1; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_router_resp_vc_sel_1_2; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_router_resp_vc_sel_1_3; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_router_resp_vc_sel_0_0; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_router_resp_vc_sel_0_1; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_router_resp_vc_sel_0_2; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_router_resp_vc_sel_0_3; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_vcalloc_req_ready; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_vcalloc_req_valid; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_vcalloc_req_bits_vc_sel_1_0; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_vcalloc_req_bits_vc_sel_1_1; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_vcalloc_req_bits_vc_sel_1_2; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_vcalloc_req_bits_vc_sel_1_3; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_vcalloc_req_bits_vc_sel_0_0; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_vcalloc_req_bits_vc_sel_0_1; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_vcalloc_req_bits_vc_sel_0_2; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_vcalloc_req_bits_vc_sel_0_3; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_vcalloc_resp_vc_sel_1_0; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_vcalloc_resp_vc_sel_1_1; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_vcalloc_resp_vc_sel_1_2; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_vcalloc_resp_vc_sel_1_3; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_vcalloc_resp_vc_sel_0_0; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_vcalloc_resp_vc_sel_0_1; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_vcalloc_resp_vc_sel_0_2; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_vcalloc_resp_vc_sel_0_3; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_out_credit_available_1_1; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_out_credit_available_1_2; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_out_credit_available_1_3; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_out_credit_available_0_1; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_out_credit_available_0_2; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_out_credit_available_0_3; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_salloc_req_0_ready; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_salloc_req_0_valid; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_salloc_req_0_bits_vc_sel_1_0; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_salloc_req_0_bits_vc_sel_1_1; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_salloc_req_0_bits_vc_sel_1_2; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_salloc_req_0_bits_vc_sel_1_3; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_salloc_req_0_bits_vc_sel_0_0; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_salloc_req_0_bits_vc_sel_0_1; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_salloc_req_0_bits_vc_sel_0_2; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_salloc_req_0_bits_vc_sel_0_3; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_salloc_req_0_bits_tail; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_out_0_valid; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_out_0_bits_flit_head; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_out_0_bits_flit_tail; // @[Router.scala 116:13]
  wire [63:0] ingress_unit_0_from_1_io_out_0_bits_flit_payload; // @[Router.scala 116:13]
  wire [1:0] ingress_unit_0_from_1_io_out_0_bits_flit_flow_ingress_node; // @[Router.scala 116:13]
  wire [1:0] ingress_unit_0_from_1_io_out_0_bits_flit_flow_egress_node; // @[Router.scala 116:13]
  wire [1:0] ingress_unit_0_from_1_io_out_0_bits_out_virt_channel; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_in_ready; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_in_valid; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_in_bits_head; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_in_bits_tail; // @[Router.scala 116:13]
  wire [63:0] ingress_unit_0_from_1_io_in_bits_payload; // @[Router.scala 116:13]
  wire  ingress_unit_0_from_1_io_in_bits_egress_id; // @[Router.scala 116:13]
  wire  output_unit_0_to_1_clock; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_reset; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_in_0_valid; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_in_0_bits_head; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_in_0_bits_tail; // @[Router.scala 122:13]
  wire [63:0] output_unit_0_to_1_io_in_0_bits_payload; // @[Router.scala 122:13]
  wire [1:0] output_unit_0_to_1_io_in_0_bits_flow_ingress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_0_to_1_io_in_0_bits_flow_egress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_0_to_1_io_in_0_bits_virt_channel_id; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_credit_available_1; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_credit_available_2; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_credit_available_3; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_channel_status_1_occupied; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_channel_status_2_occupied; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_channel_status_3_occupied; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_allocs_1_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_allocs_2_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_allocs_3_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_credit_alloc_1_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_credit_alloc_2_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_credit_alloc_3_alloc; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_out_flit_0_valid; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_out_flit_0_bits_head; // @[Router.scala 122:13]
  wire  output_unit_0_to_1_io_out_flit_0_bits_tail; // @[Router.scala 122:13]
  wire [63:0] output_unit_0_to_1_io_out_flit_0_bits_payload; // @[Router.scala 122:13]
  wire [1:0] output_unit_0_to_1_io_out_flit_0_bits_flow_ingress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_0_to_1_io_out_flit_0_bits_flow_egress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_0_to_1_io_out_flit_0_bits_virt_channel_id; // @[Router.scala 122:13]
  wire [3:0] output_unit_0_to_1_io_out_credit_return; // @[Router.scala 122:13]
  wire [3:0] output_unit_0_to_1_io_out_vc_free; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_clock; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_reset; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_in_0_valid; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_in_0_bits_head; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_in_0_bits_tail; // @[Router.scala 122:13]
  wire [63:0] output_unit_1_to_3_io_in_0_bits_payload; // @[Router.scala 122:13]
  wire [1:0] output_unit_1_to_3_io_in_0_bits_flow_ingress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_1_to_3_io_in_0_bits_flow_egress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_1_to_3_io_in_0_bits_virt_channel_id; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_credit_available_1; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_credit_available_2; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_credit_available_3; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_channel_status_1_occupied; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_channel_status_2_occupied; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_channel_status_3_occupied; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_allocs_1_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_allocs_2_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_allocs_3_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_credit_alloc_1_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_credit_alloc_2_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_credit_alloc_3_alloc; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_out_flit_0_valid; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_out_flit_0_bits_head; // @[Router.scala 122:13]
  wire  output_unit_1_to_3_io_out_flit_0_bits_tail; // @[Router.scala 122:13]
  wire [63:0] output_unit_1_to_3_io_out_flit_0_bits_payload; // @[Router.scala 122:13]
  wire [1:0] output_unit_1_to_3_io_out_flit_0_bits_flow_ingress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_1_to_3_io_out_flit_0_bits_flow_egress_node; // @[Router.scala 122:13]
  wire [1:0] output_unit_1_to_3_io_out_flit_0_bits_virt_channel_id; // @[Router.scala 122:13]
  wire [3:0] output_unit_1_to_3_io_out_credit_return; // @[Router.scala 122:13]
  wire [3:0] output_unit_1_to_3_io_out_vc_free; // @[Router.scala 122:13]
  wire  switch_clock; // @[Router.scala 129:24]
  wire  switch_reset; // @[Router.scala 129:24]
  wire  switch_io_in_0_0_valid; // @[Router.scala 129:24]
  wire  switch_io_in_0_0_bits_flit_head; // @[Router.scala 129:24]
  wire  switch_io_in_0_0_bits_flit_tail; // @[Router.scala 129:24]
  wire [63:0] switch_io_in_0_0_bits_flit_payload; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_0_0_bits_flit_flow_ingress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_0_0_bits_flit_flow_egress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_0_0_bits_out_virt_channel; // @[Router.scala 129:24]
  wire  switch_io_out_1_0_valid; // @[Router.scala 129:24]
  wire  switch_io_out_1_0_bits_head; // @[Router.scala 129:24]
  wire  switch_io_out_1_0_bits_tail; // @[Router.scala 129:24]
  wire [63:0] switch_io_out_1_0_bits_payload; // @[Router.scala 129:24]
  wire [1:0] switch_io_out_1_0_bits_flow_ingress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_out_1_0_bits_flow_egress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_out_1_0_bits_virt_channel_id; // @[Router.scala 129:24]
  wire  switch_io_out_0_0_valid; // @[Router.scala 129:24]
  wire  switch_io_out_0_0_bits_head; // @[Router.scala 129:24]
  wire  switch_io_out_0_0_bits_tail; // @[Router.scala 129:24]
  wire [63:0] switch_io_out_0_0_bits_payload; // @[Router.scala 129:24]
  wire [1:0] switch_io_out_0_0_bits_flow_ingress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_out_0_0_bits_flow_egress_node; // @[Router.scala 129:24]
  wire [1:0] switch_io_out_0_0_bits_virt_channel_id; // @[Router.scala 129:24]
  wire  switch_io_sel_1_0_0_0; // @[Router.scala 129:24]
  wire  switch_io_sel_0_0_0_0; // @[Router.scala 129:24]
  wire  switch_allocator_clock; // @[Router.scala 130:34]
  wire  switch_allocator_reset; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_ready; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_valid; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_1_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_1_1; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_1_2; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_1_3; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_0_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_0_1; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_0_2; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_0_3; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_tail; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_1_1_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_1_2_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_1_3_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_0_1_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_0_2_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_0_3_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_1_0_0_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_0_0_0_0; // @[Router.scala 130:34]
  wire  vc_allocator_clock; // @[Router.scala 131:30]
  wire  vc_allocator_reset; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_ready; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_valid; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_1_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_1_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_1_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_1_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_0_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_0_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_0_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_0_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_1_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_1_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_1_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_1_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_0_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_0_1; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_0_2; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_0_3; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_1_1_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_1_2_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_1_3_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_0_1_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_0_2_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_0_3_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_1_1_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_1_2_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_1_3_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_0_1_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_0_2_alloc; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_0_3_alloc; // @[Router.scala 131:30]
  wire [1:0] route_computer_io_req_0_bits_flow_ingress_node; // @[Router.scala 134:32]
  wire [1:0] route_computer_io_req_0_bits_flow_egress_node; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_1_0; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_1_1; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_1_2; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_1_3; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_0_0; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_0_1; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_0_2; // @[Router.scala 134:32]
  wire  route_computer_io_resp_0_vc_sel_0_3; // @[Router.scala 134:32]
  wire [19:0] plusarg_reader_out; // @[PlusArg.scala 80:11]
  reg  switch_io_sel_REG_1_0_0_0; // @[Router.scala 176:14]
  reg  switch_io_sel_REG_0_0_0_0; // @[Router.scala 176:14]
  reg [63:0] debug_tsc; // @[Router.scala 193:28]
  wire [63:0] _debug_tsc_T_1 = debug_tsc + 64'h1; // @[Router.scala 194:28]
  reg [63:0] debug_sample; // @[Router.scala 195:31]
  wire [63:0] _debug_sample_T_1 = debug_sample + 64'h1; // @[Router.scala 196:34]
  wire [19:0] _T_1 = plusarg_reader_out - 20'h1; // @[Router.scala 198:40]
  wire [63:0] _GEN_2 = {{44'd0}, _T_1}; // @[Router.scala 198:24]
  wire  _T_2 = debug_sample == _GEN_2; // @[Router.scala 198:24]
  wire  bundleIn_0_flit_ready = ingress_unit_0_from_1_io_in_ready; // @[Nodes.scala 1215:84 Router.scala 142:68]
  wire  _T_3 = bundleIn_0_flit_ready & auto_ingress_nodes_in_flit_valid; // @[Decoupled.scala 51:35]
  reg [63:0] util_ctr; // @[Router.scala 201:29]
  reg  fired; // @[Router.scala 202:26]
  wire [63:0] _GEN_3 = {{63'd0}, _T_3}; // @[Router.scala 203:28]
  wire [63:0] _util_ctr_T_1 = util_ctr + _GEN_3; // @[Router.scala 203:28]
  wire  _T_9 = plusarg_reader_out != 20'h0 & _T_2 & fired; // @[Router.scala 205:71]
  wire  fires_count = vc_allocator_io_req_0_ready & vc_allocator_io_req_0_valid; // @[Decoupled.scala 51:35]
  IngressUnit_1 ingress_unit_0_from_1 ( // @[Router.scala 116:13]
    .clock(ingress_unit_0_from_1_clock),
    .reset(ingress_unit_0_from_1_reset),
    .io_router_req_valid(ingress_unit_0_from_1_io_router_req_valid),
    .io_router_req_bits_flow_ingress_node(ingress_unit_0_from_1_io_router_req_bits_flow_ingress_node),
    .io_router_req_bits_flow_egress_node(ingress_unit_0_from_1_io_router_req_bits_flow_egress_node),
    .io_router_resp_vc_sel_1_0(ingress_unit_0_from_1_io_router_resp_vc_sel_1_0),
    .io_router_resp_vc_sel_1_1(ingress_unit_0_from_1_io_router_resp_vc_sel_1_1),
    .io_router_resp_vc_sel_1_2(ingress_unit_0_from_1_io_router_resp_vc_sel_1_2),
    .io_router_resp_vc_sel_1_3(ingress_unit_0_from_1_io_router_resp_vc_sel_1_3),
    .io_router_resp_vc_sel_0_0(ingress_unit_0_from_1_io_router_resp_vc_sel_0_0),
    .io_router_resp_vc_sel_0_1(ingress_unit_0_from_1_io_router_resp_vc_sel_0_1),
    .io_router_resp_vc_sel_0_2(ingress_unit_0_from_1_io_router_resp_vc_sel_0_2),
    .io_router_resp_vc_sel_0_3(ingress_unit_0_from_1_io_router_resp_vc_sel_0_3),
    .io_vcalloc_req_ready(ingress_unit_0_from_1_io_vcalloc_req_ready),
    .io_vcalloc_req_valid(ingress_unit_0_from_1_io_vcalloc_req_valid),
    .io_vcalloc_req_bits_vc_sel_1_0(ingress_unit_0_from_1_io_vcalloc_req_bits_vc_sel_1_0),
    .io_vcalloc_req_bits_vc_sel_1_1(ingress_unit_0_from_1_io_vcalloc_req_bits_vc_sel_1_1),
    .io_vcalloc_req_bits_vc_sel_1_2(ingress_unit_0_from_1_io_vcalloc_req_bits_vc_sel_1_2),
    .io_vcalloc_req_bits_vc_sel_1_3(ingress_unit_0_from_1_io_vcalloc_req_bits_vc_sel_1_3),
    .io_vcalloc_req_bits_vc_sel_0_0(ingress_unit_0_from_1_io_vcalloc_req_bits_vc_sel_0_0),
    .io_vcalloc_req_bits_vc_sel_0_1(ingress_unit_0_from_1_io_vcalloc_req_bits_vc_sel_0_1),
    .io_vcalloc_req_bits_vc_sel_0_2(ingress_unit_0_from_1_io_vcalloc_req_bits_vc_sel_0_2),
    .io_vcalloc_req_bits_vc_sel_0_3(ingress_unit_0_from_1_io_vcalloc_req_bits_vc_sel_0_3),
    .io_vcalloc_resp_vc_sel_1_0(ingress_unit_0_from_1_io_vcalloc_resp_vc_sel_1_0),
    .io_vcalloc_resp_vc_sel_1_1(ingress_unit_0_from_1_io_vcalloc_resp_vc_sel_1_1),
    .io_vcalloc_resp_vc_sel_1_2(ingress_unit_0_from_1_io_vcalloc_resp_vc_sel_1_2),
    .io_vcalloc_resp_vc_sel_1_3(ingress_unit_0_from_1_io_vcalloc_resp_vc_sel_1_3),
    .io_vcalloc_resp_vc_sel_0_0(ingress_unit_0_from_1_io_vcalloc_resp_vc_sel_0_0),
    .io_vcalloc_resp_vc_sel_0_1(ingress_unit_0_from_1_io_vcalloc_resp_vc_sel_0_1),
    .io_vcalloc_resp_vc_sel_0_2(ingress_unit_0_from_1_io_vcalloc_resp_vc_sel_0_2),
    .io_vcalloc_resp_vc_sel_0_3(ingress_unit_0_from_1_io_vcalloc_resp_vc_sel_0_3),
    .io_out_credit_available_1_1(ingress_unit_0_from_1_io_out_credit_available_1_1),
    .io_out_credit_available_1_2(ingress_unit_0_from_1_io_out_credit_available_1_2),
    .io_out_credit_available_1_3(ingress_unit_0_from_1_io_out_credit_available_1_3),
    .io_out_credit_available_0_1(ingress_unit_0_from_1_io_out_credit_available_0_1),
    .io_out_credit_available_0_2(ingress_unit_0_from_1_io_out_credit_available_0_2),
    .io_out_credit_available_0_3(ingress_unit_0_from_1_io_out_credit_available_0_3),
    .io_salloc_req_0_ready(ingress_unit_0_from_1_io_salloc_req_0_ready),
    .io_salloc_req_0_valid(ingress_unit_0_from_1_io_salloc_req_0_valid),
    .io_salloc_req_0_bits_vc_sel_1_0(ingress_unit_0_from_1_io_salloc_req_0_bits_vc_sel_1_0),
    .io_salloc_req_0_bits_vc_sel_1_1(ingress_unit_0_from_1_io_salloc_req_0_bits_vc_sel_1_1),
    .io_salloc_req_0_bits_vc_sel_1_2(ingress_unit_0_from_1_io_salloc_req_0_bits_vc_sel_1_2),
    .io_salloc_req_0_bits_vc_sel_1_3(ingress_unit_0_from_1_io_salloc_req_0_bits_vc_sel_1_3),
    .io_salloc_req_0_bits_vc_sel_0_0(ingress_unit_0_from_1_io_salloc_req_0_bits_vc_sel_0_0),
    .io_salloc_req_0_bits_vc_sel_0_1(ingress_unit_0_from_1_io_salloc_req_0_bits_vc_sel_0_1),
    .io_salloc_req_0_bits_vc_sel_0_2(ingress_unit_0_from_1_io_salloc_req_0_bits_vc_sel_0_2),
    .io_salloc_req_0_bits_vc_sel_0_3(ingress_unit_0_from_1_io_salloc_req_0_bits_vc_sel_0_3),
    .io_salloc_req_0_bits_tail(ingress_unit_0_from_1_io_salloc_req_0_bits_tail),
    .io_out_0_valid(ingress_unit_0_from_1_io_out_0_valid),
    .io_out_0_bits_flit_head(ingress_unit_0_from_1_io_out_0_bits_flit_head),
    .io_out_0_bits_flit_tail(ingress_unit_0_from_1_io_out_0_bits_flit_tail),
    .io_out_0_bits_flit_payload(ingress_unit_0_from_1_io_out_0_bits_flit_payload),
    .io_out_0_bits_flit_flow_ingress_node(ingress_unit_0_from_1_io_out_0_bits_flit_flow_ingress_node),
    .io_out_0_bits_flit_flow_egress_node(ingress_unit_0_from_1_io_out_0_bits_flit_flow_egress_node),
    .io_out_0_bits_out_virt_channel(ingress_unit_0_from_1_io_out_0_bits_out_virt_channel),
    .io_in_ready(ingress_unit_0_from_1_io_in_ready),
    .io_in_valid(ingress_unit_0_from_1_io_in_valid),
    .io_in_bits_head(ingress_unit_0_from_1_io_in_bits_head),
    .io_in_bits_tail(ingress_unit_0_from_1_io_in_bits_tail),
    .io_in_bits_payload(ingress_unit_0_from_1_io_in_bits_payload),
    .io_in_bits_egress_id(ingress_unit_0_from_1_io_in_bits_egress_id)
  );
  OutputUnit output_unit_0_to_1 ( // @[Router.scala 122:13]
    .clock(output_unit_0_to_1_clock),
    .reset(output_unit_0_to_1_reset),
    .io_in_0_valid(output_unit_0_to_1_io_in_0_valid),
    .io_in_0_bits_head(output_unit_0_to_1_io_in_0_bits_head),
    .io_in_0_bits_tail(output_unit_0_to_1_io_in_0_bits_tail),
    .io_in_0_bits_payload(output_unit_0_to_1_io_in_0_bits_payload),
    .io_in_0_bits_flow_ingress_node(output_unit_0_to_1_io_in_0_bits_flow_ingress_node),
    .io_in_0_bits_flow_egress_node(output_unit_0_to_1_io_in_0_bits_flow_egress_node),
    .io_in_0_bits_virt_channel_id(output_unit_0_to_1_io_in_0_bits_virt_channel_id),
    .io_credit_available_1(output_unit_0_to_1_io_credit_available_1),
    .io_credit_available_2(output_unit_0_to_1_io_credit_available_2),
    .io_credit_available_3(output_unit_0_to_1_io_credit_available_3),
    .io_channel_status_1_occupied(output_unit_0_to_1_io_channel_status_1_occupied),
    .io_channel_status_2_occupied(output_unit_0_to_1_io_channel_status_2_occupied),
    .io_channel_status_3_occupied(output_unit_0_to_1_io_channel_status_3_occupied),
    .io_allocs_1_alloc(output_unit_0_to_1_io_allocs_1_alloc),
    .io_allocs_2_alloc(output_unit_0_to_1_io_allocs_2_alloc),
    .io_allocs_3_alloc(output_unit_0_to_1_io_allocs_3_alloc),
    .io_credit_alloc_1_alloc(output_unit_0_to_1_io_credit_alloc_1_alloc),
    .io_credit_alloc_2_alloc(output_unit_0_to_1_io_credit_alloc_2_alloc),
    .io_credit_alloc_3_alloc(output_unit_0_to_1_io_credit_alloc_3_alloc),
    .io_out_flit_0_valid(output_unit_0_to_1_io_out_flit_0_valid),
    .io_out_flit_0_bits_head(output_unit_0_to_1_io_out_flit_0_bits_head),
    .io_out_flit_0_bits_tail(output_unit_0_to_1_io_out_flit_0_bits_tail),
    .io_out_flit_0_bits_payload(output_unit_0_to_1_io_out_flit_0_bits_payload),
    .io_out_flit_0_bits_flow_ingress_node(output_unit_0_to_1_io_out_flit_0_bits_flow_ingress_node),
    .io_out_flit_0_bits_flow_egress_node(output_unit_0_to_1_io_out_flit_0_bits_flow_egress_node),
    .io_out_flit_0_bits_virt_channel_id(output_unit_0_to_1_io_out_flit_0_bits_virt_channel_id),
    .io_out_credit_return(output_unit_0_to_1_io_out_credit_return),
    .io_out_vc_free(output_unit_0_to_1_io_out_vc_free)
  );
  OutputUnit output_unit_1_to_3 ( // @[Router.scala 122:13]
    .clock(output_unit_1_to_3_clock),
    .reset(output_unit_1_to_3_reset),
    .io_in_0_valid(output_unit_1_to_3_io_in_0_valid),
    .io_in_0_bits_head(output_unit_1_to_3_io_in_0_bits_head),
    .io_in_0_bits_tail(output_unit_1_to_3_io_in_0_bits_tail),
    .io_in_0_bits_payload(output_unit_1_to_3_io_in_0_bits_payload),
    .io_in_0_bits_flow_ingress_node(output_unit_1_to_3_io_in_0_bits_flow_ingress_node),
    .io_in_0_bits_flow_egress_node(output_unit_1_to_3_io_in_0_bits_flow_egress_node),
    .io_in_0_bits_virt_channel_id(output_unit_1_to_3_io_in_0_bits_virt_channel_id),
    .io_credit_available_1(output_unit_1_to_3_io_credit_available_1),
    .io_credit_available_2(output_unit_1_to_3_io_credit_available_2),
    .io_credit_available_3(output_unit_1_to_3_io_credit_available_3),
    .io_channel_status_1_occupied(output_unit_1_to_3_io_channel_status_1_occupied),
    .io_channel_status_2_occupied(output_unit_1_to_3_io_channel_status_2_occupied),
    .io_channel_status_3_occupied(output_unit_1_to_3_io_channel_status_3_occupied),
    .io_allocs_1_alloc(output_unit_1_to_3_io_allocs_1_alloc),
    .io_allocs_2_alloc(output_unit_1_to_3_io_allocs_2_alloc),
    .io_allocs_3_alloc(output_unit_1_to_3_io_allocs_3_alloc),
    .io_credit_alloc_1_alloc(output_unit_1_to_3_io_credit_alloc_1_alloc),
    .io_credit_alloc_2_alloc(output_unit_1_to_3_io_credit_alloc_2_alloc),
    .io_credit_alloc_3_alloc(output_unit_1_to_3_io_credit_alloc_3_alloc),
    .io_out_flit_0_valid(output_unit_1_to_3_io_out_flit_0_valid),
    .io_out_flit_0_bits_head(output_unit_1_to_3_io_out_flit_0_bits_head),
    .io_out_flit_0_bits_tail(output_unit_1_to_3_io_out_flit_0_bits_tail),
    .io_out_flit_0_bits_payload(output_unit_1_to_3_io_out_flit_0_bits_payload),
    .io_out_flit_0_bits_flow_ingress_node(output_unit_1_to_3_io_out_flit_0_bits_flow_ingress_node),
    .io_out_flit_0_bits_flow_egress_node(output_unit_1_to_3_io_out_flit_0_bits_flow_egress_node),
    .io_out_flit_0_bits_virt_channel_id(output_unit_1_to_3_io_out_flit_0_bits_virt_channel_id),
    .io_out_credit_return(output_unit_1_to_3_io_out_credit_return),
    .io_out_vc_free(output_unit_1_to_3_io_out_vc_free)
  );
  Switch switch ( // @[Router.scala 129:24]
    .clock(switch_clock),
    .reset(switch_reset),
    .io_in_0_0_valid(switch_io_in_0_0_valid),
    .io_in_0_0_bits_flit_head(switch_io_in_0_0_bits_flit_head),
    .io_in_0_0_bits_flit_tail(switch_io_in_0_0_bits_flit_tail),
    .io_in_0_0_bits_flit_payload(switch_io_in_0_0_bits_flit_payload),
    .io_in_0_0_bits_flit_flow_ingress_node(switch_io_in_0_0_bits_flit_flow_ingress_node),
    .io_in_0_0_bits_flit_flow_egress_node(switch_io_in_0_0_bits_flit_flow_egress_node),
    .io_in_0_0_bits_out_virt_channel(switch_io_in_0_0_bits_out_virt_channel),
    .io_out_1_0_valid(switch_io_out_1_0_valid),
    .io_out_1_0_bits_head(switch_io_out_1_0_bits_head),
    .io_out_1_0_bits_tail(switch_io_out_1_0_bits_tail),
    .io_out_1_0_bits_payload(switch_io_out_1_0_bits_payload),
    .io_out_1_0_bits_flow_ingress_node(switch_io_out_1_0_bits_flow_ingress_node),
    .io_out_1_0_bits_flow_egress_node(switch_io_out_1_0_bits_flow_egress_node),
    .io_out_1_0_bits_virt_channel_id(switch_io_out_1_0_bits_virt_channel_id),
    .io_out_0_0_valid(switch_io_out_0_0_valid),
    .io_out_0_0_bits_head(switch_io_out_0_0_bits_head),
    .io_out_0_0_bits_tail(switch_io_out_0_0_bits_tail),
    .io_out_0_0_bits_payload(switch_io_out_0_0_bits_payload),
    .io_out_0_0_bits_flow_ingress_node(switch_io_out_0_0_bits_flow_ingress_node),
    .io_out_0_0_bits_flow_egress_node(switch_io_out_0_0_bits_flow_egress_node),
    .io_out_0_0_bits_virt_channel_id(switch_io_out_0_0_bits_virt_channel_id),
    .io_sel_1_0_0_0(switch_io_sel_1_0_0_0),
    .io_sel_0_0_0_0(switch_io_sel_0_0_0_0)
  );
  SwitchAllocator switch_allocator ( // @[Router.scala 130:34]
    .clock(switch_allocator_clock),
    .reset(switch_allocator_reset),
    .io_req_0_0_ready(switch_allocator_io_req_0_0_ready),
    .io_req_0_0_valid(switch_allocator_io_req_0_0_valid),
    .io_req_0_0_bits_vc_sel_1_0(switch_allocator_io_req_0_0_bits_vc_sel_1_0),
    .io_req_0_0_bits_vc_sel_1_1(switch_allocator_io_req_0_0_bits_vc_sel_1_1),
    .io_req_0_0_bits_vc_sel_1_2(switch_allocator_io_req_0_0_bits_vc_sel_1_2),
    .io_req_0_0_bits_vc_sel_1_3(switch_allocator_io_req_0_0_bits_vc_sel_1_3),
    .io_req_0_0_bits_vc_sel_0_0(switch_allocator_io_req_0_0_bits_vc_sel_0_0),
    .io_req_0_0_bits_vc_sel_0_1(switch_allocator_io_req_0_0_bits_vc_sel_0_1),
    .io_req_0_0_bits_vc_sel_0_2(switch_allocator_io_req_0_0_bits_vc_sel_0_2),
    .io_req_0_0_bits_vc_sel_0_3(switch_allocator_io_req_0_0_bits_vc_sel_0_3),
    .io_req_0_0_bits_tail(switch_allocator_io_req_0_0_bits_tail),
    .io_credit_alloc_1_1_alloc(switch_allocator_io_credit_alloc_1_1_alloc),
    .io_credit_alloc_1_2_alloc(switch_allocator_io_credit_alloc_1_2_alloc),
    .io_credit_alloc_1_3_alloc(switch_allocator_io_credit_alloc_1_3_alloc),
    .io_credit_alloc_0_1_alloc(switch_allocator_io_credit_alloc_0_1_alloc),
    .io_credit_alloc_0_2_alloc(switch_allocator_io_credit_alloc_0_2_alloc),
    .io_credit_alloc_0_3_alloc(switch_allocator_io_credit_alloc_0_3_alloc),
    .io_switch_sel_1_0_0_0(switch_allocator_io_switch_sel_1_0_0_0),
    .io_switch_sel_0_0_0_0(switch_allocator_io_switch_sel_0_0_0_0)
  );
  RotatingSingleVCAllocator vc_allocator ( // @[Router.scala 131:30]
    .clock(vc_allocator_clock),
    .reset(vc_allocator_reset),
    .io_req_0_ready(vc_allocator_io_req_0_ready),
    .io_req_0_valid(vc_allocator_io_req_0_valid),
    .io_req_0_bits_vc_sel_1_0(vc_allocator_io_req_0_bits_vc_sel_1_0),
    .io_req_0_bits_vc_sel_1_1(vc_allocator_io_req_0_bits_vc_sel_1_1),
    .io_req_0_bits_vc_sel_1_2(vc_allocator_io_req_0_bits_vc_sel_1_2),
    .io_req_0_bits_vc_sel_1_3(vc_allocator_io_req_0_bits_vc_sel_1_3),
    .io_req_0_bits_vc_sel_0_0(vc_allocator_io_req_0_bits_vc_sel_0_0),
    .io_req_0_bits_vc_sel_0_1(vc_allocator_io_req_0_bits_vc_sel_0_1),
    .io_req_0_bits_vc_sel_0_2(vc_allocator_io_req_0_bits_vc_sel_0_2),
    .io_req_0_bits_vc_sel_0_3(vc_allocator_io_req_0_bits_vc_sel_0_3),
    .io_resp_0_vc_sel_1_0(vc_allocator_io_resp_0_vc_sel_1_0),
    .io_resp_0_vc_sel_1_1(vc_allocator_io_resp_0_vc_sel_1_1),
    .io_resp_0_vc_sel_1_2(vc_allocator_io_resp_0_vc_sel_1_2),
    .io_resp_0_vc_sel_1_3(vc_allocator_io_resp_0_vc_sel_1_3),
    .io_resp_0_vc_sel_0_0(vc_allocator_io_resp_0_vc_sel_0_0),
    .io_resp_0_vc_sel_0_1(vc_allocator_io_resp_0_vc_sel_0_1),
    .io_resp_0_vc_sel_0_2(vc_allocator_io_resp_0_vc_sel_0_2),
    .io_resp_0_vc_sel_0_3(vc_allocator_io_resp_0_vc_sel_0_3),
    .io_channel_status_1_1_occupied(vc_allocator_io_channel_status_1_1_occupied),
    .io_channel_status_1_2_occupied(vc_allocator_io_channel_status_1_2_occupied),
    .io_channel_status_1_3_occupied(vc_allocator_io_channel_status_1_3_occupied),
    .io_channel_status_0_1_occupied(vc_allocator_io_channel_status_0_1_occupied),
    .io_channel_status_0_2_occupied(vc_allocator_io_channel_status_0_2_occupied),
    .io_channel_status_0_3_occupied(vc_allocator_io_channel_status_0_3_occupied),
    .io_out_allocs_1_1_alloc(vc_allocator_io_out_allocs_1_1_alloc),
    .io_out_allocs_1_2_alloc(vc_allocator_io_out_allocs_1_2_alloc),
    .io_out_allocs_1_3_alloc(vc_allocator_io_out_allocs_1_3_alloc),
    .io_out_allocs_0_1_alloc(vc_allocator_io_out_allocs_0_1_alloc),
    .io_out_allocs_0_2_alloc(vc_allocator_io_out_allocs_0_2_alloc),
    .io_out_allocs_0_3_alloc(vc_allocator_io_out_allocs_0_3_alloc)
  );
  RouteComputer_2 route_computer ( // @[Router.scala 134:32]
    .io_req_0_bits_flow_ingress_node(route_computer_io_req_0_bits_flow_ingress_node),
    .io_req_0_bits_flow_egress_node(route_computer_io_req_0_bits_flow_egress_node),
    .io_resp_0_vc_sel_1_0(route_computer_io_resp_0_vc_sel_1_0),
    .io_resp_0_vc_sel_1_1(route_computer_io_resp_0_vc_sel_1_1),
    .io_resp_0_vc_sel_1_2(route_computer_io_resp_0_vc_sel_1_2),
    .io_resp_0_vc_sel_1_3(route_computer_io_resp_0_vc_sel_1_3),
    .io_resp_0_vc_sel_0_0(route_computer_io_resp_0_vc_sel_0_0),
    .io_resp_0_vc_sel_0_1(route_computer_io_resp_0_vc_sel_0_1),
    .io_resp_0_vc_sel_0_2(route_computer_io_resp_0_vc_sel_0_2),
    .io_resp_0_vc_sel_0_3(route_computer_io_resp_0_vc_sel_0_3)
  );
  plusarg_reader #(.FORMAT("noc_util_sample_rate=%d"), .DEFAULT(0), .WIDTH(20)) plusarg_reader ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_out)
  );
  assign auto_ingress_nodes_in_flit_ready = ingress_unit_0_from_1_io_in_ready; // @[Nodes.scala 1215:84 Router.scala 142:68]
  assign auto_source_nodes_out_1_flit_0_valid = output_unit_1_to_3_io_out_flit_0_valid; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_1_flit_0_bits_head = output_unit_1_to_3_io_out_flit_0_bits_head; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_1_flit_0_bits_tail = output_unit_1_to_3_io_out_flit_0_bits_tail; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_1_flit_0_bits_payload = output_unit_1_to_3_io_out_flit_0_bits_payload; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_1_flit_0_bits_flow_ingress_node = output_unit_1_to_3_io_out_flit_0_bits_flow_ingress_node
    ; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_1_flit_0_bits_flow_egress_node = output_unit_1_to_3_io_out_flit_0_bits_flow_egress_node; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_1_flit_0_bits_virt_channel_id = output_unit_1_to_3_io_out_flit_0_bits_virt_channel_id; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_0_flit_0_valid = output_unit_0_to_1_io_out_flit_0_valid; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_0_flit_0_bits_head = output_unit_0_to_1_io_out_flit_0_bits_head; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_0_flit_0_bits_tail = output_unit_0_to_1_io_out_flit_0_bits_tail; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_0_flit_0_bits_payload = output_unit_0_to_1_io_out_flit_0_bits_payload; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_0_flit_0_bits_flow_ingress_node = output_unit_0_to_1_io_out_flit_0_bits_flow_ingress_node
    ; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_0_flit_0_bits_flow_egress_node = output_unit_0_to_1_io_out_flit_0_bits_flow_egress_node; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign auto_source_nodes_out_0_flit_0_bits_virt_channel_id = output_unit_0_to_1_io_out_flit_0_bits_virt_channel_id; // @[Nodes.scala 1212:84 Router.scala 143:60]
  assign ingress_unit_0_from_1_clock = clock;
  assign ingress_unit_0_from_1_reset = reset;
  assign ingress_unit_0_from_1_io_router_resp_vc_sel_1_0 = route_computer_io_resp_0_vc_sel_1_0; // @[Router.scala 148:38]
  assign ingress_unit_0_from_1_io_router_resp_vc_sel_1_1 = route_computer_io_resp_0_vc_sel_1_1; // @[Router.scala 148:38]
  assign ingress_unit_0_from_1_io_router_resp_vc_sel_1_2 = route_computer_io_resp_0_vc_sel_1_2; // @[Router.scala 148:38]
  assign ingress_unit_0_from_1_io_router_resp_vc_sel_1_3 = route_computer_io_resp_0_vc_sel_1_3; // @[Router.scala 148:38]
  assign ingress_unit_0_from_1_io_router_resp_vc_sel_0_0 = route_computer_io_resp_0_vc_sel_0_0; // @[Router.scala 148:38]
  assign ingress_unit_0_from_1_io_router_resp_vc_sel_0_1 = route_computer_io_resp_0_vc_sel_0_1; // @[Router.scala 148:38]
  assign ingress_unit_0_from_1_io_router_resp_vc_sel_0_2 = route_computer_io_resp_0_vc_sel_0_2; // @[Router.scala 148:38]
  assign ingress_unit_0_from_1_io_router_resp_vc_sel_0_3 = route_computer_io_resp_0_vc_sel_0_3; // @[Router.scala 148:38]
  assign ingress_unit_0_from_1_io_vcalloc_req_ready = vc_allocator_io_req_0_ready; // @[Router.scala 151:23]
  assign ingress_unit_0_from_1_io_vcalloc_resp_vc_sel_1_0 = vc_allocator_io_resp_0_vc_sel_1_0; // @[Router.scala 153:39]
  assign ingress_unit_0_from_1_io_vcalloc_resp_vc_sel_1_1 = vc_allocator_io_resp_0_vc_sel_1_1; // @[Router.scala 153:39]
  assign ingress_unit_0_from_1_io_vcalloc_resp_vc_sel_1_2 = vc_allocator_io_resp_0_vc_sel_1_2; // @[Router.scala 153:39]
  assign ingress_unit_0_from_1_io_vcalloc_resp_vc_sel_1_3 = vc_allocator_io_resp_0_vc_sel_1_3; // @[Router.scala 153:39]
  assign ingress_unit_0_from_1_io_vcalloc_resp_vc_sel_0_0 = vc_allocator_io_resp_0_vc_sel_0_0; // @[Router.scala 153:39]
  assign ingress_unit_0_from_1_io_vcalloc_resp_vc_sel_0_1 = vc_allocator_io_resp_0_vc_sel_0_1; // @[Router.scala 153:39]
  assign ingress_unit_0_from_1_io_vcalloc_resp_vc_sel_0_2 = vc_allocator_io_resp_0_vc_sel_0_2; // @[Router.scala 153:39]
  assign ingress_unit_0_from_1_io_vcalloc_resp_vc_sel_0_3 = vc_allocator_io_resp_0_vc_sel_0_3; // @[Router.scala 153:39]
  assign ingress_unit_0_from_1_io_out_credit_available_1_1 = output_unit_1_to_3_io_credit_available_1; // @[Router.scala 162:42]
  assign ingress_unit_0_from_1_io_out_credit_available_1_2 = output_unit_1_to_3_io_credit_available_2; // @[Router.scala 162:42]
  assign ingress_unit_0_from_1_io_out_credit_available_1_3 = output_unit_1_to_3_io_credit_available_3; // @[Router.scala 162:42]
  assign ingress_unit_0_from_1_io_out_credit_available_0_1 = output_unit_0_to_1_io_credit_available_1; // @[Router.scala 162:42]
  assign ingress_unit_0_from_1_io_out_credit_available_0_2 = output_unit_0_to_1_io_credit_available_2; // @[Router.scala 162:42]
  assign ingress_unit_0_from_1_io_out_credit_available_0_3 = output_unit_0_to_1_io_credit_available_3; // @[Router.scala 162:42]
  assign ingress_unit_0_from_1_io_salloc_req_0_ready = switch_allocator_io_req_0_0_ready; // @[Router.scala 165:23]
  assign ingress_unit_0_from_1_io_in_valid = auto_ingress_nodes_in_flit_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign ingress_unit_0_from_1_io_in_bits_head = auto_ingress_nodes_in_flit_bits_head; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign ingress_unit_0_from_1_io_in_bits_tail = auto_ingress_nodes_in_flit_bits_tail; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign ingress_unit_0_from_1_io_in_bits_payload = auto_ingress_nodes_in_flit_bits_payload; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign ingress_unit_0_from_1_io_in_bits_egress_id = auto_ingress_nodes_in_flit_bits_egress_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign output_unit_0_to_1_clock = clock;
  assign output_unit_0_to_1_reset = reset;
  assign output_unit_0_to_1_io_in_0_valid = switch_io_out_0_0_valid; // @[Router.scala 172:29]
  assign output_unit_0_to_1_io_in_0_bits_head = switch_io_out_0_0_bits_head; // @[Router.scala 172:29]
  assign output_unit_0_to_1_io_in_0_bits_tail = switch_io_out_0_0_bits_tail; // @[Router.scala 172:29]
  assign output_unit_0_to_1_io_in_0_bits_payload = switch_io_out_0_0_bits_payload; // @[Router.scala 172:29]
  assign output_unit_0_to_1_io_in_0_bits_flow_ingress_node = switch_io_out_0_0_bits_flow_ingress_node; // @[Router.scala 172:29]
  assign output_unit_0_to_1_io_in_0_bits_flow_egress_node = switch_io_out_0_0_bits_flow_egress_node; // @[Router.scala 172:29]
  assign output_unit_0_to_1_io_in_0_bits_virt_channel_id = switch_io_out_0_0_bits_virt_channel_id; // @[Router.scala 172:29]
  assign output_unit_0_to_1_io_allocs_1_alloc = vc_allocator_io_out_allocs_0_1_alloc; // @[Router.scala 157:33]
  assign output_unit_0_to_1_io_allocs_2_alloc = vc_allocator_io_out_allocs_0_2_alloc; // @[Router.scala 157:33]
  assign output_unit_0_to_1_io_allocs_3_alloc = vc_allocator_io_out_allocs_0_3_alloc; // @[Router.scala 157:33]
  assign output_unit_0_to_1_io_credit_alloc_1_alloc = switch_allocator_io_credit_alloc_0_1_alloc; // @[Router.scala 167:39]
  assign output_unit_0_to_1_io_credit_alloc_2_alloc = switch_allocator_io_credit_alloc_0_2_alloc; // @[Router.scala 167:39]
  assign output_unit_0_to_1_io_credit_alloc_3_alloc = switch_allocator_io_credit_alloc_0_3_alloc; // @[Router.scala 167:39]
  assign output_unit_0_to_1_io_out_credit_return = auto_source_nodes_out_0_credit_return; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign output_unit_0_to_1_io_out_vc_free = auto_source_nodes_out_0_vc_free; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign output_unit_1_to_3_clock = clock;
  assign output_unit_1_to_3_reset = reset;
  assign output_unit_1_to_3_io_in_0_valid = switch_io_out_1_0_valid; // @[Router.scala 172:29]
  assign output_unit_1_to_3_io_in_0_bits_head = switch_io_out_1_0_bits_head; // @[Router.scala 172:29]
  assign output_unit_1_to_3_io_in_0_bits_tail = switch_io_out_1_0_bits_tail; // @[Router.scala 172:29]
  assign output_unit_1_to_3_io_in_0_bits_payload = switch_io_out_1_0_bits_payload; // @[Router.scala 172:29]
  assign output_unit_1_to_3_io_in_0_bits_flow_ingress_node = switch_io_out_1_0_bits_flow_ingress_node; // @[Router.scala 172:29]
  assign output_unit_1_to_3_io_in_0_bits_flow_egress_node = switch_io_out_1_0_bits_flow_egress_node; // @[Router.scala 172:29]
  assign output_unit_1_to_3_io_in_0_bits_virt_channel_id = switch_io_out_1_0_bits_virt_channel_id; // @[Router.scala 172:29]
  assign output_unit_1_to_3_io_allocs_1_alloc = vc_allocator_io_out_allocs_1_1_alloc; // @[Router.scala 157:33]
  assign output_unit_1_to_3_io_allocs_2_alloc = vc_allocator_io_out_allocs_1_2_alloc; // @[Router.scala 157:33]
  assign output_unit_1_to_3_io_allocs_3_alloc = vc_allocator_io_out_allocs_1_3_alloc; // @[Router.scala 157:33]
  assign output_unit_1_to_3_io_credit_alloc_1_alloc = switch_allocator_io_credit_alloc_1_1_alloc; // @[Router.scala 167:39]
  assign output_unit_1_to_3_io_credit_alloc_2_alloc = switch_allocator_io_credit_alloc_1_2_alloc; // @[Router.scala 167:39]
  assign output_unit_1_to_3_io_credit_alloc_3_alloc = switch_allocator_io_credit_alloc_1_3_alloc; // @[Router.scala 167:39]
  assign output_unit_1_to_3_io_out_credit_return = auto_source_nodes_out_1_credit_return; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign output_unit_1_to_3_io_out_vc_free = auto_source_nodes_out_1_vc_free; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign switch_clock = clock;
  assign switch_reset = reset;
  assign switch_io_in_0_0_valid = ingress_unit_0_from_1_io_out_0_valid; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_head = ingress_unit_0_from_1_io_out_0_bits_flit_head; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_tail = ingress_unit_0_from_1_io_out_0_bits_flit_tail; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_payload = ingress_unit_0_from_1_io_out_0_bits_flit_payload; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_flow_ingress_node = ingress_unit_0_from_1_io_out_0_bits_flit_flow_ingress_node; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_flow_egress_node = ingress_unit_0_from_1_io_out_0_bits_flit_flow_egress_node; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_out_virt_channel = ingress_unit_0_from_1_io_out_0_bits_out_virt_channel; // @[Router.scala 170:23]
  assign switch_io_sel_1_0_0_0 = switch_io_sel_REG_1_0_0_0; // @[Router.scala 173:19]
  assign switch_io_sel_0_0_0_0 = switch_io_sel_REG_0_0_0_0; // @[Router.scala 173:19]
  assign switch_allocator_clock = clock;
  assign switch_allocator_reset = reset;
  assign switch_allocator_io_req_0_0_valid = ingress_unit_0_from_1_io_salloc_req_0_valid; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_1_0 = ingress_unit_0_from_1_io_salloc_req_0_bits_vc_sel_1_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_1_1 = ingress_unit_0_from_1_io_salloc_req_0_bits_vc_sel_1_1; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_1_2 = ingress_unit_0_from_1_io_salloc_req_0_bits_vc_sel_1_2; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_1_3 = ingress_unit_0_from_1_io_salloc_req_0_bits_vc_sel_1_3; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_0_0 = ingress_unit_0_from_1_io_salloc_req_0_bits_vc_sel_0_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_0_1 = ingress_unit_0_from_1_io_salloc_req_0_bits_vc_sel_0_1; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_0_2 = ingress_unit_0_from_1_io_salloc_req_0_bits_vc_sel_0_2; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_0_3 = ingress_unit_0_from_1_io_salloc_req_0_bits_vc_sel_0_3; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_tail = ingress_unit_0_from_1_io_salloc_req_0_bits_tail; // @[Router.scala 165:23]
  assign vc_allocator_clock = clock;
  assign vc_allocator_reset = reset;
  assign vc_allocator_io_req_0_valid = ingress_unit_0_from_1_io_vcalloc_req_valid; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_1_0 = ingress_unit_0_from_1_io_vcalloc_req_bits_vc_sel_1_0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_1_1 = ingress_unit_0_from_1_io_vcalloc_req_bits_vc_sel_1_1; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_1_2 = ingress_unit_0_from_1_io_vcalloc_req_bits_vc_sel_1_2; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_1_3 = ingress_unit_0_from_1_io_vcalloc_req_bits_vc_sel_1_3; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_0_0 = ingress_unit_0_from_1_io_vcalloc_req_bits_vc_sel_0_0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_0_1 = ingress_unit_0_from_1_io_vcalloc_req_bits_vc_sel_0_1; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_0_2 = ingress_unit_0_from_1_io_vcalloc_req_bits_vc_sel_0_2; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_0_3 = ingress_unit_0_from_1_io_vcalloc_req_bits_vc_sel_0_3; // @[Router.scala 151:23]
  assign vc_allocator_io_channel_status_1_1_occupied = output_unit_1_to_3_io_channel_status_1_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_1_2_occupied = output_unit_1_to_3_io_channel_status_2_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_1_3_occupied = output_unit_1_to_3_io_channel_status_3_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_0_1_occupied = output_unit_0_to_1_io_channel_status_1_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_0_2_occupied = output_unit_0_to_1_io_channel_status_2_occupied; // @[Router.scala 159:23]
  assign vc_allocator_io_channel_status_0_3_occupied = output_unit_0_to_1_io_channel_status_3_occupied; // @[Router.scala 159:23]
  assign route_computer_io_req_0_bits_flow_ingress_node = ingress_unit_0_from_1_io_router_req_bits_flow_ingress_node; // @[Router.scala 146:23]
  assign route_computer_io_req_0_bits_flow_egress_node = ingress_unit_0_from_1_io_router_req_bits_flow_egress_node; // @[Router.scala 146:23]
  always @(posedge clock) begin
    switch_io_sel_REG_1_0_0_0 <= switch_allocator_io_switch_sel_1_0_0_0; // @[Router.scala 176:14]
    switch_io_sel_REG_0_0_0_0 <= switch_allocator_io_switch_sel_0_0_0_0; // @[Router.scala 176:14]
    if (reset) begin // @[Router.scala 193:28]
      debug_tsc <= 64'h0; // @[Router.scala 193:28]
    end else begin
      debug_tsc <= _debug_tsc_T_1; // @[Router.scala 194:15]
    end
    if (reset) begin // @[Router.scala 195:31]
      debug_sample <= 64'h0; // @[Router.scala 195:31]
    end else if (debug_sample == _GEN_2) begin // @[Router.scala 198:47]
      debug_sample <= 64'h0; // @[Router.scala 198:62]
    end else begin
      debug_sample <= _debug_sample_T_1; // @[Router.scala 196:18]
    end
    if (reset) begin // @[Router.scala 201:29]
      util_ctr <= 64'h0; // @[Router.scala 201:29]
    end else begin
      util_ctr <= _util_ctr_T_1; // @[Router.scala 203:16]
    end
    if (reset) begin // @[Router.scala 202:26]
      fired <= 1'h0; // @[Router.scala 202:26]
    end else if (plusarg_reader_out != 20'h0 & _T_2 & fired) begin // @[Router.scala 205:81]
      fired <= _T_3; // @[Router.scala 208:15]
    end else begin
      fired <= fired | _T_3; // @[Router.scala 204:13]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9 & ~reset) begin
          $fwrite(32'h80000002,"nocsample %d i1 2 %d\n",debug_tsc,util_ctr); // @[Router.scala 207:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  switch_io_sel_REG_1_0_0_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  switch_io_sel_REG_0_0_0_0 = _RAND_1[0:0];
  _RAND_2 = {2{`RANDOM}};
  debug_tsc = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  debug_sample = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  util_ctr = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  fired = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ClockSinkDomain_2(
  output        auto_routers_ingress_nodes_in_flit_ready,
  input         auto_routers_ingress_nodes_in_flit_valid,
  input         auto_routers_ingress_nodes_in_flit_bits_head,
  input         auto_routers_ingress_nodes_in_flit_bits_tail,
  input  [63:0] auto_routers_ingress_nodes_in_flit_bits_payload,
  input         auto_routers_ingress_nodes_in_flit_bits_egress_id,
  output        auto_routers_source_nodes_out_1_flit_0_valid,
  output        auto_routers_source_nodes_out_1_flit_0_bits_head,
  output        auto_routers_source_nodes_out_1_flit_0_bits_tail,
  output [63:0] auto_routers_source_nodes_out_1_flit_0_bits_payload,
  output [1:0]  auto_routers_source_nodes_out_1_flit_0_bits_flow_ingress_node,
  output [1:0]  auto_routers_source_nodes_out_1_flit_0_bits_flow_egress_node,
  output [1:0]  auto_routers_source_nodes_out_1_flit_0_bits_virt_channel_id,
  input  [3:0]  auto_routers_source_nodes_out_1_credit_return,
  input  [3:0]  auto_routers_source_nodes_out_1_vc_free,
  output        auto_routers_source_nodes_out_0_flit_0_valid,
  output        auto_routers_source_nodes_out_0_flit_0_bits_head,
  output        auto_routers_source_nodes_out_0_flit_0_bits_tail,
  output [63:0] auto_routers_source_nodes_out_0_flit_0_bits_payload,
  output [1:0]  auto_routers_source_nodes_out_0_flit_0_bits_flow_ingress_node,
  output [1:0]  auto_routers_source_nodes_out_0_flit_0_bits_flow_egress_node,
  output [1:0]  auto_routers_source_nodes_out_0_flit_0_bits_virt_channel_id,
  input  [3:0]  auto_routers_source_nodes_out_0_credit_return,
  input  [3:0]  auto_routers_source_nodes_out_0_vc_free,
  input         auto_clock_in_clock,
  input         auto_clock_in_reset
);
  wire  routers_clock; // @[NoC.scala 64:22]
  wire  routers_reset; // @[NoC.scala 64:22]
  wire  routers_auto_ingress_nodes_in_flit_ready; // @[NoC.scala 64:22]
  wire  routers_auto_ingress_nodes_in_flit_valid; // @[NoC.scala 64:22]
  wire  routers_auto_ingress_nodes_in_flit_bits_head; // @[NoC.scala 64:22]
  wire  routers_auto_ingress_nodes_in_flit_bits_tail; // @[NoC.scala 64:22]
  wire [63:0] routers_auto_ingress_nodes_in_flit_bits_payload; // @[NoC.scala 64:22]
  wire  routers_auto_ingress_nodes_in_flit_bits_egress_id; // @[NoC.scala 64:22]
  wire  routers_auto_source_nodes_out_1_flit_0_valid; // @[NoC.scala 64:22]
  wire  routers_auto_source_nodes_out_1_flit_0_bits_head; // @[NoC.scala 64:22]
  wire  routers_auto_source_nodes_out_1_flit_0_bits_tail; // @[NoC.scala 64:22]
  wire [63:0] routers_auto_source_nodes_out_1_flit_0_bits_payload; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_source_nodes_out_1_flit_0_bits_flow_ingress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_source_nodes_out_1_flit_0_bits_flow_egress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_source_nodes_out_1_flit_0_bits_virt_channel_id; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_source_nodes_out_1_credit_return; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_source_nodes_out_1_vc_free; // @[NoC.scala 64:22]
  wire  routers_auto_source_nodes_out_0_flit_0_valid; // @[NoC.scala 64:22]
  wire  routers_auto_source_nodes_out_0_flit_0_bits_head; // @[NoC.scala 64:22]
  wire  routers_auto_source_nodes_out_0_flit_0_bits_tail; // @[NoC.scala 64:22]
  wire [63:0] routers_auto_source_nodes_out_0_flit_0_bits_payload; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_source_nodes_out_0_flit_0_bits_flow_ingress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_source_nodes_out_0_flit_0_bits_flow_egress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_source_nodes_out_0_flit_0_bits_virt_channel_id; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_source_nodes_out_0_credit_return; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_source_nodes_out_0_vc_free; // @[NoC.scala 64:22]
  Router_2 routers ( // @[NoC.scala 64:22]
    .clock(routers_clock),
    .reset(routers_reset),
    .auto_ingress_nodes_in_flit_ready(routers_auto_ingress_nodes_in_flit_ready),
    .auto_ingress_nodes_in_flit_valid(routers_auto_ingress_nodes_in_flit_valid),
    .auto_ingress_nodes_in_flit_bits_head(routers_auto_ingress_nodes_in_flit_bits_head),
    .auto_ingress_nodes_in_flit_bits_tail(routers_auto_ingress_nodes_in_flit_bits_tail),
    .auto_ingress_nodes_in_flit_bits_payload(routers_auto_ingress_nodes_in_flit_bits_payload),
    .auto_ingress_nodes_in_flit_bits_egress_id(routers_auto_ingress_nodes_in_flit_bits_egress_id),
    .auto_source_nodes_out_1_flit_0_valid(routers_auto_source_nodes_out_1_flit_0_valid),
    .auto_source_nodes_out_1_flit_0_bits_head(routers_auto_source_nodes_out_1_flit_0_bits_head),
    .auto_source_nodes_out_1_flit_0_bits_tail(routers_auto_source_nodes_out_1_flit_0_bits_tail),
    .auto_source_nodes_out_1_flit_0_bits_payload(routers_auto_source_nodes_out_1_flit_0_bits_payload),
    .auto_source_nodes_out_1_flit_0_bits_flow_ingress_node(routers_auto_source_nodes_out_1_flit_0_bits_flow_ingress_node
      ),
    .auto_source_nodes_out_1_flit_0_bits_flow_egress_node(routers_auto_source_nodes_out_1_flit_0_bits_flow_egress_node),
    .auto_source_nodes_out_1_flit_0_bits_virt_channel_id(routers_auto_source_nodes_out_1_flit_0_bits_virt_channel_id),
    .auto_source_nodes_out_1_credit_return(routers_auto_source_nodes_out_1_credit_return),
    .auto_source_nodes_out_1_vc_free(routers_auto_source_nodes_out_1_vc_free),
    .auto_source_nodes_out_0_flit_0_valid(routers_auto_source_nodes_out_0_flit_0_valid),
    .auto_source_nodes_out_0_flit_0_bits_head(routers_auto_source_nodes_out_0_flit_0_bits_head),
    .auto_source_nodes_out_0_flit_0_bits_tail(routers_auto_source_nodes_out_0_flit_0_bits_tail),
    .auto_source_nodes_out_0_flit_0_bits_payload(routers_auto_source_nodes_out_0_flit_0_bits_payload),
    .auto_source_nodes_out_0_flit_0_bits_flow_ingress_node(routers_auto_source_nodes_out_0_flit_0_bits_flow_ingress_node
      ),
    .auto_source_nodes_out_0_flit_0_bits_flow_egress_node(routers_auto_source_nodes_out_0_flit_0_bits_flow_egress_node),
    .auto_source_nodes_out_0_flit_0_bits_virt_channel_id(routers_auto_source_nodes_out_0_flit_0_bits_virt_channel_id),
    .auto_source_nodes_out_0_credit_return(routers_auto_source_nodes_out_0_credit_return),
    .auto_source_nodes_out_0_vc_free(routers_auto_source_nodes_out_0_vc_free)
  );
  assign auto_routers_ingress_nodes_in_flit_ready = routers_auto_ingress_nodes_in_flit_ready; // @[LazyModule.scala 366:16]
  assign auto_routers_source_nodes_out_1_flit_0_valid = routers_auto_source_nodes_out_1_flit_0_valid; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_1_flit_0_bits_head = routers_auto_source_nodes_out_1_flit_0_bits_head; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_1_flit_0_bits_tail = routers_auto_source_nodes_out_1_flit_0_bits_tail; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_1_flit_0_bits_payload = routers_auto_source_nodes_out_1_flit_0_bits_payload; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_1_flit_0_bits_flow_ingress_node =
    routers_auto_source_nodes_out_1_flit_0_bits_flow_ingress_node; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_1_flit_0_bits_flow_egress_node =
    routers_auto_source_nodes_out_1_flit_0_bits_flow_egress_node; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_1_flit_0_bits_virt_channel_id =
    routers_auto_source_nodes_out_1_flit_0_bits_virt_channel_id; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_0_flit_0_valid = routers_auto_source_nodes_out_0_flit_0_valid; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_0_flit_0_bits_head = routers_auto_source_nodes_out_0_flit_0_bits_head; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_0_flit_0_bits_tail = routers_auto_source_nodes_out_0_flit_0_bits_tail; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_0_flit_0_bits_payload = routers_auto_source_nodes_out_0_flit_0_bits_payload; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_0_flit_0_bits_flow_ingress_node =
    routers_auto_source_nodes_out_0_flit_0_bits_flow_ingress_node; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_0_flit_0_bits_flow_egress_node =
    routers_auto_source_nodes_out_0_flit_0_bits_flow_egress_node; // @[LazyModule.scala 368:12]
  assign auto_routers_source_nodes_out_0_flit_0_bits_virt_channel_id =
    routers_auto_source_nodes_out_0_flit_0_bits_virt_channel_id; // @[LazyModule.scala 368:12]
  assign routers_clock = auto_clock_in_clock; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign routers_reset = auto_clock_in_reset; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign routers_auto_ingress_nodes_in_flit_valid = auto_routers_ingress_nodes_in_flit_valid; // @[LazyModule.scala 366:16]
  assign routers_auto_ingress_nodes_in_flit_bits_head = auto_routers_ingress_nodes_in_flit_bits_head; // @[LazyModule.scala 366:16]
  assign routers_auto_ingress_nodes_in_flit_bits_tail = auto_routers_ingress_nodes_in_flit_bits_tail; // @[LazyModule.scala 366:16]
  assign routers_auto_ingress_nodes_in_flit_bits_payload = auto_routers_ingress_nodes_in_flit_bits_payload; // @[LazyModule.scala 366:16]
  assign routers_auto_ingress_nodes_in_flit_bits_egress_id = auto_routers_ingress_nodes_in_flit_bits_egress_id; // @[LazyModule.scala 366:16]
  assign routers_auto_source_nodes_out_1_credit_return = auto_routers_source_nodes_out_1_credit_return; // @[LazyModule.scala 368:12]
  assign routers_auto_source_nodes_out_1_vc_free = auto_routers_source_nodes_out_1_vc_free; // @[LazyModule.scala 368:12]
  assign routers_auto_source_nodes_out_0_credit_return = auto_routers_source_nodes_out_0_credit_return; // @[LazyModule.scala 368:12]
  assign routers_auto_source_nodes_out_0_vc_free = auto_routers_source_nodes_out_0_vc_free; // @[LazyModule.scala 368:12]
endmodule
module NoCMonitor_2(
  input        clock,
  input        reset,
  input        io_in_flit_0_valid,
  input        io_in_flit_0_bits_head,
  input        io_in_flit_0_bits_tail,
  input  [1:0] io_in_flit_0_bits_flow_ingress_node,
  input  [1:0] io_in_flit_0_bits_flow_egress_node,
  input  [1:0] io_in_flit_0_bits_virt_channel_id
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg  in_flight_0; // @[Monitor.scala 16:26]
  reg  in_flight_1; // @[Monitor.scala 16:26]
  reg  in_flight_2; // @[Monitor.scala 16:26]
  reg  in_flight_3; // @[Monitor.scala 16:26]
  wire  _GEN_0 = 2'h0 == io_in_flit_0_bits_virt_channel_id | in_flight_0; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_1 = 2'h1 == io_in_flit_0_bits_virt_channel_id | in_flight_1; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_2 = 2'h2 == io_in_flit_0_bits_virt_channel_id | in_flight_2; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_3 = 2'h3 == io_in_flit_0_bits_virt_channel_id | in_flight_3; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_5 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? in_flight_1 : in_flight_0; // @[Monitor.scala 22:{17,17}]
  wire  _GEN_6 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? in_flight_2 : _GEN_5; // @[Monitor.scala 22:{17,17}]
  wire  _GEN_7 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? in_flight_3 : _GEN_6; // @[Monitor.scala 22:{17,17}]
  wire  _T_2 = ~reset; // @[Monitor.scala 22:16]
  wire  _GEN_8 = io_in_flit_0_bits_head ? _GEN_0 : in_flight_0; // @[Monitor.scala 16:26 20:29]
  wire  _GEN_9 = io_in_flit_0_bits_head ? _GEN_1 : in_flight_1; // @[Monitor.scala 16:26 20:29]
  wire  _GEN_10 = io_in_flit_0_bits_head ? _GEN_2 : in_flight_2; // @[Monitor.scala 16:26 20:29]
  wire  _GEN_11 = io_in_flit_0_bits_head ? _GEN_3 : in_flight_3; // @[Monitor.scala 16:26 20:29]
  wire  _T_4 = io_in_flit_0_valid & io_in_flit_0_bits_head; // @[Monitor.scala 29:22]
  wire  _T_12 = io_in_flit_0_bits_flow_egress_node == 2'h3; // @[Types.scala 54:21]
  wire  _T_13 = io_in_flit_0_bits_flow_ingress_node == 2'h0 & _T_12; // @[Types.scala 53:39]
  wire  _GEN_29 = _T_4 & ~reset; // @[Monitor.scala 22:16]
  always @(posedge clock) begin
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_0 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h0 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_0 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_0 <= _GEN_8;
        end
      end else begin
        in_flight_0 <= _GEN_8;
      end
    end
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_1 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h1 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_1 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_1 <= _GEN_9;
        end
      end else begin
        in_flight_1 <= _GEN_9;
      end
    end
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_2 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h2 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_2 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_2 <= _GEN_10;
        end
      end else begin
        in_flight_2 <= _GEN_10;
      end
    end
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_3 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h3 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_3 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_3 <= _GEN_11;
        end
      end else begin
        in_flight_3 <= _GEN_11;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4 & ~reset & ~(~_GEN_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed: Flit head/tail sequencing is broken\n    at Monitor.scala:22 assert (!in_flight(flit.bits.virt_channel_id), \"Flit head/tail sequencing is broken\")\n"
            ); // @[Monitor.scala 22:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h1 | _T_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h2 | _T_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h3 | _T_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  in_flight_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  in_flight_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  in_flight_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  in_flight_3 = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (_T_4 & ~reset) begin
      assert(~_GEN_7); // @[Monitor.scala 22:16]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h0); // @[Monitor.scala 32:17]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h1 | _T_13); // @[Monitor.scala 32:17]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h2 | _T_13); // @[Monitor.scala 32:17]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h3 | _T_13); // @[Monitor.scala 32:17]
    end
  end
endmodule
module NoCMonitor_3(
  input        clock,
  input        reset,
  input        io_in_flit_0_valid,
  input        io_in_flit_0_bits_head,
  input        io_in_flit_0_bits_tail,
  input  [1:0] io_in_flit_0_bits_flow_ingress_node,
  input  [1:0] io_in_flit_0_bits_flow_egress_node,
  input  [1:0] io_in_flit_0_bits_virt_channel_id
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg  in_flight_0; // @[Monitor.scala 16:26]
  reg  in_flight_1; // @[Monitor.scala 16:26]
  reg  in_flight_2; // @[Monitor.scala 16:26]
  reg  in_flight_3; // @[Monitor.scala 16:26]
  wire  _GEN_0 = 2'h0 == io_in_flit_0_bits_virt_channel_id | in_flight_0; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_1 = 2'h1 == io_in_flit_0_bits_virt_channel_id | in_flight_1; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_2 = 2'h2 == io_in_flit_0_bits_virt_channel_id | in_flight_2; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_3 = 2'h3 == io_in_flit_0_bits_virt_channel_id | in_flight_3; // @[Monitor.scala 16:26 21:{46,46}]
  wire  _GEN_5 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? in_flight_1 : in_flight_0; // @[Monitor.scala 22:{17,17}]
  wire  _GEN_6 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? in_flight_2 : _GEN_5; // @[Monitor.scala 22:{17,17}]
  wire  _GEN_7 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? in_flight_3 : _GEN_6; // @[Monitor.scala 22:{17,17}]
  wire  _T_2 = ~reset; // @[Monitor.scala 22:16]
  wire  _GEN_8 = io_in_flit_0_bits_head ? _GEN_0 : in_flight_0; // @[Monitor.scala 16:26 20:29]
  wire  _GEN_9 = io_in_flit_0_bits_head ? _GEN_1 : in_flight_1; // @[Monitor.scala 16:26 20:29]
  wire  _GEN_10 = io_in_flit_0_bits_head ? _GEN_2 : in_flight_2; // @[Monitor.scala 16:26 20:29]
  wire  _GEN_11 = io_in_flit_0_bits_head ? _GEN_3 : in_flight_3; // @[Monitor.scala 16:26 20:29]
  wire  _T_4 = io_in_flit_0_valid & io_in_flit_0_bits_head; // @[Monitor.scala 29:22]
  wire  _T_12 = io_in_flit_0_bits_flow_egress_node == 2'h3; // @[Types.scala 54:21]
  wire  _T_13 = io_in_flit_0_bits_flow_ingress_node == 2'h2 & _T_12; // @[Types.scala 53:39]
  wire  _GEN_29 = _T_4 & ~reset; // @[Monitor.scala 22:16]
  always @(posedge clock) begin
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_0 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h0 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_0 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_0 <= _GEN_8;
        end
      end else begin
        in_flight_0 <= _GEN_8;
      end
    end
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_1 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h1 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_1 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_1 <= _GEN_9;
        end
      end else begin
        in_flight_1 <= _GEN_9;
      end
    end
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_2 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h2 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_2 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_2 <= _GEN_10;
        end
      end else begin
        in_flight_2 <= _GEN_10;
      end
    end
    if (reset) begin // @[Monitor.scala 16:26]
      in_flight_3 <= 1'h0; // @[Monitor.scala 16:26]
    end else if (io_in_flit_0_valid) begin // @[Monitor.scala 19:23]
      if (io_in_flit_0_bits_tail) begin // @[Monitor.scala 24:29]
        if (2'h3 == io_in_flit_0_bits_virt_channel_id) begin // @[Monitor.scala 25:46]
          in_flight_3 <= 1'h0; // @[Monitor.scala 25:46]
        end else begin
          in_flight_3 <= _GEN_11;
        end
      end else begin
        in_flight_3 <= _GEN_11;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4 & ~reset & ~(~_GEN_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed: Flit head/tail sequencing is broken\n    at Monitor.scala:22 assert (!in_flight(flit.bits.virt_channel_id), \"Flit head/tail sequencing is broken\")\n"
            ); // @[Monitor.scala 22:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h1 | _T_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h2 | _T_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & ~(io_in_flit_0_bits_virt_channel_id != 2'h3 | _T_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Monitor.scala:32 assert(flit.bits.virt_channel_id =/= i.U || v.possibleFlows.toSeq.map(_.isFlow(flit.bits.flow)).orR)\n"
            ); // @[Monitor.scala 32:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  in_flight_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  in_flight_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  in_flight_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  in_flight_3 = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (_T_4 & ~reset) begin
      assert(~_GEN_7); // @[Monitor.scala 22:16]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h0); // @[Monitor.scala 32:17]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h1 | _T_13); // @[Monitor.scala 32:17]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h2 | _T_13); // @[Monitor.scala 32:17]
    end
    //
    if (_T_4 & _T_2) begin
      assert(io_in_flit_0_bits_virt_channel_id != 2'h3 | _T_13); // @[Monitor.scala 32:17]
    end
  end
endmodule
module InputUnit_2(
  input         clock,
  input         reset,
  output        io_router_req_valid,
  output [1:0]  io_router_req_bits_src_virt_id,
  input         io_vcalloc_req_ready,
  output        io_vcalloc_req_valid,
  output        io_vcalloc_req_bits_vc_sel_0_0,
  input         io_vcalloc_resp_vc_sel_0_0,
  input         io_out_credit_available_0_0,
  input         io_salloc_req_0_ready,
  output        io_salloc_req_0_valid,
  output        io_salloc_req_0_bits_vc_sel_0_0,
  output        io_salloc_req_0_bits_tail,
  output        io_out_0_valid,
  output        io_out_0_bits_flit_head,
  output        io_out_0_bits_flit_tail,
  output [63:0] io_out_0_bits_flit_payload,
  output [1:0]  io_out_0_bits_flit_flow_ingress_node,
  output [1:0]  io_debug_va_stall,
  output [1:0]  io_debug_sa_stall,
  input         io_in_flit_0_valid,
  input         io_in_flit_0_bits_head,
  input         io_in_flit_0_bits_tail,
  input  [63:0] io_in_flit_0_bits_payload,
  input  [1:0]  io_in_flit_0_bits_flow_ingress_node,
  input  [1:0]  io_in_flit_0_bits_flow_egress_node,
  input  [1:0]  io_in_flit_0_bits_virt_channel_id,
  output [3:0]  io_in_credit_return,
  output [3:0]  io_in_vc_free
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
`endif // RANDOMIZE_REG_INIT
  wire  input_buffer_clock; // @[InputUnit.scala 180:28]
  wire  input_buffer_reset; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_enq_0_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_enq_0_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_enq_0_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_enq_0_bits_payload; // @[InputUnit.scala 180:28]
  wire [1:0] input_buffer_io_enq_0_bits_virt_channel_id; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_0_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_0_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_deq_0_bits_payload; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_ready; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_1_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_deq_1_bits_payload; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_ready; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_2_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_deq_2_bits_payload; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_3_ready; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_3_valid; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_3_bits_head; // @[InputUnit.scala 180:28]
  wire  input_buffer_io_deq_3_bits_tail; // @[InputUnit.scala 180:28]
  wire [63:0] input_buffer_io_deq_3_bits_payload; // @[InputUnit.scala 180:28]
  wire  route_arbiter_io_in_1_valid; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_2_ready; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_2_valid; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_3_ready; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_in_3_valid; // @[InputUnit.scala 186:29]
  wire  route_arbiter_io_out_valid; // @[InputUnit.scala 186:29]
  wire [1:0] route_arbiter_io_out_bits_src_virt_id; // @[InputUnit.scala 186:29]
  wire  salloc_arb_clock; // @[InputUnit.scala 279:26]
  wire  salloc_arb_reset; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_0_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_1_bits_tail; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_2_bits_tail; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_in_3_bits_tail; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_ready; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_valid; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_vc_sel_0_0; // @[InputUnit.scala 279:26]
  wire  salloc_arb_io_out_0_bits_tail; // @[InputUnit.scala 279:26]
  wire [3:0] salloc_arb_io_chosen_oh_0; // @[InputUnit.scala 279:26]
  reg [2:0] states_1_g; // @[InputUnit.scala 191:19]
  reg  states_1_vc_sel_0_0; // @[InputUnit.scala 191:19]
  reg [1:0] states_1_flow_ingress_node; // @[InputUnit.scala 191:19]
  reg [2:0] states_2_g; // @[InputUnit.scala 191:19]
  reg  states_2_vc_sel_0_0; // @[InputUnit.scala 191:19]
  reg [1:0] states_2_flow_ingress_node; // @[InputUnit.scala 191:19]
  reg [2:0] states_3_g; // @[InputUnit.scala 191:19]
  reg  states_3_vc_sel_0_0; // @[InputUnit.scala 191:19]
  reg [1:0] states_3_flow_ingress_node; // @[InputUnit.scala 191:19]
  wire  _T = io_in_flit_0_valid & io_in_flit_0_bits_head; // @[InputUnit.scala 194:32]
  wire  _T_3 = ~reset; // @[InputUnit.scala 196:13]
  wire [2:0] _GEN_1 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? states_1_g : 3'h0; // @[InputUnit.scala 197:{27,27}]
  wire [2:0] _GEN_2 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? states_2_g : _GEN_1; // @[InputUnit.scala 197:{27,27}]
  wire [2:0] _GEN_3 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? states_3_g : _GEN_2; // @[InputUnit.scala 197:{27,27}]
  wire  at_dest = io_in_flit_0_bits_flow_egress_node == 2'h3; // @[InputUnit.scala 198:57]
  wire [2:0] _states_g_T = at_dest ? 3'h2 : 3'h1; // @[InputUnit.scala 199:26]
  wire [2:0] _GEN_5 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? _states_g_T : states_1_g; // @[InputUnit.scala 191:19 199:{20,20}]
  wire [2:0] _GEN_6 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? _states_g_T : states_2_g; // @[InputUnit.scala 191:19 199:{20,20}]
  wire [2:0] _GEN_7 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? _states_g_T : states_3_g; // @[InputUnit.scala 191:19 199:{20,20}]
  wire  _GEN_9 = 2'h1 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_1_vc_sel_0_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_10 = 2'h2 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_2_vc_sel_0_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_11 = 2'h3 == io_in_flit_0_bits_virt_channel_id ? 1'h0 : states_3_vc_sel_0_0; // @[InputUnit.scala 191:19 200:{45,45}]
  wire  _GEN_13 = 2'h1 == io_in_flit_0_bits_virt_channel_id | _GEN_9; // @[InputUnit.scala 203:{44,44}]
  wire  _GEN_14 = 2'h2 == io_in_flit_0_bits_virt_channel_id | _GEN_10; // @[InputUnit.scala 203:{44,44}]
  wire  _GEN_15 = 2'h3 == io_in_flit_0_bits_virt_channel_id | _GEN_11; // @[InputUnit.scala 203:{44,44}]
  wire [2:0] _GEN_41 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_5 : states_1_g; // @[InputUnit.scala 191:19 194:60]
  wire [2:0] _GEN_42 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_6 : states_2_g; // @[InputUnit.scala 191:19 194:60]
  wire [2:0] _GEN_43 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_7 : states_3_g; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_45 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_13 : states_1_vc_sel_0_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_46 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_14 : states_2_vc_sel_0_0; // @[InputUnit.scala 191:19 194:60]
  wire  _GEN_47 = io_in_flit_0_valid & io_in_flit_0_bits_head ? _GEN_15 : states_3_vc_sel_0_0; // @[InputUnit.scala 191:19 194:60]
  wire  _T_10 = route_arbiter_io_in_1_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_68 = _T_10 ? 3'h2 : _GEN_41; // @[InputUnit.scala 215:{23,29}]
  wire  _T_11 = route_arbiter_io_in_2_ready & route_arbiter_io_in_2_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_69 = _T_11 ? 3'h2 : _GEN_42; // @[InputUnit.scala 215:{23,29}]
  wire  _T_12 = route_arbiter_io_in_3_ready & route_arbiter_io_in_3_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_70 = _T_12 ? 3'h2 : _GEN_43; // @[InputUnit.scala 215:{23,29}]
  wire [2:0] _GEN_72 = 2'h1 == io_router_req_bits_src_virt_id ? states_1_g : 3'h0; // @[InputUnit.scala 224:{25,25}]
  wire [2:0] _GEN_73 = 2'h2 == io_router_req_bits_src_virt_id ? states_2_g : _GEN_72; // @[InputUnit.scala 224:{25,25}]
  wire [2:0] _GEN_74 = 2'h3 == io_router_req_bits_src_virt_id ? states_3_g : _GEN_73; // @[InputUnit.scala 224:{25,25}]
  wire [2:0] _GEN_76 = 2'h1 == io_router_req_bits_src_virt_id ? 3'h2 : _GEN_68; // @[InputUnit.scala 225:{18,18}]
  wire [2:0] _GEN_77 = 2'h2 == io_router_req_bits_src_virt_id ? 3'h2 : _GEN_69; // @[InputUnit.scala 225:{18,18}]
  wire [2:0] _GEN_78 = 2'h3 == io_router_req_bits_src_virt_id ? 3'h2 : _GEN_70; // @[InputUnit.scala 225:{18,18}]
  wire  _GEN_80 = 2'h1 == io_router_req_bits_src_virt_id ? 1'h0 : _GEN_45; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_81 = 2'h2 == io_router_req_bits_src_virt_id ? 1'h0 : _GEN_46; // @[InputUnit.scala 227:25 228:26]
  wire  _GEN_82 = 2'h3 == io_router_req_bits_src_virt_id ? 1'h0 : _GEN_47; // @[InputUnit.scala 227:25 228:26]
  wire [2:0] _GEN_84 = io_router_req_valid ? _GEN_76 : _GEN_68; // @[InputUnit.scala 222:31]
  wire [2:0] _GEN_85 = io_router_req_valid ? _GEN_77 : _GEN_69; // @[InputUnit.scala 222:31]
  wire [2:0] _GEN_86 = io_router_req_valid ? _GEN_78 : _GEN_70; // @[InputUnit.scala 222:31]
  wire  _GEN_88 = io_router_req_valid ? _GEN_80 : _GEN_45; // @[InputUnit.scala 222:31]
  wire  _GEN_89 = io_router_req_valid ? _GEN_81 : _GEN_46; // @[InputUnit.scala 222:31]
  wire  _GEN_90 = io_router_req_valid ? _GEN_82 : _GEN_47; // @[InputUnit.scala 222:31]
  reg [3:0] mask; // @[InputUnit.scala 233:21]
  wire  vcalloc_vals_1 = states_1_g == 3'h2; // @[InputUnit.scala 249:32]
  wire  vcalloc_vals_3 = states_3_g == 3'h2; // @[InputUnit.scala 249:32]
  wire  vcalloc_vals_2 = states_2_g == 3'h2; // @[InputUnit.scala 249:32]
  wire [3:0] _vcalloc_filter_T = {vcalloc_vals_3,vcalloc_vals_2,vcalloc_vals_1,1'h0}; // @[InputUnit.scala 236:59]
  wire [3:0] _vcalloc_filter_T_2 = ~mask; // @[InputUnit.scala 236:89]
  wire [3:0] _vcalloc_filter_T_3 = _vcalloc_filter_T & _vcalloc_filter_T_2; // @[InputUnit.scala 236:87]
  wire [7:0] _vcalloc_filter_T_4 = {vcalloc_vals_3,vcalloc_vals_2,vcalloc_vals_1,1'h0,_vcalloc_filter_T_3}; // @[Cat.scala 33:92]
  wire [7:0] _vcalloc_filter_T_13 = _vcalloc_filter_T_4[7] ? 8'h80 : 8'h0; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_14 = _vcalloc_filter_T_4[6] ? 8'h40 : _vcalloc_filter_T_13; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_15 = _vcalloc_filter_T_4[5] ? 8'h20 : _vcalloc_filter_T_14; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_16 = _vcalloc_filter_T_4[4] ? 8'h10 : _vcalloc_filter_T_15; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_17 = _vcalloc_filter_T_4[3] ? 8'h8 : _vcalloc_filter_T_16; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_18 = _vcalloc_filter_T_4[2] ? 8'h4 : _vcalloc_filter_T_17; // @[Mux.scala 47:70]
  wire [7:0] _vcalloc_filter_T_19 = _vcalloc_filter_T_4[1] ? 8'h2 : _vcalloc_filter_T_18; // @[Mux.scala 47:70]
  wire [7:0] vcalloc_filter = _vcalloc_filter_T_4[0] ? 8'h1 : _vcalloc_filter_T_19; // @[Mux.scala 47:70]
  wire [3:0] vcalloc_sel = vcalloc_filter[3:0] | vcalloc_filter[7:4]; // @[InputUnit.scala 237:58]
  wire [3:0] _mask_T = 4'h1 << io_router_req_bits_src_virt_id; // @[InputUnit.scala 240:18]
  wire [3:0] _mask_T_2 = _mask_T - 4'h1; // @[InputUnit.scala 240:53]
  wire  _T_25 = vcalloc_vals_1 | vcalloc_vals_2 | vcalloc_vals_3; // @[package.scala 73:59]
  wire [1:0] _mask_T_12 = vcalloc_sel[1] ? 2'h3 : 2'h0; // @[Mux.scala 27:73]
  wire [2:0] _mask_T_13 = vcalloc_sel[2] ? 3'h7 : 3'h0; // @[Mux.scala 27:73]
  wire [3:0] _mask_T_14 = vcalloc_sel[3] ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [1:0] _GEN_23 = {{1'd0}, vcalloc_sel[0]}; // @[Mux.scala 27:73]
  wire [1:0] _mask_T_15 = _GEN_23 | _mask_T_12; // @[Mux.scala 27:73]
  wire [2:0] _GEN_28 = {{1'd0}, _mask_T_15}; // @[Mux.scala 27:73]
  wire [2:0] _mask_T_16 = _GEN_28 | _mask_T_13; // @[Mux.scala 27:73]
  wire [3:0] _GEN_29 = {{1'd0}, _mask_T_16}; // @[Mux.scala 27:73]
  wire [3:0] _mask_T_17 = _GEN_29 | _mask_T_14; // @[Mux.scala 27:73]
  wire [2:0] _GEN_93 = vcalloc_vals_1 & vcalloc_sel[1] & io_vcalloc_req_ready ? 3'h3 : _GEN_84; // @[InputUnit.scala 253:{76,82}]
  wire [2:0] _GEN_94 = vcalloc_vals_2 & vcalloc_sel[2] & io_vcalloc_req_ready ? 3'h3 : _GEN_85; // @[InputUnit.scala 253:{76,82}]
  wire [2:0] _GEN_95 = vcalloc_vals_3 & vcalloc_sel[3] & io_vcalloc_req_ready ? 3'h3 : _GEN_86; // @[InputUnit.scala 253:{76,82}]
  wire [1:0] _io_debug_va_stall_T = {{1'd0}, vcalloc_vals_1}; // @[Bitwise.scala 51:90]
  wire [1:0] _io_debug_va_stall_T_2 = vcalloc_vals_2 + vcalloc_vals_3; // @[Bitwise.scala 51:90]
  wire [2:0] _io_debug_va_stall_T_4 = _io_debug_va_stall_T + _io_debug_va_stall_T_2; // @[Bitwise.scala 51:90]
  wire [2:0] _GEN_30 = {{2'd0}, io_vcalloc_req_ready}; // @[InputUnit.scala 266:47]
  wire [2:0] _io_debug_va_stall_T_7 = _io_debug_va_stall_T_4 - _GEN_30; // @[InputUnit.scala 266:47]
  wire  _T_35 = io_vcalloc_req_ready & io_vcalloc_req_valid; // @[Decoupled.scala 51:35]
  wire  credit_available = states_1_vc_sel_0_0 & io_out_credit_available_0_0; // @[InputUnit.scala 287:47]
  wire  _T_56 = salloc_arb_io_in_1_ready & salloc_arb_io_in_1_valid; // @[Decoupled.scala 51:35]
  wire  credit_available_1 = states_2_vc_sel_0_0 & io_out_credit_available_0_0; // @[InputUnit.scala 287:47]
  wire  _T_58 = salloc_arb_io_in_2_ready & salloc_arb_io_in_2_valid; // @[Decoupled.scala 51:35]
  wire  credit_available_2 = states_3_vc_sel_0_0 & io_out_credit_available_0_0; // @[InputUnit.scala 287:47]
  wire  _T_60 = salloc_arb_io_in_3_ready & salloc_arb_io_in_3_valid; // @[Decoupled.scala 51:35]
  wire  _io_debug_sa_stall_T_1 = salloc_arb_io_in_0_valid & ~salloc_arb_io_in_0_ready; // @[InputUnit.scala 301:67]
  wire  _io_debug_sa_stall_T_3 = salloc_arb_io_in_1_valid & ~salloc_arb_io_in_1_ready; // @[InputUnit.scala 301:67]
  wire  _io_debug_sa_stall_T_5 = salloc_arb_io_in_2_valid & ~salloc_arb_io_in_2_ready; // @[InputUnit.scala 301:67]
  wire  _io_debug_sa_stall_T_7 = salloc_arb_io_in_3_valid & ~salloc_arb_io_in_3_ready; // @[InputUnit.scala 301:67]
  wire [1:0] _io_debug_sa_stall_T_8 = _io_debug_sa_stall_T_1 + _io_debug_sa_stall_T_3; // @[Bitwise.scala 51:90]
  wire [1:0] _io_debug_sa_stall_T_10 = _io_debug_sa_stall_T_5 + _io_debug_sa_stall_T_7; // @[Bitwise.scala 51:90]
  wire [2:0] _io_debug_sa_stall_T_12 = _io_debug_sa_stall_T_8 + _io_debug_sa_stall_T_10; // @[Bitwise.scala 51:90]
  reg  salloc_outs_0_valid; // @[InputUnit.scala 318:8]
  reg  salloc_outs_0_flit_head; // @[InputUnit.scala 318:8]
  reg  salloc_outs_0_flit_tail; // @[InputUnit.scala 318:8]
  reg [63:0] salloc_outs_0_flit_payload; // @[InputUnit.scala 318:8]
  reg [1:0] salloc_outs_0_flit_flow_ingress_node; // @[InputUnit.scala 318:8]
  wire  _io_in_credit_return_T = salloc_arb_io_out_0_ready & salloc_arb_io_out_0_valid; // @[Decoupled.scala 51:35]
  wire  _io_in_vc_free_T_11 = salloc_arb_io_chosen_oh_0[0] & input_buffer_io_deq_0_bits_tail | salloc_arb_io_chosen_oh_0
    [1] & input_buffer_io_deq_1_bits_tail | salloc_arb_io_chosen_oh_0[2] & input_buffer_io_deq_2_bits_tail |
    salloc_arb_io_chosen_oh_0[3] & input_buffer_io_deq_3_bits_tail; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_4 = salloc_arb_io_chosen_oh_0[0] ? input_buffer_io_deq_0_bits_payload : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_5 = salloc_arb_io_chosen_oh_0[1] ? input_buffer_io_deq_1_bits_payload : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_6 = salloc_arb_io_chosen_oh_0[2] ? input_buffer_io_deq_2_bits_payload : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_7 = salloc_arb_io_chosen_oh_0[3] ? input_buffer_io_deq_3_bits_payload : 64'h0
    ; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_8 = _salloc_outs_0_flit_payload_T_4 | _salloc_outs_0_flit_payload_T_5; // @[Mux.scala 27:73]
  wire [63:0] _salloc_outs_0_flit_payload_T_9 = _salloc_outs_0_flit_payload_T_8 | _salloc_outs_0_flit_payload_T_6; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_26 = salloc_arb_io_chosen_oh_0[1] ? states_1_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_27 = salloc_arb_io_chosen_oh_0[2] ? states_2_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_28 = salloc_arb_io_chosen_oh_0[3] ? states_3_flow_ingress_node : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _salloc_outs_0_flit_flow_T_30 = _salloc_outs_0_flit_flow_T_26 | _salloc_outs_0_flit_flow_T_27; // @[Mux.scala 27:73]
  InputBuffer input_buffer ( // @[InputUnit.scala 180:28]
    .clock(input_buffer_clock),
    .reset(input_buffer_reset),
    .io_enq_0_valid(input_buffer_io_enq_0_valid),
    .io_enq_0_bits_head(input_buffer_io_enq_0_bits_head),
    .io_enq_0_bits_tail(input_buffer_io_enq_0_bits_tail),
    .io_enq_0_bits_payload(input_buffer_io_enq_0_bits_payload),
    .io_enq_0_bits_virt_channel_id(input_buffer_io_enq_0_bits_virt_channel_id),
    .io_deq_0_bits_head(input_buffer_io_deq_0_bits_head),
    .io_deq_0_bits_tail(input_buffer_io_deq_0_bits_tail),
    .io_deq_0_bits_payload(input_buffer_io_deq_0_bits_payload),
    .io_deq_1_ready(input_buffer_io_deq_1_ready),
    .io_deq_1_valid(input_buffer_io_deq_1_valid),
    .io_deq_1_bits_head(input_buffer_io_deq_1_bits_head),
    .io_deq_1_bits_tail(input_buffer_io_deq_1_bits_tail),
    .io_deq_1_bits_payload(input_buffer_io_deq_1_bits_payload),
    .io_deq_2_ready(input_buffer_io_deq_2_ready),
    .io_deq_2_valid(input_buffer_io_deq_2_valid),
    .io_deq_2_bits_head(input_buffer_io_deq_2_bits_head),
    .io_deq_2_bits_tail(input_buffer_io_deq_2_bits_tail),
    .io_deq_2_bits_payload(input_buffer_io_deq_2_bits_payload),
    .io_deq_3_ready(input_buffer_io_deq_3_ready),
    .io_deq_3_valid(input_buffer_io_deq_3_valid),
    .io_deq_3_bits_head(input_buffer_io_deq_3_bits_head),
    .io_deq_3_bits_tail(input_buffer_io_deq_3_bits_tail),
    .io_deq_3_bits_payload(input_buffer_io_deq_3_bits_payload)
  );
  Arbiter route_arbiter ( // @[InputUnit.scala 186:29]
    .io_in_1_valid(route_arbiter_io_in_1_valid),
    .io_in_2_ready(route_arbiter_io_in_2_ready),
    .io_in_2_valid(route_arbiter_io_in_2_valid),
    .io_in_3_ready(route_arbiter_io_in_3_ready),
    .io_in_3_valid(route_arbiter_io_in_3_valid),
    .io_out_valid(route_arbiter_io_out_valid),
    .io_out_bits_src_virt_id(route_arbiter_io_out_bits_src_virt_id)
  );
  SwitchArbiter_2 salloc_arb ( // @[InputUnit.scala 279:26]
    .clock(salloc_arb_clock),
    .reset(salloc_arb_reset),
    .io_in_0_ready(salloc_arb_io_in_0_ready),
    .io_in_0_valid(salloc_arb_io_in_0_valid),
    .io_in_1_ready(salloc_arb_io_in_1_ready),
    .io_in_1_valid(salloc_arb_io_in_1_valid),
    .io_in_1_bits_vc_sel_0_0(salloc_arb_io_in_1_bits_vc_sel_0_0),
    .io_in_1_bits_tail(salloc_arb_io_in_1_bits_tail),
    .io_in_2_ready(salloc_arb_io_in_2_ready),
    .io_in_2_valid(salloc_arb_io_in_2_valid),
    .io_in_2_bits_vc_sel_0_0(salloc_arb_io_in_2_bits_vc_sel_0_0),
    .io_in_2_bits_tail(salloc_arb_io_in_2_bits_tail),
    .io_in_3_ready(salloc_arb_io_in_3_ready),
    .io_in_3_valid(salloc_arb_io_in_3_valid),
    .io_in_3_bits_vc_sel_0_0(salloc_arb_io_in_3_bits_vc_sel_0_0),
    .io_in_3_bits_tail(salloc_arb_io_in_3_bits_tail),
    .io_out_0_ready(salloc_arb_io_out_0_ready),
    .io_out_0_valid(salloc_arb_io_out_0_valid),
    .io_out_0_bits_vc_sel_0_0(salloc_arb_io_out_0_bits_vc_sel_0_0),
    .io_out_0_bits_tail(salloc_arb_io_out_0_bits_tail),
    .io_chosen_oh_0(salloc_arb_io_chosen_oh_0)
  );
  assign io_router_req_valid = route_arbiter_io_out_valid; // @[InputUnit.scala 189:17]
  assign io_router_req_bits_src_virt_id = route_arbiter_io_out_bits_src_virt_id; // @[InputUnit.scala 189:17]
  assign io_vcalloc_req_valid = vcalloc_vals_1 | vcalloc_vals_2 | vcalloc_vals_3; // @[package.scala 73:59]
  assign io_vcalloc_req_bits_vc_sel_0_0 = vcalloc_sel[1] & states_1_vc_sel_0_0 | vcalloc_sel[2] & states_2_vc_sel_0_0 |
    vcalloc_sel[3] & states_3_vc_sel_0_0; // @[Mux.scala 27:73]
  assign io_salloc_req_0_valid = salloc_arb_io_out_0_valid; // @[InputUnit.scala 302:17 303:19 305:35]
  assign io_salloc_req_0_bits_vc_sel_0_0 = salloc_arb_io_out_0_bits_vc_sel_0_0; // @[InputUnit.scala 302:17]
  assign io_salloc_req_0_bits_tail = salloc_arb_io_out_0_bits_tail; // @[InputUnit.scala 302:17]
  assign io_out_0_valid = salloc_outs_0_valid; // @[InputUnit.scala 349:21]
  assign io_out_0_bits_flit_head = salloc_outs_0_flit_head; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_flit_tail = salloc_outs_0_flit_tail; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_flit_payload = salloc_outs_0_flit_payload; // @[InputUnit.scala 350:25]
  assign io_out_0_bits_flit_flow_ingress_node = salloc_outs_0_flit_flow_ingress_node; // @[InputUnit.scala 350:25]
  assign io_debug_va_stall = _io_debug_va_stall_T_7[1:0]; // @[InputUnit.scala 266:21]
  assign io_debug_sa_stall = _io_debug_sa_stall_T_12[1:0]; // @[InputUnit.scala 301:21]
  assign io_in_credit_return = _io_in_credit_return_T ? salloc_arb_io_chosen_oh_0 : 4'h0; // @[InputUnit.scala 322:8]
  assign io_in_vc_free = _io_in_credit_return_T & _io_in_vc_free_T_11 ? salloc_arb_io_chosen_oh_0 : 4'h0; // @[InputUnit.scala 325:8]
  assign input_buffer_clock = clock;
  assign input_buffer_reset = reset;
  assign input_buffer_io_enq_0_valid = io_in_flit_0_valid; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_head = io_in_flit_0_bits_head; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_tail = io_in_flit_0_bits_tail; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_payload = io_in_flit_0_bits_payload; // @[InputUnit.scala 182:28]
  assign input_buffer_io_enq_0_bits_virt_channel_id = io_in_flit_0_bits_virt_channel_id; // @[InputUnit.scala 182:28]
  assign input_buffer_io_deq_1_ready = salloc_arb_io_in_1_ready; // @[InputUnit.scala 295:36]
  assign input_buffer_io_deq_2_ready = salloc_arb_io_in_2_ready; // @[InputUnit.scala 295:36]
  assign input_buffer_io_deq_3_ready = salloc_arb_io_in_3_ready; // @[InputUnit.scala 295:36]
  assign route_arbiter_io_in_1_valid = states_1_g == 3'h1; // @[InputUnit.scala 212:22]
  assign route_arbiter_io_in_2_valid = states_2_g == 3'h1; // @[InputUnit.scala 212:22]
  assign route_arbiter_io_in_3_valid = states_3_g == 3'h1; // @[InputUnit.scala 212:22]
  assign salloc_arb_clock = clock;
  assign salloc_arb_reset = reset;
  assign salloc_arb_io_in_0_valid = 1'h0; // @[InputUnit.scala 297:15]
  assign salloc_arb_io_in_1_valid = states_1_g == 3'h3 & credit_available & input_buffer_io_deq_1_valid; // @[InputUnit.scala 288:50]
  assign salloc_arb_io_in_1_bits_vc_sel_0_0 = states_1_vc_sel_0_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_1_bits_tail = input_buffer_io_deq_1_bits_tail; // @[InputUnit.scala 291:19]
  assign salloc_arb_io_in_2_valid = states_2_g == 3'h3 & credit_available_1 & input_buffer_io_deq_2_valid; // @[InputUnit.scala 288:50]
  assign salloc_arb_io_in_2_bits_vc_sel_0_0 = states_2_vc_sel_0_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_2_bits_tail = input_buffer_io_deq_2_bits_tail; // @[InputUnit.scala 291:19]
  assign salloc_arb_io_in_3_valid = states_3_g == 3'h3 & credit_available_2 & input_buffer_io_deq_3_valid; // @[InputUnit.scala 288:50]
  assign salloc_arb_io_in_3_bits_vc_sel_0_0 = states_3_vc_sel_0_0; // @[InputUnit.scala 289:21]
  assign salloc_arb_io_in_3_bits_tail = input_buffer_io_deq_3_bits_tail; // @[InputUnit.scala 291:19]
  assign salloc_arb_io_out_0_ready = io_salloc_req_0_ready; // @[InputUnit.scala 302:17 303:19 304:39]
  always @(posedge clock) begin
    if (reset) begin // @[InputUnit.scala 377:23]
      states_1_g <= 3'h0; // @[InputUnit.scala 378:24]
    end else if (_T_56 & input_buffer_io_deq_1_bits_tail) begin // @[InputUnit.scala 292:35]
      states_1_g <= 3'h0; // @[InputUnit.scala 293:13]
    end else if (_T_35) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_g <= 3'h3; // @[InputUnit.scala 272:21]
      end else begin
        states_1_g <= _GEN_93;
      end
    end else begin
      states_1_g <= _GEN_93;
    end
    if (_T_35) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[1]) begin // @[InputUnit.scala 270:29]
        states_1_vc_sel_0_0 <= io_vcalloc_resp_vc_sel_0_0; // @[InputUnit.scala 271:26]
      end else begin
        states_1_vc_sel_0_0 <= _GEN_88;
      end
    end else begin
      states_1_vc_sel_0_0 <= _GEN_88;
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h1 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_1_flow_ingress_node <= io_in_flit_0_bits_flow_ingress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (reset) begin // @[InputUnit.scala 377:23]
      states_2_g <= 3'h0; // @[InputUnit.scala 378:24]
    end else if (_T_58 & input_buffer_io_deq_2_bits_tail) begin // @[InputUnit.scala 292:35]
      states_2_g <= 3'h0; // @[InputUnit.scala 293:13]
    end else if (_T_35) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_g <= 3'h3; // @[InputUnit.scala 272:21]
      end else begin
        states_2_g <= _GEN_94;
      end
    end else begin
      states_2_g <= _GEN_94;
    end
    if (_T_35) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[2]) begin // @[InputUnit.scala 270:29]
        states_2_vc_sel_0_0 <= io_vcalloc_resp_vc_sel_0_0; // @[InputUnit.scala 271:26]
      end else begin
        states_2_vc_sel_0_0 <= _GEN_89;
      end
    end else begin
      states_2_vc_sel_0_0 <= _GEN_89;
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h2 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_2_flow_ingress_node <= io_in_flit_0_bits_flow_ingress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (reset) begin // @[InputUnit.scala 377:23]
      states_3_g <= 3'h0; // @[InputUnit.scala 378:24]
    end else if (_T_60 & input_buffer_io_deq_3_bits_tail) begin // @[InputUnit.scala 292:35]
      states_3_g <= 3'h0; // @[InputUnit.scala 293:13]
    end else if (_T_35) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_g <= 3'h3; // @[InputUnit.scala 272:21]
      end else begin
        states_3_g <= _GEN_95;
      end
    end else begin
      states_3_g <= _GEN_95;
    end
    if (_T_35) begin // @[InputUnit.scala 268:32]
      if (vcalloc_sel[3]) begin // @[InputUnit.scala 270:29]
        states_3_vc_sel_0_0 <= io_vcalloc_resp_vc_sel_0_0; // @[InputUnit.scala 271:26]
      end else begin
        states_3_vc_sel_0_0 <= _GEN_90;
      end
    end else begin
      states_3_vc_sel_0_0 <= _GEN_90;
    end
    if (io_in_flit_0_valid & io_in_flit_0_bits_head) begin // @[InputUnit.scala 194:60]
      if (2'h3 == io_in_flit_0_bits_virt_channel_id) begin // @[InputUnit.scala 206:23]
        states_3_flow_ingress_node <= io_in_flit_0_bits_flow_ingress_node; // @[InputUnit.scala 206:23]
      end
    end
    if (reset) begin // @[InputUnit.scala 233:21]
      mask <= 4'h0; // @[InputUnit.scala 233:21]
    end else if (io_router_req_valid) begin // @[InputUnit.scala 239:31]
      mask <= _mask_T_2; // @[InputUnit.scala 240:10]
    end else if (_T_25) begin // @[InputUnit.scala 241:34]
      mask <= _mask_T_17; // @[InputUnit.scala 242:10]
    end
    salloc_outs_0_valid <= salloc_arb_io_out_0_ready & salloc_arb_io_out_0_valid; // @[Decoupled.scala 51:35]
    salloc_outs_0_flit_head <= salloc_arb_io_chosen_oh_0[0] & input_buffer_io_deq_0_bits_head |
      salloc_arb_io_chosen_oh_0[1] & input_buffer_io_deq_1_bits_head | salloc_arb_io_chosen_oh_0[2] &
      input_buffer_io_deq_2_bits_head | salloc_arb_io_chosen_oh_0[3] & input_buffer_io_deq_3_bits_head; // @[Mux.scala 27:73]
    salloc_outs_0_flit_tail <= salloc_arb_io_chosen_oh_0[0] & input_buffer_io_deq_0_bits_tail |
      salloc_arb_io_chosen_oh_0[1] & input_buffer_io_deq_1_bits_tail | salloc_arb_io_chosen_oh_0[2] &
      input_buffer_io_deq_2_bits_tail | salloc_arb_io_chosen_oh_0[3] & input_buffer_io_deq_3_bits_tail; // @[Mux.scala 27:73]
    salloc_outs_0_flit_payload <= _salloc_outs_0_flit_payload_T_9 | _salloc_outs_0_flit_payload_T_7; // @[Mux.scala 27:73]
    salloc_outs_0_flit_flow_ingress_node <= _salloc_outs_0_flit_flow_T_30 | _salloc_outs_0_flit_flow_T_28; // @[Mux.scala 27:73]
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T & _T_3 & ~(_GEN_3 == 3'h0)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:197 assert(states(id).g === g_i)\n"); // @[InputUnit.scala 197:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_router_req_valid & _T_3 & ~(_GEN_74 == 3'h1)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:224 assert(states(id).g === g_r)\n"); // @[InputUnit.scala 224:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_35 & vcalloc_sel[0] & _T_3) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:274 assert(states(i).g === g_v)\n"); // @[InputUnit.scala 274:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_35 & vcalloc_sel[1] & _T_3 & ~vcalloc_vals_1) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:274 assert(states(i).g === g_v)\n"); // @[InputUnit.scala 274:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_35 & vcalloc_sel[2] & _T_3 & ~vcalloc_vals_2) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:274 assert(states(i).g === g_v)\n"); // @[InputUnit.scala 274:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_35 & vcalloc_sel[3] & _T_3 & ~vcalloc_vals_3) begin
          $fwrite(32'h80000002,"Assertion failed\n    at InputUnit.scala:274 assert(states(i).g === g_v)\n"); // @[InputUnit.scala 274:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  states_1_g = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  states_1_vc_sel_0_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  states_1_flow_ingress_node = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  states_2_g = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  states_2_vc_sel_0_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  states_2_flow_ingress_node = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  states_3_g = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  states_3_vc_sel_0_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  states_3_flow_ingress_node = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  mask = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  salloc_outs_0_valid = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  salloc_outs_0_flit_head = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  salloc_outs_0_flit_tail = _RAND_12[0:0];
  _RAND_13 = {2{`RANDOM}};
  salloc_outs_0_flit_payload = _RAND_13[63:0];
  _RAND_14 = {1{`RANDOM}};
  salloc_outs_0_flit_flow_ingress_node = _RAND_14[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (_T & ~reset) begin
      assert(1'h1); // @[InputUnit.scala 196:13]
    end
    //
    if (_T & _T_3) begin
      assert(_GEN_3 == 3'h0); // @[InputUnit.scala 197:13]
    end
    //
    if (io_router_req_valid & _T_3) begin
      assert(_GEN_74 == 3'h1); // @[InputUnit.scala 224:11]
    end
    //
    if (_T_35 & vcalloc_sel[0] & _T_3) begin
      assert(1'h0); // @[InputUnit.scala 274:17]
    end
    //
    if (_T_35 & vcalloc_sel[1] & _T_3) begin
      assert(vcalloc_vals_1); // @[InputUnit.scala 274:17]
    end
    //
    if (_T_35 & vcalloc_sel[2] & _T_3) begin
      assert(vcalloc_vals_2); // @[InputUnit.scala 274:17]
    end
    //
    if (_T_35 & vcalloc_sel[3] & _T_3) begin
      assert(vcalloc_vals_3); // @[InputUnit.scala 274:17]
    end
  end
endmodule
module Router_3(
  input         clock,
  input         reset,
  output [1:0]  auto_debug_out_va_stall_0,
  output [1:0]  auto_debug_out_va_stall_1,
  output [1:0]  auto_debug_out_sa_stall_0,
  output [1:0]  auto_debug_out_sa_stall_1,
  output        auto_egress_nodes_out_flit_valid,
  output        auto_egress_nodes_out_flit_bits_head,
  output        auto_egress_nodes_out_flit_bits_tail,
  output [63:0] auto_egress_nodes_out_flit_bits_payload,
  output        auto_egress_nodes_out_flit_bits_ingress_id,
  input         auto_dest_nodes_in_1_flit_0_valid,
  input         auto_dest_nodes_in_1_flit_0_bits_head,
  input         auto_dest_nodes_in_1_flit_0_bits_tail,
  input  [63:0] auto_dest_nodes_in_1_flit_0_bits_payload,
  input  [1:0]  auto_dest_nodes_in_1_flit_0_bits_flow_ingress_node,
  input  [1:0]  auto_dest_nodes_in_1_flit_0_bits_flow_egress_node,
  input  [1:0]  auto_dest_nodes_in_1_flit_0_bits_virt_channel_id,
  output [3:0]  auto_dest_nodes_in_1_credit_return,
  output [3:0]  auto_dest_nodes_in_1_vc_free,
  input         auto_dest_nodes_in_0_flit_0_valid,
  input         auto_dest_nodes_in_0_flit_0_bits_head,
  input         auto_dest_nodes_in_0_flit_0_bits_tail,
  input  [63:0] auto_dest_nodes_in_0_flit_0_bits_payload,
  input  [1:0]  auto_dest_nodes_in_0_flit_0_bits_flow_ingress_node,
  input  [1:0]  auto_dest_nodes_in_0_flit_0_bits_flow_egress_node,
  input  [1:0]  auto_dest_nodes_in_0_flit_0_bits_virt_channel_id,
  output [3:0]  auto_dest_nodes_in_0_credit_return,
  output [3:0]  auto_dest_nodes_in_0_vc_free
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  monitor_clock; // @[Nodes.scala 24:25]
  wire  monitor_reset; // @[Nodes.scala 24:25]
  wire  monitor_io_in_flit_0_valid; // @[Nodes.scala 24:25]
  wire  monitor_io_in_flit_0_bits_head; // @[Nodes.scala 24:25]
  wire  monitor_io_in_flit_0_bits_tail; // @[Nodes.scala 24:25]
  wire [1:0] monitor_io_in_flit_0_bits_flow_ingress_node; // @[Nodes.scala 24:25]
  wire [1:0] monitor_io_in_flit_0_bits_flow_egress_node; // @[Nodes.scala 24:25]
  wire [1:0] monitor_io_in_flit_0_bits_virt_channel_id; // @[Nodes.scala 24:25]
  wire  monitor_1_clock; // @[Nodes.scala 24:25]
  wire  monitor_1_reset; // @[Nodes.scala 24:25]
  wire  monitor_1_io_in_flit_0_valid; // @[Nodes.scala 24:25]
  wire  monitor_1_io_in_flit_0_bits_head; // @[Nodes.scala 24:25]
  wire  monitor_1_io_in_flit_0_bits_tail; // @[Nodes.scala 24:25]
  wire [1:0] monitor_1_io_in_flit_0_bits_flow_ingress_node; // @[Nodes.scala 24:25]
  wire [1:0] monitor_1_io_in_flit_0_bits_flow_egress_node; // @[Nodes.scala 24:25]
  wire [1:0] monitor_1_io_in_flit_0_bits_virt_channel_id; // @[Nodes.scala 24:25]
  wire  input_unit_0_from_0_clock; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_reset; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_router_req_valid; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_0_io_router_req_bits_src_virt_id; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_req_ready; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_req_valid; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_vcalloc_resp_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_out_credit_available_0_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_salloc_req_0_ready; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_salloc_req_0_valid; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_salloc_req_0_bits_tail; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_out_0_valid; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_out_0_bits_flit_head; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_out_0_bits_flit_tail; // @[Router.scala 112:13]
  wire [63:0] input_unit_0_from_0_io_out_0_bits_flit_payload; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_0_io_out_0_bits_flit_flow_ingress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_0_io_debug_va_stall; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_0_io_debug_sa_stall; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_in_flit_0_valid; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_in_flit_0_bits_head; // @[Router.scala 112:13]
  wire  input_unit_0_from_0_io_in_flit_0_bits_tail; // @[Router.scala 112:13]
  wire [63:0] input_unit_0_from_0_io_in_flit_0_bits_payload; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_0_io_in_flit_0_bits_flow_ingress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_0_io_in_flit_0_bits_flow_egress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_0_from_0_io_in_flit_0_bits_virt_channel_id; // @[Router.scala 112:13]
  wire [3:0] input_unit_0_from_0_io_in_credit_return; // @[Router.scala 112:13]
  wire [3:0] input_unit_0_from_0_io_in_vc_free; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_clock; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_reset; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_router_req_valid; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_2_io_router_req_bits_src_virt_id; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_req_ready; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_req_valid; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_vcalloc_resp_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_out_credit_available_0_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_salloc_req_0_ready; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_salloc_req_0_valid; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_0_0; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_salloc_req_0_bits_tail; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_out_0_valid; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_out_0_bits_flit_head; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_out_0_bits_flit_tail; // @[Router.scala 112:13]
  wire [63:0] input_unit_1_from_2_io_out_0_bits_flit_payload; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_2_io_out_0_bits_flit_flow_ingress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_2_io_debug_va_stall; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_2_io_debug_sa_stall; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_in_flit_0_valid; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_in_flit_0_bits_head; // @[Router.scala 112:13]
  wire  input_unit_1_from_2_io_in_flit_0_bits_tail; // @[Router.scala 112:13]
  wire [63:0] input_unit_1_from_2_io_in_flit_0_bits_payload; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_2_io_in_flit_0_bits_flow_ingress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_2_io_in_flit_0_bits_flow_egress_node; // @[Router.scala 112:13]
  wire [1:0] input_unit_1_from_2_io_in_flit_0_bits_virt_channel_id; // @[Router.scala 112:13]
  wire [3:0] input_unit_1_from_2_io_in_credit_return; // @[Router.scala 112:13]
  wire [3:0] input_unit_1_from_2_io_in_vc_free; // @[Router.scala 112:13]
  wire  egress_unit_0_to_1_clock; // @[Router.scala 125:13]
  wire  egress_unit_0_to_1_reset; // @[Router.scala 125:13]
  wire  egress_unit_0_to_1_io_in_0_valid; // @[Router.scala 125:13]
  wire  egress_unit_0_to_1_io_in_0_bits_head; // @[Router.scala 125:13]
  wire  egress_unit_0_to_1_io_in_0_bits_tail; // @[Router.scala 125:13]
  wire [63:0] egress_unit_0_to_1_io_in_0_bits_payload; // @[Router.scala 125:13]
  wire [1:0] egress_unit_0_to_1_io_in_0_bits_flow_ingress_node; // @[Router.scala 125:13]
  wire  egress_unit_0_to_1_io_credit_available_0; // @[Router.scala 125:13]
  wire  egress_unit_0_to_1_io_channel_status_0_occupied; // @[Router.scala 125:13]
  wire  egress_unit_0_to_1_io_allocs_0_alloc; // @[Router.scala 125:13]
  wire  egress_unit_0_to_1_io_credit_alloc_0_alloc; // @[Router.scala 125:13]
  wire  egress_unit_0_to_1_io_credit_alloc_0_tail; // @[Router.scala 125:13]
  wire  egress_unit_0_to_1_io_out_valid; // @[Router.scala 125:13]
  wire  egress_unit_0_to_1_io_out_bits_head; // @[Router.scala 125:13]
  wire  egress_unit_0_to_1_io_out_bits_tail; // @[Router.scala 125:13]
  wire [63:0] egress_unit_0_to_1_io_out_bits_payload; // @[Router.scala 125:13]
  wire  egress_unit_0_to_1_io_out_bits_ingress_id; // @[Router.scala 125:13]
  wire  switch_clock; // @[Router.scala 129:24]
  wire  switch_reset; // @[Router.scala 129:24]
  wire  switch_io_in_1_0_valid; // @[Router.scala 129:24]
  wire  switch_io_in_1_0_bits_flit_head; // @[Router.scala 129:24]
  wire  switch_io_in_1_0_bits_flit_tail; // @[Router.scala 129:24]
  wire [63:0] switch_io_in_1_0_bits_flit_payload; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_1_0_bits_flit_flow_ingress_node; // @[Router.scala 129:24]
  wire  switch_io_in_0_0_valid; // @[Router.scala 129:24]
  wire  switch_io_in_0_0_bits_flit_head; // @[Router.scala 129:24]
  wire  switch_io_in_0_0_bits_flit_tail; // @[Router.scala 129:24]
  wire [63:0] switch_io_in_0_0_bits_flit_payload; // @[Router.scala 129:24]
  wire [1:0] switch_io_in_0_0_bits_flit_flow_ingress_node; // @[Router.scala 129:24]
  wire  switch_io_out_0_0_valid; // @[Router.scala 129:24]
  wire  switch_io_out_0_0_bits_head; // @[Router.scala 129:24]
  wire  switch_io_out_0_0_bits_tail; // @[Router.scala 129:24]
  wire [63:0] switch_io_out_0_0_bits_payload; // @[Router.scala 129:24]
  wire [1:0] switch_io_out_0_0_bits_flow_ingress_node; // @[Router.scala 129:24]
  wire  switch_io_sel_0_0_1_0; // @[Router.scala 129:24]
  wire  switch_io_sel_0_0_0_0; // @[Router.scala 129:24]
  wire  switch_allocator_clock; // @[Router.scala 130:34]
  wire  switch_allocator_reset; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_ready; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_valid; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_vc_sel_0_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_1_0_bits_tail; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_ready; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_valid; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_vc_sel_0_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_req_0_0_bits_tail; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_0_0_alloc; // @[Router.scala 130:34]
  wire  switch_allocator_io_credit_alloc_0_0_tail; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_0_0_1_0; // @[Router.scala 130:34]
  wire  switch_allocator_io_switch_sel_0_0_0_0; // @[Router.scala 130:34]
  wire  vc_allocator_clock; // @[Router.scala 131:30]
  wire  vc_allocator_reset; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_ready; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_valid; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_1_bits_vc_sel_0_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_ready; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_valid; // @[Router.scala 131:30]
  wire  vc_allocator_io_req_0_bits_vc_sel_0_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_1_vc_sel_0_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_resp_0_vc_sel_0_0; // @[Router.scala 131:30]
  wire  vc_allocator_io_channel_status_0_0_occupied; // @[Router.scala 131:30]
  wire  vc_allocator_io_out_allocs_0_0_alloc; // @[Router.scala 131:30]
  wire  route_computer_clock; // @[Router.scala 134:32]
  wire  route_computer_reset; // @[Router.scala 134:32]
  wire  route_computer_io_req_1_valid; // @[Router.scala 134:32]
  wire  route_computer_io_req_0_valid; // @[Router.scala 134:32]
  wire [19:0] plusarg_reader_out; // @[PlusArg.scala 80:11]
  wire  _fires_count_T = vc_allocator_io_req_0_ready & vc_allocator_io_req_0_valid; // @[Decoupled.scala 51:35]
  wire  _fires_count_T_1 = vc_allocator_io_req_1_ready & vc_allocator_io_req_1_valid; // @[Decoupled.scala 51:35]
  reg  switch_io_sel_REG_0_0_1_0; // @[Router.scala 176:14]
  reg  switch_io_sel_REG_0_0_0_0; // @[Router.scala 176:14]
  reg [63:0] debug_tsc; // @[Router.scala 193:28]
  wire [63:0] _debug_tsc_T_1 = debug_tsc + 64'h1; // @[Router.scala 194:28]
  reg [63:0] debug_sample; // @[Router.scala 195:31]
  wire [63:0] _debug_sample_T_1 = debug_sample + 64'h1; // @[Router.scala 196:34]
  wire [19:0] _T_1 = plusarg_reader_out - 20'h1; // @[Router.scala 198:40]
  wire [63:0] _GEN_4 = {{44'd0}, _T_1}; // @[Router.scala 198:24]
  wire  _T_2 = debug_sample == _GEN_4; // @[Router.scala 198:24]
  reg [63:0] util_ctr; // @[Router.scala 201:29]
  reg  fired; // @[Router.scala 202:26]
  wire [63:0] _GEN_5 = {{63'd0}, auto_dest_nodes_in_0_flit_0_valid}; // @[Router.scala 203:28]
  wire [63:0] _util_ctr_T_1 = util_ctr + _GEN_5; // @[Router.scala 203:28]
  wire  _T_8 = plusarg_reader_out != 20'h0 & _T_2 & fired; // @[Router.scala 205:71]
  reg [63:0] util_ctr_1; // @[Router.scala 201:29]
  reg  fired_1; // @[Router.scala 202:26]
  wire [63:0] _GEN_7 = {{63'd0}, auto_dest_nodes_in_1_flit_0_valid}; // @[Router.scala 203:28]
  wire [63:0] _util_ctr_T_3 = util_ctr_1 + _GEN_7; // @[Router.scala 203:28]
  wire  _T_16 = plusarg_reader_out != 20'h0 & _T_2 & fired_1; // @[Router.scala 205:71]
  wire  x1_flit_valid = egress_unit_0_to_1_io_out_valid; // @[Nodes.scala 1212:84 Router.scala 144:65]
  reg [63:0] util_ctr_2; // @[Router.scala 201:29]
  reg  fired_2; // @[Router.scala 202:26]
  wire [63:0] _GEN_9 = {{63'd0}, x1_flit_valid}; // @[Router.scala 203:28]
  wire [63:0] _util_ctr_T_5 = util_ctr_2 + _GEN_9; // @[Router.scala 203:28]
  wire  _T_25 = plusarg_reader_out != 20'h0 & _T_2 & fired_2; // @[Router.scala 205:71]
  wire [1:0] fires_count = _fires_count_T + _fires_count_T_1; // @[Bitwise.scala 51:90]
  NoCMonitor_2 monitor ( // @[Nodes.scala 24:25]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_flit_0_valid(monitor_io_in_flit_0_valid),
    .io_in_flit_0_bits_head(monitor_io_in_flit_0_bits_head),
    .io_in_flit_0_bits_tail(monitor_io_in_flit_0_bits_tail),
    .io_in_flit_0_bits_flow_ingress_node(monitor_io_in_flit_0_bits_flow_ingress_node),
    .io_in_flit_0_bits_flow_egress_node(monitor_io_in_flit_0_bits_flow_egress_node),
    .io_in_flit_0_bits_virt_channel_id(monitor_io_in_flit_0_bits_virt_channel_id)
  );
  NoCMonitor_3 monitor_1 ( // @[Nodes.scala 24:25]
    .clock(monitor_1_clock),
    .reset(monitor_1_reset),
    .io_in_flit_0_valid(monitor_1_io_in_flit_0_valid),
    .io_in_flit_0_bits_head(monitor_1_io_in_flit_0_bits_head),
    .io_in_flit_0_bits_tail(monitor_1_io_in_flit_0_bits_tail),
    .io_in_flit_0_bits_flow_ingress_node(monitor_1_io_in_flit_0_bits_flow_ingress_node),
    .io_in_flit_0_bits_flow_egress_node(monitor_1_io_in_flit_0_bits_flow_egress_node),
    .io_in_flit_0_bits_virt_channel_id(monitor_1_io_in_flit_0_bits_virt_channel_id)
  );
  InputUnit_2 input_unit_0_from_0 ( // @[Router.scala 112:13]
    .clock(input_unit_0_from_0_clock),
    .reset(input_unit_0_from_0_reset),
    .io_router_req_valid(input_unit_0_from_0_io_router_req_valid),
    .io_router_req_bits_src_virt_id(input_unit_0_from_0_io_router_req_bits_src_virt_id),
    .io_vcalloc_req_ready(input_unit_0_from_0_io_vcalloc_req_ready),
    .io_vcalloc_req_valid(input_unit_0_from_0_io_vcalloc_req_valid),
    .io_vcalloc_req_bits_vc_sel_0_0(input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_0),
    .io_vcalloc_resp_vc_sel_0_0(input_unit_0_from_0_io_vcalloc_resp_vc_sel_0_0),
    .io_out_credit_available_0_0(input_unit_0_from_0_io_out_credit_available_0_0),
    .io_salloc_req_0_ready(input_unit_0_from_0_io_salloc_req_0_ready),
    .io_salloc_req_0_valid(input_unit_0_from_0_io_salloc_req_0_valid),
    .io_salloc_req_0_bits_vc_sel_0_0(input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_0),
    .io_salloc_req_0_bits_tail(input_unit_0_from_0_io_salloc_req_0_bits_tail),
    .io_out_0_valid(input_unit_0_from_0_io_out_0_valid),
    .io_out_0_bits_flit_head(input_unit_0_from_0_io_out_0_bits_flit_head),
    .io_out_0_bits_flit_tail(input_unit_0_from_0_io_out_0_bits_flit_tail),
    .io_out_0_bits_flit_payload(input_unit_0_from_0_io_out_0_bits_flit_payload),
    .io_out_0_bits_flit_flow_ingress_node(input_unit_0_from_0_io_out_0_bits_flit_flow_ingress_node),
    .io_debug_va_stall(input_unit_0_from_0_io_debug_va_stall),
    .io_debug_sa_stall(input_unit_0_from_0_io_debug_sa_stall),
    .io_in_flit_0_valid(input_unit_0_from_0_io_in_flit_0_valid),
    .io_in_flit_0_bits_head(input_unit_0_from_0_io_in_flit_0_bits_head),
    .io_in_flit_0_bits_tail(input_unit_0_from_0_io_in_flit_0_bits_tail),
    .io_in_flit_0_bits_payload(input_unit_0_from_0_io_in_flit_0_bits_payload),
    .io_in_flit_0_bits_flow_ingress_node(input_unit_0_from_0_io_in_flit_0_bits_flow_ingress_node),
    .io_in_flit_0_bits_flow_egress_node(input_unit_0_from_0_io_in_flit_0_bits_flow_egress_node),
    .io_in_flit_0_bits_virt_channel_id(input_unit_0_from_0_io_in_flit_0_bits_virt_channel_id),
    .io_in_credit_return(input_unit_0_from_0_io_in_credit_return),
    .io_in_vc_free(input_unit_0_from_0_io_in_vc_free)
  );
  InputUnit_2 input_unit_1_from_2 ( // @[Router.scala 112:13]
    .clock(input_unit_1_from_2_clock),
    .reset(input_unit_1_from_2_reset),
    .io_router_req_valid(input_unit_1_from_2_io_router_req_valid),
    .io_router_req_bits_src_virt_id(input_unit_1_from_2_io_router_req_bits_src_virt_id),
    .io_vcalloc_req_ready(input_unit_1_from_2_io_vcalloc_req_ready),
    .io_vcalloc_req_valid(input_unit_1_from_2_io_vcalloc_req_valid),
    .io_vcalloc_req_bits_vc_sel_0_0(input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_0_0),
    .io_vcalloc_resp_vc_sel_0_0(input_unit_1_from_2_io_vcalloc_resp_vc_sel_0_0),
    .io_out_credit_available_0_0(input_unit_1_from_2_io_out_credit_available_0_0),
    .io_salloc_req_0_ready(input_unit_1_from_2_io_salloc_req_0_ready),
    .io_salloc_req_0_valid(input_unit_1_from_2_io_salloc_req_0_valid),
    .io_salloc_req_0_bits_vc_sel_0_0(input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_0_0),
    .io_salloc_req_0_bits_tail(input_unit_1_from_2_io_salloc_req_0_bits_tail),
    .io_out_0_valid(input_unit_1_from_2_io_out_0_valid),
    .io_out_0_bits_flit_head(input_unit_1_from_2_io_out_0_bits_flit_head),
    .io_out_0_bits_flit_tail(input_unit_1_from_2_io_out_0_bits_flit_tail),
    .io_out_0_bits_flit_payload(input_unit_1_from_2_io_out_0_bits_flit_payload),
    .io_out_0_bits_flit_flow_ingress_node(input_unit_1_from_2_io_out_0_bits_flit_flow_ingress_node),
    .io_debug_va_stall(input_unit_1_from_2_io_debug_va_stall),
    .io_debug_sa_stall(input_unit_1_from_2_io_debug_sa_stall),
    .io_in_flit_0_valid(input_unit_1_from_2_io_in_flit_0_valid),
    .io_in_flit_0_bits_head(input_unit_1_from_2_io_in_flit_0_bits_head),
    .io_in_flit_0_bits_tail(input_unit_1_from_2_io_in_flit_0_bits_tail),
    .io_in_flit_0_bits_payload(input_unit_1_from_2_io_in_flit_0_bits_payload),
    .io_in_flit_0_bits_flow_ingress_node(input_unit_1_from_2_io_in_flit_0_bits_flow_ingress_node),
    .io_in_flit_0_bits_flow_egress_node(input_unit_1_from_2_io_in_flit_0_bits_flow_egress_node),
    .io_in_flit_0_bits_virt_channel_id(input_unit_1_from_2_io_in_flit_0_bits_virt_channel_id),
    .io_in_credit_return(input_unit_1_from_2_io_in_credit_return),
    .io_in_vc_free(input_unit_1_from_2_io_in_vc_free)
  );
  EgressUnit egress_unit_0_to_1 ( // @[Router.scala 125:13]
    .clock(egress_unit_0_to_1_clock),
    .reset(egress_unit_0_to_1_reset),
    .io_in_0_valid(egress_unit_0_to_1_io_in_0_valid),
    .io_in_0_bits_head(egress_unit_0_to_1_io_in_0_bits_head),
    .io_in_0_bits_tail(egress_unit_0_to_1_io_in_0_bits_tail),
    .io_in_0_bits_payload(egress_unit_0_to_1_io_in_0_bits_payload),
    .io_in_0_bits_flow_ingress_node(egress_unit_0_to_1_io_in_0_bits_flow_ingress_node),
    .io_credit_available_0(egress_unit_0_to_1_io_credit_available_0),
    .io_channel_status_0_occupied(egress_unit_0_to_1_io_channel_status_0_occupied),
    .io_allocs_0_alloc(egress_unit_0_to_1_io_allocs_0_alloc),
    .io_credit_alloc_0_alloc(egress_unit_0_to_1_io_credit_alloc_0_alloc),
    .io_credit_alloc_0_tail(egress_unit_0_to_1_io_credit_alloc_0_tail),
    .io_out_valid(egress_unit_0_to_1_io_out_valid),
    .io_out_bits_head(egress_unit_0_to_1_io_out_bits_head),
    .io_out_bits_tail(egress_unit_0_to_1_io_out_bits_tail),
    .io_out_bits_payload(egress_unit_0_to_1_io_out_bits_payload),
    .io_out_bits_ingress_id(egress_unit_0_to_1_io_out_bits_ingress_id)
  );
  Switch_1 switch ( // @[Router.scala 129:24]
    .clock(switch_clock),
    .reset(switch_reset),
    .io_in_1_0_valid(switch_io_in_1_0_valid),
    .io_in_1_0_bits_flit_head(switch_io_in_1_0_bits_flit_head),
    .io_in_1_0_bits_flit_tail(switch_io_in_1_0_bits_flit_tail),
    .io_in_1_0_bits_flit_payload(switch_io_in_1_0_bits_flit_payload),
    .io_in_1_0_bits_flit_flow_ingress_node(switch_io_in_1_0_bits_flit_flow_ingress_node),
    .io_in_0_0_valid(switch_io_in_0_0_valid),
    .io_in_0_0_bits_flit_head(switch_io_in_0_0_bits_flit_head),
    .io_in_0_0_bits_flit_tail(switch_io_in_0_0_bits_flit_tail),
    .io_in_0_0_bits_flit_payload(switch_io_in_0_0_bits_flit_payload),
    .io_in_0_0_bits_flit_flow_ingress_node(switch_io_in_0_0_bits_flit_flow_ingress_node),
    .io_out_0_0_valid(switch_io_out_0_0_valid),
    .io_out_0_0_bits_head(switch_io_out_0_0_bits_head),
    .io_out_0_0_bits_tail(switch_io_out_0_0_bits_tail),
    .io_out_0_0_bits_payload(switch_io_out_0_0_bits_payload),
    .io_out_0_0_bits_flow_ingress_node(switch_io_out_0_0_bits_flow_ingress_node),
    .io_sel_0_0_1_0(switch_io_sel_0_0_1_0),
    .io_sel_0_0_0_0(switch_io_sel_0_0_0_0)
  );
  SwitchAllocator_1 switch_allocator ( // @[Router.scala 130:34]
    .clock(switch_allocator_clock),
    .reset(switch_allocator_reset),
    .io_req_1_0_ready(switch_allocator_io_req_1_0_ready),
    .io_req_1_0_valid(switch_allocator_io_req_1_0_valid),
    .io_req_1_0_bits_vc_sel_0_0(switch_allocator_io_req_1_0_bits_vc_sel_0_0),
    .io_req_1_0_bits_tail(switch_allocator_io_req_1_0_bits_tail),
    .io_req_0_0_ready(switch_allocator_io_req_0_0_ready),
    .io_req_0_0_valid(switch_allocator_io_req_0_0_valid),
    .io_req_0_0_bits_vc_sel_0_0(switch_allocator_io_req_0_0_bits_vc_sel_0_0),
    .io_req_0_0_bits_tail(switch_allocator_io_req_0_0_bits_tail),
    .io_credit_alloc_0_0_alloc(switch_allocator_io_credit_alloc_0_0_alloc),
    .io_credit_alloc_0_0_tail(switch_allocator_io_credit_alloc_0_0_tail),
    .io_switch_sel_0_0_1_0(switch_allocator_io_switch_sel_0_0_1_0),
    .io_switch_sel_0_0_0_0(switch_allocator_io_switch_sel_0_0_0_0)
  );
  RotatingSingleVCAllocator_1 vc_allocator ( // @[Router.scala 131:30]
    .clock(vc_allocator_clock),
    .reset(vc_allocator_reset),
    .io_req_1_ready(vc_allocator_io_req_1_ready),
    .io_req_1_valid(vc_allocator_io_req_1_valid),
    .io_req_1_bits_vc_sel_0_0(vc_allocator_io_req_1_bits_vc_sel_0_0),
    .io_req_0_ready(vc_allocator_io_req_0_ready),
    .io_req_0_valid(vc_allocator_io_req_0_valid),
    .io_req_0_bits_vc_sel_0_0(vc_allocator_io_req_0_bits_vc_sel_0_0),
    .io_resp_1_vc_sel_0_0(vc_allocator_io_resp_1_vc_sel_0_0),
    .io_resp_0_vc_sel_0_0(vc_allocator_io_resp_0_vc_sel_0_0),
    .io_channel_status_0_0_occupied(vc_allocator_io_channel_status_0_0_occupied),
    .io_out_allocs_0_0_alloc(vc_allocator_io_out_allocs_0_0_alloc)
  );
  RouteComputer_1 route_computer ( // @[Router.scala 134:32]
    .clock(route_computer_clock),
    .reset(route_computer_reset),
    .io_req_1_valid(route_computer_io_req_1_valid),
    .io_req_0_valid(route_computer_io_req_0_valid)
  );
  plusarg_reader #(.FORMAT("noc_util_sample_rate=%d"), .DEFAULT(0), .WIDTH(20)) plusarg_reader ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_out)
  );
  assign auto_debug_out_va_stall_0 = input_unit_0_from_0_io_debug_va_stall; // @[Nodes.scala 1212:84 Router.scala 190:92]
  assign auto_debug_out_va_stall_1 = input_unit_1_from_2_io_debug_va_stall; // @[Nodes.scala 1212:84 Router.scala 190:92]
  assign auto_debug_out_sa_stall_0 = input_unit_0_from_0_io_debug_sa_stall; // @[Nodes.scala 1212:84 Router.scala 191:92]
  assign auto_debug_out_sa_stall_1 = input_unit_1_from_2_io_debug_sa_stall; // @[Nodes.scala 1212:84 Router.scala 191:92]
  assign auto_egress_nodes_out_flit_valid = egress_unit_0_to_1_io_out_valid; // @[Nodes.scala 1212:84 Router.scala 144:65]
  assign auto_egress_nodes_out_flit_bits_head = egress_unit_0_to_1_io_out_bits_head; // @[Nodes.scala 1212:84 Router.scala 144:65]
  assign auto_egress_nodes_out_flit_bits_tail = egress_unit_0_to_1_io_out_bits_tail; // @[Nodes.scala 1212:84 Router.scala 144:65]
  assign auto_egress_nodes_out_flit_bits_payload = egress_unit_0_to_1_io_out_bits_payload; // @[Nodes.scala 1212:84 Router.scala 144:65]
  assign auto_egress_nodes_out_flit_bits_ingress_id = egress_unit_0_to_1_io_out_bits_ingress_id; // @[Nodes.scala 1212:84 Router.scala 144:65]
  assign auto_dest_nodes_in_1_credit_return = input_unit_1_from_2_io_in_credit_return; // @[Nodes.scala 1215:84 Router.scala 141:68]
  assign auto_dest_nodes_in_1_vc_free = input_unit_1_from_2_io_in_vc_free; // @[Nodes.scala 1215:84 Router.scala 141:68]
  assign auto_dest_nodes_in_0_credit_return = input_unit_0_from_0_io_in_credit_return; // @[Nodes.scala 1215:84 Router.scala 141:68]
  assign auto_dest_nodes_in_0_vc_free = input_unit_0_from_0_io_in_vc_free; // @[Nodes.scala 1215:84 Router.scala 141:68]
  assign monitor_clock = clock;
  assign monitor_reset = reset;
  assign monitor_io_in_flit_0_valid = auto_dest_nodes_in_0_flit_0_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_io_in_flit_0_bits_head = auto_dest_nodes_in_0_flit_0_bits_head; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_io_in_flit_0_bits_tail = auto_dest_nodes_in_0_flit_0_bits_tail; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_io_in_flit_0_bits_flow_ingress_node = auto_dest_nodes_in_0_flit_0_bits_flow_ingress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_io_in_flit_0_bits_flow_egress_node = auto_dest_nodes_in_0_flit_0_bits_flow_egress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_io_in_flit_0_bits_virt_channel_id = auto_dest_nodes_in_0_flit_0_bits_virt_channel_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_1_clock = clock;
  assign monitor_1_reset = reset;
  assign monitor_1_io_in_flit_0_valid = auto_dest_nodes_in_1_flit_0_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_1_io_in_flit_0_bits_head = auto_dest_nodes_in_1_flit_0_bits_head; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_1_io_in_flit_0_bits_tail = auto_dest_nodes_in_1_flit_0_bits_tail; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_1_io_in_flit_0_bits_flow_ingress_node = auto_dest_nodes_in_1_flit_0_bits_flow_ingress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_1_io_in_flit_0_bits_flow_egress_node = auto_dest_nodes_in_1_flit_0_bits_flow_egress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign monitor_1_io_in_flit_0_bits_virt_channel_id = auto_dest_nodes_in_1_flit_0_bits_virt_channel_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_0_clock = clock;
  assign input_unit_0_from_0_reset = reset;
  assign input_unit_0_from_0_io_vcalloc_req_ready = vc_allocator_io_req_0_ready; // @[Router.scala 151:23]
  assign input_unit_0_from_0_io_vcalloc_resp_vc_sel_0_0 = vc_allocator_io_resp_0_vc_sel_0_0; // @[Router.scala 153:39]
  assign input_unit_0_from_0_io_out_credit_available_0_0 = egress_unit_0_to_1_io_credit_available_0; // @[Router.scala 162:42]
  assign input_unit_0_from_0_io_salloc_req_0_ready = switch_allocator_io_req_0_0_ready; // @[Router.scala 165:23]
  assign input_unit_0_from_0_io_in_flit_0_valid = auto_dest_nodes_in_0_flit_0_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_0_io_in_flit_0_bits_head = auto_dest_nodes_in_0_flit_0_bits_head; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_0_io_in_flit_0_bits_tail = auto_dest_nodes_in_0_flit_0_bits_tail; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_0_io_in_flit_0_bits_payload = auto_dest_nodes_in_0_flit_0_bits_payload; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_0_io_in_flit_0_bits_flow_ingress_node = auto_dest_nodes_in_0_flit_0_bits_flow_ingress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_0_io_in_flit_0_bits_flow_egress_node = auto_dest_nodes_in_0_flit_0_bits_flow_egress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_0_from_0_io_in_flit_0_bits_virt_channel_id = auto_dest_nodes_in_0_flit_0_bits_virt_channel_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_1_from_2_clock = clock;
  assign input_unit_1_from_2_reset = reset;
  assign input_unit_1_from_2_io_vcalloc_req_ready = vc_allocator_io_req_1_ready; // @[Router.scala 151:23]
  assign input_unit_1_from_2_io_vcalloc_resp_vc_sel_0_0 = vc_allocator_io_resp_1_vc_sel_0_0; // @[Router.scala 153:39]
  assign input_unit_1_from_2_io_out_credit_available_0_0 = egress_unit_0_to_1_io_credit_available_0; // @[Router.scala 162:42]
  assign input_unit_1_from_2_io_salloc_req_0_ready = switch_allocator_io_req_1_0_ready; // @[Router.scala 165:23]
  assign input_unit_1_from_2_io_in_flit_0_valid = auto_dest_nodes_in_1_flit_0_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_1_from_2_io_in_flit_0_bits_head = auto_dest_nodes_in_1_flit_0_bits_head; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_1_from_2_io_in_flit_0_bits_tail = auto_dest_nodes_in_1_flit_0_bits_tail; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_1_from_2_io_in_flit_0_bits_payload = auto_dest_nodes_in_1_flit_0_bits_payload; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_1_from_2_io_in_flit_0_bits_flow_ingress_node = auto_dest_nodes_in_1_flit_0_bits_flow_ingress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_1_from_2_io_in_flit_0_bits_flow_egress_node = auto_dest_nodes_in_1_flit_0_bits_flow_egress_node; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign input_unit_1_from_2_io_in_flit_0_bits_virt_channel_id = auto_dest_nodes_in_1_flit_0_bits_virt_channel_id; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign egress_unit_0_to_1_clock = clock;
  assign egress_unit_0_to_1_reset = reset;
  assign egress_unit_0_to_1_io_in_0_valid = switch_io_out_0_0_valid; // @[Router.scala 172:29]
  assign egress_unit_0_to_1_io_in_0_bits_head = switch_io_out_0_0_bits_head; // @[Router.scala 172:29]
  assign egress_unit_0_to_1_io_in_0_bits_tail = switch_io_out_0_0_bits_tail; // @[Router.scala 172:29]
  assign egress_unit_0_to_1_io_in_0_bits_payload = switch_io_out_0_0_bits_payload; // @[Router.scala 172:29]
  assign egress_unit_0_to_1_io_in_0_bits_flow_ingress_node = switch_io_out_0_0_bits_flow_ingress_node; // @[Router.scala 172:29]
  assign egress_unit_0_to_1_io_allocs_0_alloc = vc_allocator_io_out_allocs_0_0_alloc; // @[Router.scala 157:33]
  assign egress_unit_0_to_1_io_credit_alloc_0_alloc = switch_allocator_io_credit_alloc_0_0_alloc; // @[Router.scala 167:39]
  assign egress_unit_0_to_1_io_credit_alloc_0_tail = switch_allocator_io_credit_alloc_0_0_tail; // @[Router.scala 167:39]
  assign switch_clock = clock;
  assign switch_reset = reset;
  assign switch_io_in_1_0_valid = input_unit_1_from_2_io_out_0_valid; // @[Router.scala 170:23]
  assign switch_io_in_1_0_bits_flit_head = input_unit_1_from_2_io_out_0_bits_flit_head; // @[Router.scala 170:23]
  assign switch_io_in_1_0_bits_flit_tail = input_unit_1_from_2_io_out_0_bits_flit_tail; // @[Router.scala 170:23]
  assign switch_io_in_1_0_bits_flit_payload = input_unit_1_from_2_io_out_0_bits_flit_payload; // @[Router.scala 170:23]
  assign switch_io_in_1_0_bits_flit_flow_ingress_node = input_unit_1_from_2_io_out_0_bits_flit_flow_ingress_node; // @[Router.scala 170:23]
  assign switch_io_in_0_0_valid = input_unit_0_from_0_io_out_0_valid; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_head = input_unit_0_from_0_io_out_0_bits_flit_head; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_tail = input_unit_0_from_0_io_out_0_bits_flit_tail; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_payload = input_unit_0_from_0_io_out_0_bits_flit_payload; // @[Router.scala 170:23]
  assign switch_io_in_0_0_bits_flit_flow_ingress_node = input_unit_0_from_0_io_out_0_bits_flit_flow_ingress_node; // @[Router.scala 170:23]
  assign switch_io_sel_0_0_1_0 = switch_io_sel_REG_0_0_1_0; // @[Router.scala 173:19]
  assign switch_io_sel_0_0_0_0 = switch_io_sel_REG_0_0_0_0; // @[Router.scala 173:19]
  assign switch_allocator_clock = clock;
  assign switch_allocator_reset = reset;
  assign switch_allocator_io_req_1_0_valid = input_unit_1_from_2_io_salloc_req_0_valid; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_vc_sel_0_0 = input_unit_1_from_2_io_salloc_req_0_bits_vc_sel_0_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_1_0_bits_tail = input_unit_1_from_2_io_salloc_req_0_bits_tail; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_valid = input_unit_0_from_0_io_salloc_req_0_valid; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_vc_sel_0_0 = input_unit_0_from_0_io_salloc_req_0_bits_vc_sel_0_0; // @[Router.scala 165:23]
  assign switch_allocator_io_req_0_0_bits_tail = input_unit_0_from_0_io_salloc_req_0_bits_tail; // @[Router.scala 165:23]
  assign vc_allocator_clock = clock;
  assign vc_allocator_reset = reset;
  assign vc_allocator_io_req_1_valid = input_unit_1_from_2_io_vcalloc_req_valid; // @[Router.scala 151:23]
  assign vc_allocator_io_req_1_bits_vc_sel_0_0 = input_unit_1_from_2_io_vcalloc_req_bits_vc_sel_0_0; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_valid = input_unit_0_from_0_io_vcalloc_req_valid; // @[Router.scala 151:23]
  assign vc_allocator_io_req_0_bits_vc_sel_0_0 = input_unit_0_from_0_io_vcalloc_req_bits_vc_sel_0_0; // @[Router.scala 151:23]
  assign vc_allocator_io_channel_status_0_0_occupied = egress_unit_0_to_1_io_channel_status_0_occupied; // @[Router.scala 159:23]
  assign route_computer_clock = clock;
  assign route_computer_reset = reset;
  assign route_computer_io_req_1_valid = input_unit_1_from_2_io_router_req_valid; // @[Router.scala 146:23]
  assign route_computer_io_req_0_valid = input_unit_0_from_0_io_router_req_valid; // @[Router.scala 146:23]
  always @(posedge clock) begin
    switch_io_sel_REG_0_0_1_0 <= switch_allocator_io_switch_sel_0_0_1_0; // @[Router.scala 176:14]
    switch_io_sel_REG_0_0_0_0 <= switch_allocator_io_switch_sel_0_0_0_0; // @[Router.scala 176:14]
    if (reset) begin // @[Router.scala 193:28]
      debug_tsc <= 64'h0; // @[Router.scala 193:28]
    end else begin
      debug_tsc <= _debug_tsc_T_1; // @[Router.scala 194:15]
    end
    if (reset) begin // @[Router.scala 195:31]
      debug_sample <= 64'h0; // @[Router.scala 195:31]
    end else if (debug_sample == _GEN_4) begin // @[Router.scala 198:47]
      debug_sample <= 64'h0; // @[Router.scala 198:62]
    end else begin
      debug_sample <= _debug_sample_T_1; // @[Router.scala 196:18]
    end
    if (reset) begin // @[Router.scala 201:29]
      util_ctr <= 64'h0; // @[Router.scala 201:29]
    end else begin
      util_ctr <= _util_ctr_T_1; // @[Router.scala 203:16]
    end
    if (reset) begin // @[Router.scala 202:26]
      fired <= 1'h0; // @[Router.scala 202:26]
    end else if (plusarg_reader_out != 20'h0 & _T_2 & fired) begin // @[Router.scala 205:81]
      fired <= auto_dest_nodes_in_0_flit_0_valid; // @[Router.scala 208:15]
    end else begin
      fired <= fired | auto_dest_nodes_in_0_flit_0_valid; // @[Router.scala 204:13]
    end
    if (reset) begin // @[Router.scala 201:29]
      util_ctr_1 <= 64'h0; // @[Router.scala 201:29]
    end else begin
      util_ctr_1 <= _util_ctr_T_3; // @[Router.scala 203:16]
    end
    if (reset) begin // @[Router.scala 202:26]
      fired_1 <= 1'h0; // @[Router.scala 202:26]
    end else if (plusarg_reader_out != 20'h0 & _T_2 & fired_1) begin // @[Router.scala 205:81]
      fired_1 <= auto_dest_nodes_in_1_flit_0_valid; // @[Router.scala 208:15]
    end else begin
      fired_1 <= fired_1 | auto_dest_nodes_in_1_flit_0_valid; // @[Router.scala 204:13]
    end
    if (reset) begin // @[Router.scala 201:29]
      util_ctr_2 <= 64'h0; // @[Router.scala 201:29]
    end else begin
      util_ctr_2 <= _util_ctr_T_5; // @[Router.scala 203:16]
    end
    if (reset) begin // @[Router.scala 202:26]
      fired_2 <= 1'h0; // @[Router.scala 202:26]
    end else if (plusarg_reader_out != 20'h0 & _T_2 & fired_2) begin // @[Router.scala 205:81]
      fired_2 <= x1_flit_valid; // @[Router.scala 208:15]
    end else begin
      fired_2 <= fired_2 | x1_flit_valid; // @[Router.scala 204:13]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8 & ~reset) begin
          $fwrite(32'h80000002,"nocsample %d 0 3 %d\n",debug_tsc,util_ctr); // @[Router.scala 207:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_16 & ~reset) begin
          $fwrite(32'h80000002,"nocsample %d 2 3 %d\n",debug_tsc,util_ctr_1); // @[Router.scala 207:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_25 & ~reset) begin
          $fwrite(32'h80000002,"nocsample %d 3 e1 %d\n",debug_tsc,util_ctr_2); // @[Router.scala 207:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  switch_io_sel_REG_0_0_1_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  switch_io_sel_REG_0_0_0_0 = _RAND_1[0:0];
  _RAND_2 = {2{`RANDOM}};
  debug_tsc = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  debug_sample = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  util_ctr = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  fired = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  util_ctr_1 = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  fired_1 = _RAND_7[0:0];
  _RAND_8 = {2{`RANDOM}};
  util_ctr_2 = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  fired_2 = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ClockSinkDomain_3(
  output [1:0]  auto_routers_debug_out_va_stall_0,
  output [1:0]  auto_routers_debug_out_va_stall_1,
  output [1:0]  auto_routers_debug_out_sa_stall_0,
  output [1:0]  auto_routers_debug_out_sa_stall_1,
  output        auto_routers_egress_nodes_out_flit_valid,
  output        auto_routers_egress_nodes_out_flit_bits_head,
  output        auto_routers_egress_nodes_out_flit_bits_tail,
  output [63:0] auto_routers_egress_nodes_out_flit_bits_payload,
  output        auto_routers_egress_nodes_out_flit_bits_ingress_id,
  input         auto_routers_dest_nodes_in_1_flit_0_valid,
  input         auto_routers_dest_nodes_in_1_flit_0_bits_head,
  input         auto_routers_dest_nodes_in_1_flit_0_bits_tail,
  input  [63:0] auto_routers_dest_nodes_in_1_flit_0_bits_payload,
  input  [1:0]  auto_routers_dest_nodes_in_1_flit_0_bits_flow_ingress_node,
  input  [1:0]  auto_routers_dest_nodes_in_1_flit_0_bits_flow_egress_node,
  input  [1:0]  auto_routers_dest_nodes_in_1_flit_0_bits_virt_channel_id,
  output [3:0]  auto_routers_dest_nodes_in_1_credit_return,
  output [3:0]  auto_routers_dest_nodes_in_1_vc_free,
  input         auto_routers_dest_nodes_in_0_flit_0_valid,
  input         auto_routers_dest_nodes_in_0_flit_0_bits_head,
  input         auto_routers_dest_nodes_in_0_flit_0_bits_tail,
  input  [63:0] auto_routers_dest_nodes_in_0_flit_0_bits_payload,
  input  [1:0]  auto_routers_dest_nodes_in_0_flit_0_bits_flow_ingress_node,
  input  [1:0]  auto_routers_dest_nodes_in_0_flit_0_bits_flow_egress_node,
  input  [1:0]  auto_routers_dest_nodes_in_0_flit_0_bits_virt_channel_id,
  output [3:0]  auto_routers_dest_nodes_in_0_credit_return,
  output [3:0]  auto_routers_dest_nodes_in_0_vc_free,
  input         auto_clock_in_clock,
  input         auto_clock_in_reset
);
  wire  routers_clock; // @[NoC.scala 64:22]
  wire  routers_reset; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_debug_out_va_stall_0; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_debug_out_va_stall_1; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_debug_out_sa_stall_0; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_debug_out_sa_stall_1; // @[NoC.scala 64:22]
  wire  routers_auto_egress_nodes_out_flit_valid; // @[NoC.scala 64:22]
  wire  routers_auto_egress_nodes_out_flit_bits_head; // @[NoC.scala 64:22]
  wire  routers_auto_egress_nodes_out_flit_bits_tail; // @[NoC.scala 64:22]
  wire [63:0] routers_auto_egress_nodes_out_flit_bits_payload; // @[NoC.scala 64:22]
  wire  routers_auto_egress_nodes_out_flit_bits_ingress_id; // @[NoC.scala 64:22]
  wire  routers_auto_dest_nodes_in_1_flit_0_valid; // @[NoC.scala 64:22]
  wire  routers_auto_dest_nodes_in_1_flit_0_bits_head; // @[NoC.scala 64:22]
  wire  routers_auto_dest_nodes_in_1_flit_0_bits_tail; // @[NoC.scala 64:22]
  wire [63:0] routers_auto_dest_nodes_in_1_flit_0_bits_payload; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_dest_nodes_in_1_flit_0_bits_flow_ingress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_dest_nodes_in_1_flit_0_bits_flow_egress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_dest_nodes_in_1_flit_0_bits_virt_channel_id; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_dest_nodes_in_1_credit_return; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_dest_nodes_in_1_vc_free; // @[NoC.scala 64:22]
  wire  routers_auto_dest_nodes_in_0_flit_0_valid; // @[NoC.scala 64:22]
  wire  routers_auto_dest_nodes_in_0_flit_0_bits_head; // @[NoC.scala 64:22]
  wire  routers_auto_dest_nodes_in_0_flit_0_bits_tail; // @[NoC.scala 64:22]
  wire [63:0] routers_auto_dest_nodes_in_0_flit_0_bits_payload; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_dest_nodes_in_0_flit_0_bits_flow_ingress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_dest_nodes_in_0_flit_0_bits_flow_egress_node; // @[NoC.scala 64:22]
  wire [1:0] routers_auto_dest_nodes_in_0_flit_0_bits_virt_channel_id; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_dest_nodes_in_0_credit_return; // @[NoC.scala 64:22]
  wire [3:0] routers_auto_dest_nodes_in_0_vc_free; // @[NoC.scala 64:22]
  Router_3 routers ( // @[NoC.scala 64:22]
    .clock(routers_clock),
    .reset(routers_reset),
    .auto_debug_out_va_stall_0(routers_auto_debug_out_va_stall_0),
    .auto_debug_out_va_stall_1(routers_auto_debug_out_va_stall_1),
    .auto_debug_out_sa_stall_0(routers_auto_debug_out_sa_stall_0),
    .auto_debug_out_sa_stall_1(routers_auto_debug_out_sa_stall_1),
    .auto_egress_nodes_out_flit_valid(routers_auto_egress_nodes_out_flit_valid),
    .auto_egress_nodes_out_flit_bits_head(routers_auto_egress_nodes_out_flit_bits_head),
    .auto_egress_nodes_out_flit_bits_tail(routers_auto_egress_nodes_out_flit_bits_tail),
    .auto_egress_nodes_out_flit_bits_payload(routers_auto_egress_nodes_out_flit_bits_payload),
    .auto_egress_nodes_out_flit_bits_ingress_id(routers_auto_egress_nodes_out_flit_bits_ingress_id),
    .auto_dest_nodes_in_1_flit_0_valid(routers_auto_dest_nodes_in_1_flit_0_valid),
    .auto_dest_nodes_in_1_flit_0_bits_head(routers_auto_dest_nodes_in_1_flit_0_bits_head),
    .auto_dest_nodes_in_1_flit_0_bits_tail(routers_auto_dest_nodes_in_1_flit_0_bits_tail),
    .auto_dest_nodes_in_1_flit_0_bits_payload(routers_auto_dest_nodes_in_1_flit_0_bits_payload),
    .auto_dest_nodes_in_1_flit_0_bits_flow_ingress_node(routers_auto_dest_nodes_in_1_flit_0_bits_flow_ingress_node),
    .auto_dest_nodes_in_1_flit_0_bits_flow_egress_node(routers_auto_dest_nodes_in_1_flit_0_bits_flow_egress_node),
    .auto_dest_nodes_in_1_flit_0_bits_virt_channel_id(routers_auto_dest_nodes_in_1_flit_0_bits_virt_channel_id),
    .auto_dest_nodes_in_1_credit_return(routers_auto_dest_nodes_in_1_credit_return),
    .auto_dest_nodes_in_1_vc_free(routers_auto_dest_nodes_in_1_vc_free),
    .auto_dest_nodes_in_0_flit_0_valid(routers_auto_dest_nodes_in_0_flit_0_valid),
    .auto_dest_nodes_in_0_flit_0_bits_head(routers_auto_dest_nodes_in_0_flit_0_bits_head),
    .auto_dest_nodes_in_0_flit_0_bits_tail(routers_auto_dest_nodes_in_0_flit_0_bits_tail),
    .auto_dest_nodes_in_0_flit_0_bits_payload(routers_auto_dest_nodes_in_0_flit_0_bits_payload),
    .auto_dest_nodes_in_0_flit_0_bits_flow_ingress_node(routers_auto_dest_nodes_in_0_flit_0_bits_flow_ingress_node),
    .auto_dest_nodes_in_0_flit_0_bits_flow_egress_node(routers_auto_dest_nodes_in_0_flit_0_bits_flow_egress_node),
    .auto_dest_nodes_in_0_flit_0_bits_virt_channel_id(routers_auto_dest_nodes_in_0_flit_0_bits_virt_channel_id),
    .auto_dest_nodes_in_0_credit_return(routers_auto_dest_nodes_in_0_credit_return),
    .auto_dest_nodes_in_0_vc_free(routers_auto_dest_nodes_in_0_vc_free)
  );
  assign auto_routers_debug_out_va_stall_0 = routers_auto_debug_out_va_stall_0; // @[LazyModule.scala 368:12]
  assign auto_routers_debug_out_va_stall_1 = routers_auto_debug_out_va_stall_1; // @[LazyModule.scala 368:12]
  assign auto_routers_debug_out_sa_stall_0 = routers_auto_debug_out_sa_stall_0; // @[LazyModule.scala 368:12]
  assign auto_routers_debug_out_sa_stall_1 = routers_auto_debug_out_sa_stall_1; // @[LazyModule.scala 368:12]
  assign auto_routers_egress_nodes_out_flit_valid = routers_auto_egress_nodes_out_flit_valid; // @[LazyModule.scala 368:12]
  assign auto_routers_egress_nodes_out_flit_bits_head = routers_auto_egress_nodes_out_flit_bits_head; // @[LazyModule.scala 368:12]
  assign auto_routers_egress_nodes_out_flit_bits_tail = routers_auto_egress_nodes_out_flit_bits_tail; // @[LazyModule.scala 368:12]
  assign auto_routers_egress_nodes_out_flit_bits_payload = routers_auto_egress_nodes_out_flit_bits_payload; // @[LazyModule.scala 368:12]
  assign auto_routers_egress_nodes_out_flit_bits_ingress_id = routers_auto_egress_nodes_out_flit_bits_ingress_id; // @[LazyModule.scala 368:12]
  assign auto_routers_dest_nodes_in_1_credit_return = routers_auto_dest_nodes_in_1_credit_return; // @[LazyModule.scala 366:16]
  assign auto_routers_dest_nodes_in_1_vc_free = routers_auto_dest_nodes_in_1_vc_free; // @[LazyModule.scala 366:16]
  assign auto_routers_dest_nodes_in_0_credit_return = routers_auto_dest_nodes_in_0_credit_return; // @[LazyModule.scala 366:16]
  assign auto_routers_dest_nodes_in_0_vc_free = routers_auto_dest_nodes_in_0_vc_free; // @[LazyModule.scala 366:16]
  assign routers_clock = auto_clock_in_clock; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign routers_reset = auto_clock_in_reset; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_1_flit_0_valid = auto_routers_dest_nodes_in_1_flit_0_valid; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_1_flit_0_bits_head = auto_routers_dest_nodes_in_1_flit_0_bits_head; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_1_flit_0_bits_tail = auto_routers_dest_nodes_in_1_flit_0_bits_tail; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_1_flit_0_bits_payload = auto_routers_dest_nodes_in_1_flit_0_bits_payload; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_1_flit_0_bits_flow_ingress_node =
    auto_routers_dest_nodes_in_1_flit_0_bits_flow_ingress_node; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_1_flit_0_bits_flow_egress_node =
    auto_routers_dest_nodes_in_1_flit_0_bits_flow_egress_node; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_1_flit_0_bits_virt_channel_id =
    auto_routers_dest_nodes_in_1_flit_0_bits_virt_channel_id; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_0_flit_0_valid = auto_routers_dest_nodes_in_0_flit_0_valid; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_0_flit_0_bits_head = auto_routers_dest_nodes_in_0_flit_0_bits_head; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_0_flit_0_bits_tail = auto_routers_dest_nodes_in_0_flit_0_bits_tail; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_0_flit_0_bits_payload = auto_routers_dest_nodes_in_0_flit_0_bits_payload; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_0_flit_0_bits_flow_ingress_node =
    auto_routers_dest_nodes_in_0_flit_0_bits_flow_ingress_node; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_0_flit_0_bits_flow_egress_node =
    auto_routers_dest_nodes_in_0_flit_0_bits_flow_egress_node; // @[LazyModule.scala 366:16]
  assign routers_auto_dest_nodes_in_0_flit_0_bits_virt_channel_id =
    auto_routers_dest_nodes_in_0_flit_0_bits_virt_channel_id; // @[LazyModule.scala 366:16]
endmodule
module NoC(
  input         clock,
  input         reset,
  output        io_ingress_1_flit_ready,
  input         io_ingress_1_flit_valid,
  input         io_ingress_1_flit_bits_head,
  input         io_ingress_1_flit_bits_tail,
  input  [63:0] io_ingress_1_flit_bits_payload,
  input         io_ingress_1_flit_bits_egress_id,
  output        io_ingress_0_flit_ready,
  input         io_ingress_0_flit_valid,
  input         io_ingress_0_flit_bits_head,
  input         io_ingress_0_flit_bits_tail,
  input  [63:0] io_ingress_0_flit_bits_payload,
  input         io_ingress_0_flit_bits_egress_id,
  output        io_egress_1_flit_valid,
  output        io_egress_1_flit_bits_head,
  output        io_egress_1_flit_bits_tail,
  output [63:0] io_egress_1_flit_bits_payload,
  output        io_egress_1_flit_bits_ingress_id,
  output        io_egress_0_flit_valid,
  output        io_egress_0_flit_bits_head,
  output        io_egress_0_flit_bits_tail,
  output [63:0] io_egress_0_flit_bits_payload,
  output        io_egress_0_flit_bits_ingress_id,
  input         io_router_clocks_0_clock,
  input         io_router_clocks_0_reset,
  input         io_router_clocks_1_clock,
  input         io_router_clocks_1_reset,
  input         io_router_clocks_2_clock,
  input         io_router_clocks_2_reset,
  input         io_router_clocks_3_clock,
  input         io_router_clocks_3_reset
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  router_sink_domain_auto_routers_ingress_nodes_in_flit_ready; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_routers_ingress_nodes_in_flit_valid; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_routers_ingress_nodes_in_flit_bits_head; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_routers_ingress_nodes_in_flit_bits_tail; // @[NoC.scala 38:40]
  wire [63:0] router_sink_domain_auto_routers_ingress_nodes_in_flit_bits_payload; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_routers_ingress_nodes_in_flit_bits_egress_id; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_routers_source_nodes_out_1_flit_0_valid; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_routers_source_nodes_out_1_flit_0_bits_head; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_routers_source_nodes_out_1_flit_0_bits_tail; // @[NoC.scala 38:40]
  wire [63:0] router_sink_domain_auto_routers_source_nodes_out_1_flit_0_bits_payload; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_auto_routers_source_nodes_out_1_flit_0_bits_flow_ingress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_auto_routers_source_nodes_out_1_flit_0_bits_flow_egress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_auto_routers_source_nodes_out_1_flit_0_bits_virt_channel_id; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_auto_routers_source_nodes_out_1_credit_return; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_auto_routers_source_nodes_out_1_vc_free; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_routers_source_nodes_out_0_flit_0_valid; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_routers_source_nodes_out_0_flit_0_bits_head; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_routers_source_nodes_out_0_flit_0_bits_tail; // @[NoC.scala 38:40]
  wire [63:0] router_sink_domain_auto_routers_source_nodes_out_0_flit_0_bits_payload; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_auto_routers_source_nodes_out_0_flit_0_bits_flow_ingress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_auto_routers_source_nodes_out_0_flit_0_bits_flow_egress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_auto_routers_source_nodes_out_0_flit_0_bits_virt_channel_id; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_auto_routers_source_nodes_out_0_credit_return; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_auto_routers_source_nodes_out_0_vc_free; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_clock_in_clock; // @[NoC.scala 38:40]
  wire  router_sink_domain_auto_clock_in_reset; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_1_auto_routers_debug_out_va_stall_0; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_1_auto_routers_debug_out_va_stall_1; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_1_auto_routers_debug_out_sa_stall_0; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_1_auto_routers_debug_out_sa_stall_1; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_routers_egress_nodes_out_flit_valid; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_routers_egress_nodes_out_flit_bits_head; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_routers_egress_nodes_out_flit_bits_tail; // @[NoC.scala 38:40]
  wire [63:0] router_sink_domain_1_auto_routers_egress_nodes_out_flit_bits_payload; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_routers_egress_nodes_out_flit_bits_ingress_id; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_routers_dest_nodes_in_1_flit_0_valid; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_routers_dest_nodes_in_1_flit_0_bits_head; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_routers_dest_nodes_in_1_flit_0_bits_tail; // @[NoC.scala 38:40]
  wire [63:0] router_sink_domain_1_auto_routers_dest_nodes_in_1_flit_0_bits_payload; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_1_auto_routers_dest_nodes_in_1_flit_0_bits_flow_ingress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_1_auto_routers_dest_nodes_in_1_flit_0_bits_flow_egress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_1_auto_routers_dest_nodes_in_1_flit_0_bits_virt_channel_id; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_1_auto_routers_dest_nodes_in_1_credit_return; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_1_auto_routers_dest_nodes_in_1_vc_free; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_routers_dest_nodes_in_0_flit_0_valid; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_routers_dest_nodes_in_0_flit_0_bits_head; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_routers_dest_nodes_in_0_flit_0_bits_tail; // @[NoC.scala 38:40]
  wire [63:0] router_sink_domain_1_auto_routers_dest_nodes_in_0_flit_0_bits_payload; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_1_auto_routers_dest_nodes_in_0_flit_0_bits_flow_ingress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_1_auto_routers_dest_nodes_in_0_flit_0_bits_flow_egress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_1_auto_routers_dest_nodes_in_0_flit_0_bits_virt_channel_id; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_1_auto_routers_dest_nodes_in_0_credit_return; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_1_auto_routers_dest_nodes_in_0_vc_free; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_clock_in_clock; // @[NoC.scala 38:40]
  wire  router_sink_domain_1_auto_clock_in_reset; // @[NoC.scala 38:40]
  wire  router_sink_domain_2_auto_routers_ingress_nodes_in_flit_ready; // @[NoC.scala 38:40]
  wire  router_sink_domain_2_auto_routers_ingress_nodes_in_flit_valid; // @[NoC.scala 38:40]
  wire  router_sink_domain_2_auto_routers_ingress_nodes_in_flit_bits_head; // @[NoC.scala 38:40]
  wire  router_sink_domain_2_auto_routers_ingress_nodes_in_flit_bits_tail; // @[NoC.scala 38:40]
  wire [63:0] router_sink_domain_2_auto_routers_ingress_nodes_in_flit_bits_payload; // @[NoC.scala 38:40]
  wire  router_sink_domain_2_auto_routers_ingress_nodes_in_flit_bits_egress_id; // @[NoC.scala 38:40]
  wire  router_sink_domain_2_auto_routers_source_nodes_out_1_flit_0_valid; // @[NoC.scala 38:40]
  wire  router_sink_domain_2_auto_routers_source_nodes_out_1_flit_0_bits_head; // @[NoC.scala 38:40]
  wire  router_sink_domain_2_auto_routers_source_nodes_out_1_flit_0_bits_tail; // @[NoC.scala 38:40]
  wire [63:0] router_sink_domain_2_auto_routers_source_nodes_out_1_flit_0_bits_payload; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_2_auto_routers_source_nodes_out_1_flit_0_bits_flow_ingress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_2_auto_routers_source_nodes_out_1_flit_0_bits_flow_egress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_2_auto_routers_source_nodes_out_1_flit_0_bits_virt_channel_id; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_2_auto_routers_source_nodes_out_1_credit_return; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_2_auto_routers_source_nodes_out_1_vc_free; // @[NoC.scala 38:40]
  wire  router_sink_domain_2_auto_routers_source_nodes_out_0_flit_0_valid; // @[NoC.scala 38:40]
  wire  router_sink_domain_2_auto_routers_source_nodes_out_0_flit_0_bits_head; // @[NoC.scala 38:40]
  wire  router_sink_domain_2_auto_routers_source_nodes_out_0_flit_0_bits_tail; // @[NoC.scala 38:40]
  wire [63:0] router_sink_domain_2_auto_routers_source_nodes_out_0_flit_0_bits_payload; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_2_auto_routers_source_nodes_out_0_flit_0_bits_flow_ingress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_2_auto_routers_source_nodes_out_0_flit_0_bits_flow_egress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_2_auto_routers_source_nodes_out_0_flit_0_bits_virt_channel_id; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_2_auto_routers_source_nodes_out_0_credit_return; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_2_auto_routers_source_nodes_out_0_vc_free; // @[NoC.scala 38:40]
  wire  router_sink_domain_2_auto_clock_in_clock; // @[NoC.scala 38:40]
  wire  router_sink_domain_2_auto_clock_in_reset; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_3_auto_routers_debug_out_va_stall_0; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_3_auto_routers_debug_out_va_stall_1; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_3_auto_routers_debug_out_sa_stall_0; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_3_auto_routers_debug_out_sa_stall_1; // @[NoC.scala 38:40]
  wire  router_sink_domain_3_auto_routers_egress_nodes_out_flit_valid; // @[NoC.scala 38:40]
  wire  router_sink_domain_3_auto_routers_egress_nodes_out_flit_bits_head; // @[NoC.scala 38:40]
  wire  router_sink_domain_3_auto_routers_egress_nodes_out_flit_bits_tail; // @[NoC.scala 38:40]
  wire [63:0] router_sink_domain_3_auto_routers_egress_nodes_out_flit_bits_payload; // @[NoC.scala 38:40]
  wire  router_sink_domain_3_auto_routers_egress_nodes_out_flit_bits_ingress_id; // @[NoC.scala 38:40]
  wire  router_sink_domain_3_auto_routers_dest_nodes_in_1_flit_0_valid; // @[NoC.scala 38:40]
  wire  router_sink_domain_3_auto_routers_dest_nodes_in_1_flit_0_bits_head; // @[NoC.scala 38:40]
  wire  router_sink_domain_3_auto_routers_dest_nodes_in_1_flit_0_bits_tail; // @[NoC.scala 38:40]
  wire [63:0] router_sink_domain_3_auto_routers_dest_nodes_in_1_flit_0_bits_payload; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_3_auto_routers_dest_nodes_in_1_flit_0_bits_flow_ingress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_3_auto_routers_dest_nodes_in_1_flit_0_bits_flow_egress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_3_auto_routers_dest_nodes_in_1_flit_0_bits_virt_channel_id; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_3_auto_routers_dest_nodes_in_1_credit_return; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_3_auto_routers_dest_nodes_in_1_vc_free; // @[NoC.scala 38:40]
  wire  router_sink_domain_3_auto_routers_dest_nodes_in_0_flit_0_valid; // @[NoC.scala 38:40]
  wire  router_sink_domain_3_auto_routers_dest_nodes_in_0_flit_0_bits_head; // @[NoC.scala 38:40]
  wire  router_sink_domain_3_auto_routers_dest_nodes_in_0_flit_0_bits_tail; // @[NoC.scala 38:40]
  wire [63:0] router_sink_domain_3_auto_routers_dest_nodes_in_0_flit_0_bits_payload; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_3_auto_routers_dest_nodes_in_0_flit_0_bits_flow_ingress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_3_auto_routers_dest_nodes_in_0_flit_0_bits_flow_egress_node; // @[NoC.scala 38:40]
  wire [1:0] router_sink_domain_3_auto_routers_dest_nodes_in_0_flit_0_bits_virt_channel_id; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_3_auto_routers_dest_nodes_in_0_credit_return; // @[NoC.scala 38:40]
  wire [3:0] router_sink_domain_3_auto_routers_dest_nodes_in_0_vc_free; // @[NoC.scala 38:40]
  wire  router_sink_domain_3_auto_clock_in_clock; // @[NoC.scala 38:40]
  wire  router_sink_domain_3_auto_clock_in_reset; // @[NoC.scala 38:40]
  reg [63:0] debug_va_stall_ctr; // @[NoC.scala 160:37]
  reg [63:0] debug_sa_stall_ctr; // @[NoC.scala 161:37]
  wire [63:0] debug_any_stall_ctr = debug_va_stall_ctr + debug_sa_stall_ctr; // @[NoC.scala 162:50]
  wire [1:0] bundleIn_0_3_va_stall_0 = router_sink_domain_1_auto_routers_debug_out_va_stall_0; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  wire [1:0] bundleIn_0_3_va_stall_1 = router_sink_domain_1_auto_routers_debug_out_va_stall_1; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  wire [1:0] _debug_va_stall_ctr_T_1 = bundleIn_0_3_va_stall_0 + bundleIn_0_3_va_stall_1; // @[NoC.scala 163:91]
  wire [1:0] bundleIn_0_5_va_stall_0 = router_sink_domain_3_auto_routers_debug_out_va_stall_0; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  wire [1:0] bundleIn_0_5_va_stall_1 = router_sink_domain_3_auto_routers_debug_out_va_stall_1; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  wire [1:0] _debug_va_stall_ctr_T_3 = bundleIn_0_5_va_stall_0 + bundleIn_0_5_va_stall_1; // @[NoC.scala 163:91]
  wire [2:0] _debug_va_stall_ctr_T_4 = {{1'd0}, _debug_va_stall_ctr_T_1}; // @[NoC.scala 163:104]
  wire [2:0] _debug_va_stall_ctr_T_6 = {{1'd0}, _debug_va_stall_ctr_T_4[1:0]}; // @[NoC.scala 163:104]
  wire [1:0] _debug_va_stall_ctr_T_9 = _debug_va_stall_ctr_T_6[1:0] + _debug_va_stall_ctr_T_3; // @[NoC.scala 163:104]
  wire [63:0] _GEN_0 = {{62'd0}, _debug_va_stall_ctr_T_9}; // @[NoC.scala 163:46]
  wire [63:0] _debug_va_stall_ctr_T_11 = debug_va_stall_ctr + _GEN_0; // @[NoC.scala 163:46]
  wire [1:0] bundleIn_0_3_sa_stall_0 = router_sink_domain_1_auto_routers_debug_out_sa_stall_0; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  wire [1:0] bundleIn_0_3_sa_stall_1 = router_sink_domain_1_auto_routers_debug_out_sa_stall_1; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  wire [1:0] _debug_sa_stall_ctr_T_1 = bundleIn_0_3_sa_stall_0 + bundleIn_0_3_sa_stall_1; // @[NoC.scala 164:91]
  wire [1:0] bundleIn_0_5_sa_stall_0 = router_sink_domain_3_auto_routers_debug_out_sa_stall_0; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  wire [1:0] bundleIn_0_5_sa_stall_1 = router_sink_domain_3_auto_routers_debug_out_sa_stall_1; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  wire [1:0] _debug_sa_stall_ctr_T_3 = bundleIn_0_5_sa_stall_0 + bundleIn_0_5_sa_stall_1; // @[NoC.scala 164:91]
  wire [2:0] _debug_sa_stall_ctr_T_4 = {{1'd0}, _debug_sa_stall_ctr_T_1}; // @[NoC.scala 164:104]
  wire [2:0] _debug_sa_stall_ctr_T_6 = {{1'd0}, _debug_sa_stall_ctr_T_4[1:0]}; // @[NoC.scala 164:104]
  wire [1:0] _debug_sa_stall_ctr_T_9 = _debug_sa_stall_ctr_T_6[1:0] + _debug_sa_stall_ctr_T_3; // @[NoC.scala 164:104]
  wire [63:0] _GEN_1 = {{62'd0}, _debug_sa_stall_ctr_T_9}; // @[NoC.scala 164:46]
  wire [63:0] _debug_sa_stall_ctr_T_11 = debug_sa_stall_ctr + _GEN_1; // @[NoC.scala 164:46]
  ClockSinkDomain router_sink_domain ( // @[NoC.scala 38:40]
    .auto_routers_ingress_nodes_in_flit_ready(router_sink_domain_auto_routers_ingress_nodes_in_flit_ready),
    .auto_routers_ingress_nodes_in_flit_valid(router_sink_domain_auto_routers_ingress_nodes_in_flit_valid),
    .auto_routers_ingress_nodes_in_flit_bits_head(router_sink_domain_auto_routers_ingress_nodes_in_flit_bits_head),
    .auto_routers_ingress_nodes_in_flit_bits_tail(router_sink_domain_auto_routers_ingress_nodes_in_flit_bits_tail),
    .auto_routers_ingress_nodes_in_flit_bits_payload(router_sink_domain_auto_routers_ingress_nodes_in_flit_bits_payload)
      ,
    .auto_routers_ingress_nodes_in_flit_bits_egress_id(
      router_sink_domain_auto_routers_ingress_nodes_in_flit_bits_egress_id),
    .auto_routers_source_nodes_out_1_flit_0_valid(router_sink_domain_auto_routers_source_nodes_out_1_flit_0_valid),
    .auto_routers_source_nodes_out_1_flit_0_bits_head(
      router_sink_domain_auto_routers_source_nodes_out_1_flit_0_bits_head),
    .auto_routers_source_nodes_out_1_flit_0_bits_tail(
      router_sink_domain_auto_routers_source_nodes_out_1_flit_0_bits_tail),
    .auto_routers_source_nodes_out_1_flit_0_bits_payload(
      router_sink_domain_auto_routers_source_nodes_out_1_flit_0_bits_payload),
    .auto_routers_source_nodes_out_1_flit_0_bits_flow_ingress_node(
      router_sink_domain_auto_routers_source_nodes_out_1_flit_0_bits_flow_ingress_node),
    .auto_routers_source_nodes_out_1_flit_0_bits_flow_egress_node(
      router_sink_domain_auto_routers_source_nodes_out_1_flit_0_bits_flow_egress_node),
    .auto_routers_source_nodes_out_1_flit_0_bits_virt_channel_id(
      router_sink_domain_auto_routers_source_nodes_out_1_flit_0_bits_virt_channel_id),
    .auto_routers_source_nodes_out_1_credit_return(router_sink_domain_auto_routers_source_nodes_out_1_credit_return),
    .auto_routers_source_nodes_out_1_vc_free(router_sink_domain_auto_routers_source_nodes_out_1_vc_free),
    .auto_routers_source_nodes_out_0_flit_0_valid(router_sink_domain_auto_routers_source_nodes_out_0_flit_0_valid),
    .auto_routers_source_nodes_out_0_flit_0_bits_head(
      router_sink_domain_auto_routers_source_nodes_out_0_flit_0_bits_head),
    .auto_routers_source_nodes_out_0_flit_0_bits_tail(
      router_sink_domain_auto_routers_source_nodes_out_0_flit_0_bits_tail),
    .auto_routers_source_nodes_out_0_flit_0_bits_payload(
      router_sink_domain_auto_routers_source_nodes_out_0_flit_0_bits_payload),
    .auto_routers_source_nodes_out_0_flit_0_bits_flow_ingress_node(
      router_sink_domain_auto_routers_source_nodes_out_0_flit_0_bits_flow_ingress_node),
    .auto_routers_source_nodes_out_0_flit_0_bits_flow_egress_node(
      router_sink_domain_auto_routers_source_nodes_out_0_flit_0_bits_flow_egress_node),
    .auto_routers_source_nodes_out_0_flit_0_bits_virt_channel_id(
      router_sink_domain_auto_routers_source_nodes_out_0_flit_0_bits_virt_channel_id),
    .auto_routers_source_nodes_out_0_credit_return(router_sink_domain_auto_routers_source_nodes_out_0_credit_return),
    .auto_routers_source_nodes_out_0_vc_free(router_sink_domain_auto_routers_source_nodes_out_0_vc_free),
    .auto_clock_in_clock(router_sink_domain_auto_clock_in_clock),
    .auto_clock_in_reset(router_sink_domain_auto_clock_in_reset)
  );
  ClockSinkDomain_1 router_sink_domain_1 ( // @[NoC.scala 38:40]
    .auto_routers_debug_out_va_stall_0(router_sink_domain_1_auto_routers_debug_out_va_stall_0),
    .auto_routers_debug_out_va_stall_1(router_sink_domain_1_auto_routers_debug_out_va_stall_1),
    .auto_routers_debug_out_sa_stall_0(router_sink_domain_1_auto_routers_debug_out_sa_stall_0),
    .auto_routers_debug_out_sa_stall_1(router_sink_domain_1_auto_routers_debug_out_sa_stall_1),
    .auto_routers_egress_nodes_out_flit_valid(router_sink_domain_1_auto_routers_egress_nodes_out_flit_valid),
    .auto_routers_egress_nodes_out_flit_bits_head(router_sink_domain_1_auto_routers_egress_nodes_out_flit_bits_head),
    .auto_routers_egress_nodes_out_flit_bits_tail(router_sink_domain_1_auto_routers_egress_nodes_out_flit_bits_tail),
    .auto_routers_egress_nodes_out_flit_bits_payload(
      router_sink_domain_1_auto_routers_egress_nodes_out_flit_bits_payload),
    .auto_routers_egress_nodes_out_flit_bits_ingress_id(
      router_sink_domain_1_auto_routers_egress_nodes_out_flit_bits_ingress_id),
    .auto_routers_dest_nodes_in_1_flit_0_valid(router_sink_domain_1_auto_routers_dest_nodes_in_1_flit_0_valid),
    .auto_routers_dest_nodes_in_1_flit_0_bits_head(router_sink_domain_1_auto_routers_dest_nodes_in_1_flit_0_bits_head),
    .auto_routers_dest_nodes_in_1_flit_0_bits_tail(router_sink_domain_1_auto_routers_dest_nodes_in_1_flit_0_bits_tail),
    .auto_routers_dest_nodes_in_1_flit_0_bits_payload(
      router_sink_domain_1_auto_routers_dest_nodes_in_1_flit_0_bits_payload),
    .auto_routers_dest_nodes_in_1_flit_0_bits_flow_ingress_node(
      router_sink_domain_1_auto_routers_dest_nodes_in_1_flit_0_bits_flow_ingress_node),
    .auto_routers_dest_nodes_in_1_flit_0_bits_flow_egress_node(
      router_sink_domain_1_auto_routers_dest_nodes_in_1_flit_0_bits_flow_egress_node),
    .auto_routers_dest_nodes_in_1_flit_0_bits_virt_channel_id(
      router_sink_domain_1_auto_routers_dest_nodes_in_1_flit_0_bits_virt_channel_id),
    .auto_routers_dest_nodes_in_1_credit_return(router_sink_domain_1_auto_routers_dest_nodes_in_1_credit_return),
    .auto_routers_dest_nodes_in_1_vc_free(router_sink_domain_1_auto_routers_dest_nodes_in_1_vc_free),
    .auto_routers_dest_nodes_in_0_flit_0_valid(router_sink_domain_1_auto_routers_dest_nodes_in_0_flit_0_valid),
    .auto_routers_dest_nodes_in_0_flit_0_bits_head(router_sink_domain_1_auto_routers_dest_nodes_in_0_flit_0_bits_head),
    .auto_routers_dest_nodes_in_0_flit_0_bits_tail(router_sink_domain_1_auto_routers_dest_nodes_in_0_flit_0_bits_tail),
    .auto_routers_dest_nodes_in_0_flit_0_bits_payload(
      router_sink_domain_1_auto_routers_dest_nodes_in_0_flit_0_bits_payload),
    .auto_routers_dest_nodes_in_0_flit_0_bits_flow_ingress_node(
      router_sink_domain_1_auto_routers_dest_nodes_in_0_flit_0_bits_flow_ingress_node),
    .auto_routers_dest_nodes_in_0_flit_0_bits_flow_egress_node(
      router_sink_domain_1_auto_routers_dest_nodes_in_0_flit_0_bits_flow_egress_node),
    .auto_routers_dest_nodes_in_0_flit_0_bits_virt_channel_id(
      router_sink_domain_1_auto_routers_dest_nodes_in_0_flit_0_bits_virt_channel_id),
    .auto_routers_dest_nodes_in_0_credit_return(router_sink_domain_1_auto_routers_dest_nodes_in_0_credit_return),
    .auto_routers_dest_nodes_in_0_vc_free(router_sink_domain_1_auto_routers_dest_nodes_in_0_vc_free),
    .auto_clock_in_clock(router_sink_domain_1_auto_clock_in_clock),
    .auto_clock_in_reset(router_sink_domain_1_auto_clock_in_reset)
  );
  ClockSinkDomain_2 router_sink_domain_2 ( // @[NoC.scala 38:40]
    .auto_routers_ingress_nodes_in_flit_ready(router_sink_domain_2_auto_routers_ingress_nodes_in_flit_ready),
    .auto_routers_ingress_nodes_in_flit_valid(router_sink_domain_2_auto_routers_ingress_nodes_in_flit_valid),
    .auto_routers_ingress_nodes_in_flit_bits_head(router_sink_domain_2_auto_routers_ingress_nodes_in_flit_bits_head),
    .auto_routers_ingress_nodes_in_flit_bits_tail(router_sink_domain_2_auto_routers_ingress_nodes_in_flit_bits_tail),
    .auto_routers_ingress_nodes_in_flit_bits_payload(
      router_sink_domain_2_auto_routers_ingress_nodes_in_flit_bits_payload),
    .auto_routers_ingress_nodes_in_flit_bits_egress_id(
      router_sink_domain_2_auto_routers_ingress_nodes_in_flit_bits_egress_id),
    .auto_routers_source_nodes_out_1_flit_0_valid(router_sink_domain_2_auto_routers_source_nodes_out_1_flit_0_valid),
    .auto_routers_source_nodes_out_1_flit_0_bits_head(
      router_sink_domain_2_auto_routers_source_nodes_out_1_flit_0_bits_head),
    .auto_routers_source_nodes_out_1_flit_0_bits_tail(
      router_sink_domain_2_auto_routers_source_nodes_out_1_flit_0_bits_tail),
    .auto_routers_source_nodes_out_1_flit_0_bits_payload(
      router_sink_domain_2_auto_routers_source_nodes_out_1_flit_0_bits_payload),
    .auto_routers_source_nodes_out_1_flit_0_bits_flow_ingress_node(
      router_sink_domain_2_auto_routers_source_nodes_out_1_flit_0_bits_flow_ingress_node),
    .auto_routers_source_nodes_out_1_flit_0_bits_flow_egress_node(
      router_sink_domain_2_auto_routers_source_nodes_out_1_flit_0_bits_flow_egress_node),
    .auto_routers_source_nodes_out_1_flit_0_bits_virt_channel_id(
      router_sink_domain_2_auto_routers_source_nodes_out_1_flit_0_bits_virt_channel_id),
    .auto_routers_source_nodes_out_1_credit_return(router_sink_domain_2_auto_routers_source_nodes_out_1_credit_return),
    .auto_routers_source_nodes_out_1_vc_free(router_sink_domain_2_auto_routers_source_nodes_out_1_vc_free),
    .auto_routers_source_nodes_out_0_flit_0_valid(router_sink_domain_2_auto_routers_source_nodes_out_0_flit_0_valid),
    .auto_routers_source_nodes_out_0_flit_0_bits_head(
      router_sink_domain_2_auto_routers_source_nodes_out_0_flit_0_bits_head),
    .auto_routers_source_nodes_out_0_flit_0_bits_tail(
      router_sink_domain_2_auto_routers_source_nodes_out_0_flit_0_bits_tail),
    .auto_routers_source_nodes_out_0_flit_0_bits_payload(
      router_sink_domain_2_auto_routers_source_nodes_out_0_flit_0_bits_payload),
    .auto_routers_source_nodes_out_0_flit_0_bits_flow_ingress_node(
      router_sink_domain_2_auto_routers_source_nodes_out_0_flit_0_bits_flow_ingress_node),
    .auto_routers_source_nodes_out_0_flit_0_bits_flow_egress_node(
      router_sink_domain_2_auto_routers_source_nodes_out_0_flit_0_bits_flow_egress_node),
    .auto_routers_source_nodes_out_0_flit_0_bits_virt_channel_id(
      router_sink_domain_2_auto_routers_source_nodes_out_0_flit_0_bits_virt_channel_id),
    .auto_routers_source_nodes_out_0_credit_return(router_sink_domain_2_auto_routers_source_nodes_out_0_credit_return),
    .auto_routers_source_nodes_out_0_vc_free(router_sink_domain_2_auto_routers_source_nodes_out_0_vc_free),
    .auto_clock_in_clock(router_sink_domain_2_auto_clock_in_clock),
    .auto_clock_in_reset(router_sink_domain_2_auto_clock_in_reset)
  );
  ClockSinkDomain_3 router_sink_domain_3 ( // @[NoC.scala 38:40]
    .auto_routers_debug_out_va_stall_0(router_sink_domain_3_auto_routers_debug_out_va_stall_0),
    .auto_routers_debug_out_va_stall_1(router_sink_domain_3_auto_routers_debug_out_va_stall_1),
    .auto_routers_debug_out_sa_stall_0(router_sink_domain_3_auto_routers_debug_out_sa_stall_0),
    .auto_routers_debug_out_sa_stall_1(router_sink_domain_3_auto_routers_debug_out_sa_stall_1),
    .auto_routers_egress_nodes_out_flit_valid(router_sink_domain_3_auto_routers_egress_nodes_out_flit_valid),
    .auto_routers_egress_nodes_out_flit_bits_head(router_sink_domain_3_auto_routers_egress_nodes_out_flit_bits_head),
    .auto_routers_egress_nodes_out_flit_bits_tail(router_sink_domain_3_auto_routers_egress_nodes_out_flit_bits_tail),
    .auto_routers_egress_nodes_out_flit_bits_payload(
      router_sink_domain_3_auto_routers_egress_nodes_out_flit_bits_payload),
    .auto_routers_egress_nodes_out_flit_bits_ingress_id(
      router_sink_domain_3_auto_routers_egress_nodes_out_flit_bits_ingress_id),
    .auto_routers_dest_nodes_in_1_flit_0_valid(router_sink_domain_3_auto_routers_dest_nodes_in_1_flit_0_valid),
    .auto_routers_dest_nodes_in_1_flit_0_bits_head(router_sink_domain_3_auto_routers_dest_nodes_in_1_flit_0_bits_head),
    .auto_routers_dest_nodes_in_1_flit_0_bits_tail(router_sink_domain_3_auto_routers_dest_nodes_in_1_flit_0_bits_tail),
    .auto_routers_dest_nodes_in_1_flit_0_bits_payload(
      router_sink_domain_3_auto_routers_dest_nodes_in_1_flit_0_bits_payload),
    .auto_routers_dest_nodes_in_1_flit_0_bits_flow_ingress_node(
      router_sink_domain_3_auto_routers_dest_nodes_in_1_flit_0_bits_flow_ingress_node),
    .auto_routers_dest_nodes_in_1_flit_0_bits_flow_egress_node(
      router_sink_domain_3_auto_routers_dest_nodes_in_1_flit_0_bits_flow_egress_node),
    .auto_routers_dest_nodes_in_1_flit_0_bits_virt_channel_id(
      router_sink_domain_3_auto_routers_dest_nodes_in_1_flit_0_bits_virt_channel_id),
    .auto_routers_dest_nodes_in_1_credit_return(router_sink_domain_3_auto_routers_dest_nodes_in_1_credit_return),
    .auto_routers_dest_nodes_in_1_vc_free(router_sink_domain_3_auto_routers_dest_nodes_in_1_vc_free),
    .auto_routers_dest_nodes_in_0_flit_0_valid(router_sink_domain_3_auto_routers_dest_nodes_in_0_flit_0_valid),
    .auto_routers_dest_nodes_in_0_flit_0_bits_head(router_sink_domain_3_auto_routers_dest_nodes_in_0_flit_0_bits_head),
    .auto_routers_dest_nodes_in_0_flit_0_bits_tail(router_sink_domain_3_auto_routers_dest_nodes_in_0_flit_0_bits_tail),
    .auto_routers_dest_nodes_in_0_flit_0_bits_payload(
      router_sink_domain_3_auto_routers_dest_nodes_in_0_flit_0_bits_payload),
    .auto_routers_dest_nodes_in_0_flit_0_bits_flow_ingress_node(
      router_sink_domain_3_auto_routers_dest_nodes_in_0_flit_0_bits_flow_ingress_node),
    .auto_routers_dest_nodes_in_0_flit_0_bits_flow_egress_node(
      router_sink_domain_3_auto_routers_dest_nodes_in_0_flit_0_bits_flow_egress_node),
    .auto_routers_dest_nodes_in_0_flit_0_bits_virt_channel_id(
      router_sink_domain_3_auto_routers_dest_nodes_in_0_flit_0_bits_virt_channel_id),
    .auto_routers_dest_nodes_in_0_credit_return(router_sink_domain_3_auto_routers_dest_nodes_in_0_credit_return),
    .auto_routers_dest_nodes_in_0_vc_free(router_sink_domain_3_auto_routers_dest_nodes_in_0_vc_free),
    .auto_clock_in_clock(router_sink_domain_3_auto_clock_in_clock),
    .auto_clock_in_reset(router_sink_domain_3_auto_clock_in_reset)
  );
  assign io_ingress_1_flit_ready = router_sink_domain_2_auto_routers_ingress_nodes_in_flit_ready; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign io_ingress_0_flit_ready = router_sink_domain_auto_routers_ingress_nodes_in_flit_ready; // @[Nodes.scala 1212:84 LazyModule.scala 355:16]
  assign io_egress_1_flit_valid = router_sink_domain_3_auto_routers_egress_nodes_out_flit_valid; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign io_egress_1_flit_bits_head = router_sink_domain_3_auto_routers_egress_nodes_out_flit_bits_head; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign io_egress_1_flit_bits_tail = router_sink_domain_3_auto_routers_egress_nodes_out_flit_bits_tail; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign io_egress_1_flit_bits_payload = router_sink_domain_3_auto_routers_egress_nodes_out_flit_bits_payload; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign io_egress_1_flit_bits_ingress_id = router_sink_domain_3_auto_routers_egress_nodes_out_flit_bits_ingress_id; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign io_egress_0_flit_valid = router_sink_domain_1_auto_routers_egress_nodes_out_flit_valid; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign io_egress_0_flit_bits_head = router_sink_domain_1_auto_routers_egress_nodes_out_flit_bits_head; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign io_egress_0_flit_bits_tail = router_sink_domain_1_auto_routers_egress_nodes_out_flit_bits_tail; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign io_egress_0_flit_bits_payload = router_sink_domain_1_auto_routers_egress_nodes_out_flit_bits_payload; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign io_egress_0_flit_bits_ingress_id = router_sink_domain_1_auto_routers_egress_nodes_out_flit_bits_ingress_id; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign router_sink_domain_auto_routers_ingress_nodes_in_flit_valid = io_ingress_0_flit_valid; // @[Nodes.scala 1212:84 NoC.scala 145:78]
  assign router_sink_domain_auto_routers_ingress_nodes_in_flit_bits_head = io_ingress_0_flit_bits_head; // @[Nodes.scala 1212:84 NoC.scala 145:78]
  assign router_sink_domain_auto_routers_ingress_nodes_in_flit_bits_tail = io_ingress_0_flit_bits_tail; // @[Nodes.scala 1212:84 NoC.scala 145:78]
  assign router_sink_domain_auto_routers_ingress_nodes_in_flit_bits_payload = io_ingress_0_flit_bits_payload; // @[Nodes.scala 1212:84 NoC.scala 145:78]
  assign router_sink_domain_auto_routers_ingress_nodes_in_flit_bits_egress_id = io_ingress_0_flit_bits_egress_id; // @[Nodes.scala 1212:84 NoC.scala 145:78]
  assign router_sink_domain_auto_routers_source_nodes_out_1_credit_return =
    router_sink_domain_3_auto_routers_dest_nodes_in_0_credit_return; // @[LazyModule.scala 355:16]
  assign router_sink_domain_auto_routers_source_nodes_out_1_vc_free =
    router_sink_domain_3_auto_routers_dest_nodes_in_0_vc_free; // @[LazyModule.scala 355:16]
  assign router_sink_domain_auto_routers_source_nodes_out_0_credit_return =
    router_sink_domain_1_auto_routers_dest_nodes_in_0_credit_return; // @[LazyModule.scala 355:16]
  assign router_sink_domain_auto_routers_source_nodes_out_0_vc_free =
    router_sink_domain_1_auto_routers_dest_nodes_in_0_vc_free; // @[LazyModule.scala 355:16]
  assign router_sink_domain_auto_clock_in_clock = io_router_clocks_0_clock; // @[Nodes.scala 1212:84 NoC.scala 147:88]
  assign router_sink_domain_auto_clock_in_reset = io_router_clocks_0_reset; // @[Nodes.scala 1212:84 NoC.scala 147:88]
  assign router_sink_domain_1_auto_routers_dest_nodes_in_1_flit_0_valid =
    router_sink_domain_2_auto_routers_source_nodes_out_0_flit_0_valid; // @[LazyModule.scala 353:16]
  assign router_sink_domain_1_auto_routers_dest_nodes_in_1_flit_0_bits_head =
    router_sink_domain_2_auto_routers_source_nodes_out_0_flit_0_bits_head; // @[LazyModule.scala 353:16]
  assign router_sink_domain_1_auto_routers_dest_nodes_in_1_flit_0_bits_tail =
    router_sink_domain_2_auto_routers_source_nodes_out_0_flit_0_bits_tail; // @[LazyModule.scala 353:16]
  assign router_sink_domain_1_auto_routers_dest_nodes_in_1_flit_0_bits_payload =
    router_sink_domain_2_auto_routers_source_nodes_out_0_flit_0_bits_payload; // @[LazyModule.scala 353:16]
  assign router_sink_domain_1_auto_routers_dest_nodes_in_1_flit_0_bits_flow_ingress_node =
    router_sink_domain_2_auto_routers_source_nodes_out_0_flit_0_bits_flow_ingress_node; // @[LazyModule.scala 353:16]
  assign router_sink_domain_1_auto_routers_dest_nodes_in_1_flit_0_bits_flow_egress_node =
    router_sink_domain_2_auto_routers_source_nodes_out_0_flit_0_bits_flow_egress_node; // @[LazyModule.scala 353:16]
  assign router_sink_domain_1_auto_routers_dest_nodes_in_1_flit_0_bits_virt_channel_id =
    router_sink_domain_2_auto_routers_source_nodes_out_0_flit_0_bits_virt_channel_id; // @[LazyModule.scala 353:16]
  assign router_sink_domain_1_auto_routers_dest_nodes_in_0_flit_0_valid =
    router_sink_domain_auto_routers_source_nodes_out_0_flit_0_valid; // @[LazyModule.scala 355:16]
  assign router_sink_domain_1_auto_routers_dest_nodes_in_0_flit_0_bits_head =
    router_sink_domain_auto_routers_source_nodes_out_0_flit_0_bits_head; // @[LazyModule.scala 355:16]
  assign router_sink_domain_1_auto_routers_dest_nodes_in_0_flit_0_bits_tail =
    router_sink_domain_auto_routers_source_nodes_out_0_flit_0_bits_tail; // @[LazyModule.scala 355:16]
  assign router_sink_domain_1_auto_routers_dest_nodes_in_0_flit_0_bits_payload =
    router_sink_domain_auto_routers_source_nodes_out_0_flit_0_bits_payload; // @[LazyModule.scala 355:16]
  assign router_sink_domain_1_auto_routers_dest_nodes_in_0_flit_0_bits_flow_ingress_node =
    router_sink_domain_auto_routers_source_nodes_out_0_flit_0_bits_flow_ingress_node; // @[LazyModule.scala 355:16]
  assign router_sink_domain_1_auto_routers_dest_nodes_in_0_flit_0_bits_flow_egress_node =
    router_sink_domain_auto_routers_source_nodes_out_0_flit_0_bits_flow_egress_node; // @[LazyModule.scala 355:16]
  assign router_sink_domain_1_auto_routers_dest_nodes_in_0_flit_0_bits_virt_channel_id =
    router_sink_domain_auto_routers_source_nodes_out_0_flit_0_bits_virt_channel_id; // @[LazyModule.scala 355:16]
  assign router_sink_domain_1_auto_clock_in_clock = io_router_clocks_1_clock; // @[Nodes.scala 1212:84 NoC.scala 147:88]
  assign router_sink_domain_1_auto_clock_in_reset = io_router_clocks_1_reset; // @[Nodes.scala 1212:84 NoC.scala 147:88]
  assign router_sink_domain_2_auto_routers_ingress_nodes_in_flit_valid = io_ingress_1_flit_valid; // @[Nodes.scala 1212:84 NoC.scala 145:78]
  assign router_sink_domain_2_auto_routers_ingress_nodes_in_flit_bits_head = io_ingress_1_flit_bits_head; // @[Nodes.scala 1212:84 NoC.scala 145:78]
  assign router_sink_domain_2_auto_routers_ingress_nodes_in_flit_bits_tail = io_ingress_1_flit_bits_tail; // @[Nodes.scala 1212:84 NoC.scala 145:78]
  assign router_sink_domain_2_auto_routers_ingress_nodes_in_flit_bits_payload = io_ingress_1_flit_bits_payload; // @[Nodes.scala 1212:84 NoC.scala 145:78]
  assign router_sink_domain_2_auto_routers_ingress_nodes_in_flit_bits_egress_id = io_ingress_1_flit_bits_egress_id; // @[Nodes.scala 1212:84 NoC.scala 145:78]
  assign router_sink_domain_2_auto_routers_source_nodes_out_1_credit_return =
    router_sink_domain_3_auto_routers_dest_nodes_in_1_credit_return; // @[LazyModule.scala 355:16]
  assign router_sink_domain_2_auto_routers_source_nodes_out_1_vc_free =
    router_sink_domain_3_auto_routers_dest_nodes_in_1_vc_free; // @[LazyModule.scala 355:16]
  assign router_sink_domain_2_auto_routers_source_nodes_out_0_credit_return =
    router_sink_domain_1_auto_routers_dest_nodes_in_1_credit_return; // @[LazyModule.scala 353:16]
  assign router_sink_domain_2_auto_routers_source_nodes_out_0_vc_free =
    router_sink_domain_1_auto_routers_dest_nodes_in_1_vc_free; // @[LazyModule.scala 353:16]
  assign router_sink_domain_2_auto_clock_in_clock = io_router_clocks_2_clock; // @[Nodes.scala 1212:84 NoC.scala 147:88]
  assign router_sink_domain_2_auto_clock_in_reset = io_router_clocks_2_reset; // @[Nodes.scala 1212:84 NoC.scala 147:88]
  assign router_sink_domain_3_auto_routers_dest_nodes_in_1_flit_0_valid =
    router_sink_domain_2_auto_routers_source_nodes_out_1_flit_0_valid; // @[LazyModule.scala 355:16]
  assign router_sink_domain_3_auto_routers_dest_nodes_in_1_flit_0_bits_head =
    router_sink_domain_2_auto_routers_source_nodes_out_1_flit_0_bits_head; // @[LazyModule.scala 355:16]
  assign router_sink_domain_3_auto_routers_dest_nodes_in_1_flit_0_bits_tail =
    router_sink_domain_2_auto_routers_source_nodes_out_1_flit_0_bits_tail; // @[LazyModule.scala 355:16]
  assign router_sink_domain_3_auto_routers_dest_nodes_in_1_flit_0_bits_payload =
    router_sink_domain_2_auto_routers_source_nodes_out_1_flit_0_bits_payload; // @[LazyModule.scala 355:16]
  assign router_sink_domain_3_auto_routers_dest_nodes_in_1_flit_0_bits_flow_ingress_node =
    router_sink_domain_2_auto_routers_source_nodes_out_1_flit_0_bits_flow_ingress_node; // @[LazyModule.scala 355:16]
  assign router_sink_domain_3_auto_routers_dest_nodes_in_1_flit_0_bits_flow_egress_node =
    router_sink_domain_2_auto_routers_source_nodes_out_1_flit_0_bits_flow_egress_node; // @[LazyModule.scala 355:16]
  assign router_sink_domain_3_auto_routers_dest_nodes_in_1_flit_0_bits_virt_channel_id =
    router_sink_domain_2_auto_routers_source_nodes_out_1_flit_0_bits_virt_channel_id; // @[LazyModule.scala 355:16]
  assign router_sink_domain_3_auto_routers_dest_nodes_in_0_flit_0_valid =
    router_sink_domain_auto_routers_source_nodes_out_1_flit_0_valid; // @[LazyModule.scala 355:16]
  assign router_sink_domain_3_auto_routers_dest_nodes_in_0_flit_0_bits_head =
    router_sink_domain_auto_routers_source_nodes_out_1_flit_0_bits_head; // @[LazyModule.scala 355:16]
  assign router_sink_domain_3_auto_routers_dest_nodes_in_0_flit_0_bits_tail =
    router_sink_domain_auto_routers_source_nodes_out_1_flit_0_bits_tail; // @[LazyModule.scala 355:16]
  assign router_sink_domain_3_auto_routers_dest_nodes_in_0_flit_0_bits_payload =
    router_sink_domain_auto_routers_source_nodes_out_1_flit_0_bits_payload; // @[LazyModule.scala 355:16]
  assign router_sink_domain_3_auto_routers_dest_nodes_in_0_flit_0_bits_flow_ingress_node =
    router_sink_domain_auto_routers_source_nodes_out_1_flit_0_bits_flow_ingress_node; // @[LazyModule.scala 355:16]
  assign router_sink_domain_3_auto_routers_dest_nodes_in_0_flit_0_bits_flow_egress_node =
    router_sink_domain_auto_routers_source_nodes_out_1_flit_0_bits_flow_egress_node; // @[LazyModule.scala 355:16]
  assign router_sink_domain_3_auto_routers_dest_nodes_in_0_flit_0_bits_virt_channel_id =
    router_sink_domain_auto_routers_source_nodes_out_1_flit_0_bits_virt_channel_id; // @[LazyModule.scala 355:16]
  assign router_sink_domain_3_auto_clock_in_clock = io_router_clocks_3_clock; // @[Nodes.scala 1212:84 NoC.scala 147:88]
  assign router_sink_domain_3_auto_clock_in_reset = io_router_clocks_3_reset; // @[Nodes.scala 1212:84 NoC.scala 147:88]
  always @(posedge clock) begin
    if (reset) begin // @[NoC.scala 160:37]
      debug_va_stall_ctr <= 64'h0; // @[NoC.scala 160:37]
    end else begin
      debug_va_stall_ctr <= _debug_va_stall_ctr_T_11; // @[NoC.scala 163:24]
    end
    if (reset) begin // @[NoC.scala 161:37]
      debug_sa_stall_ctr <= 64'h0; // @[NoC.scala 161:37]
    end else begin
      debug_sa_stall_ctr <= _debug_sa_stall_ctr_T_11; // @[NoC.scala 164:24]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  debug_va_stall_ctr = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  debug_sa_stall_ctr = _RAND_1[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MaxPeriodFibonacciLFSR(
  input   clock,
  input   reset,
  output  io_out_0,
  output  io_out_1,
  output  io_out_2,
  output  io_out_3,
  output  io_out_4,
  output  io_out_5,
  output  io_out_6,
  output  io_out_7,
  output  io_out_8,
  output  io_out_9,
  output  io_out_10,
  output  io_out_11,
  output  io_out_12,
  output  io_out_13,
  output  io_out_14,
  output  io_out_15,
  output  io_out_16,
  output  io_out_17,
  output  io_out_18,
  output  io_out_19
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
`endif // RANDOMIZE_REG_INIT
  reg  state_0; // @[PRNG.scala 55:49]
  reg  state_1; // @[PRNG.scala 55:49]
  reg  state_2; // @[PRNG.scala 55:49]
  reg  state_3; // @[PRNG.scala 55:49]
  reg  state_4; // @[PRNG.scala 55:49]
  reg  state_5; // @[PRNG.scala 55:49]
  reg  state_6; // @[PRNG.scala 55:49]
  reg  state_7; // @[PRNG.scala 55:49]
  reg  state_8; // @[PRNG.scala 55:49]
  reg  state_9; // @[PRNG.scala 55:49]
  reg  state_10; // @[PRNG.scala 55:49]
  reg  state_11; // @[PRNG.scala 55:49]
  reg  state_12; // @[PRNG.scala 55:49]
  reg  state_13; // @[PRNG.scala 55:49]
  reg  state_14; // @[PRNG.scala 55:49]
  reg  state_15; // @[PRNG.scala 55:49]
  reg  state_16; // @[PRNG.scala 55:49]
  reg  state_17; // @[PRNG.scala 55:49]
  reg  state_18; // @[PRNG.scala 55:49]
  reg  state_19; // @[PRNG.scala 55:49]
  wire  _T = state_19 ^ state_16; // @[LFSR.scala 15:41]
  assign io_out_0 = state_0; // @[PRNG.scala 78:10]
  assign io_out_1 = state_1; // @[PRNG.scala 78:10]
  assign io_out_2 = state_2; // @[PRNG.scala 78:10]
  assign io_out_3 = state_3; // @[PRNG.scala 78:10]
  assign io_out_4 = state_4; // @[PRNG.scala 78:10]
  assign io_out_5 = state_5; // @[PRNG.scala 78:10]
  assign io_out_6 = state_6; // @[PRNG.scala 78:10]
  assign io_out_7 = state_7; // @[PRNG.scala 78:10]
  assign io_out_8 = state_8; // @[PRNG.scala 78:10]
  assign io_out_9 = state_9; // @[PRNG.scala 78:10]
  assign io_out_10 = state_10; // @[PRNG.scala 78:10]
  assign io_out_11 = state_11; // @[PRNG.scala 78:10]
  assign io_out_12 = state_12; // @[PRNG.scala 78:10]
  assign io_out_13 = state_13; // @[PRNG.scala 78:10]
  assign io_out_14 = state_14; // @[PRNG.scala 78:10]
  assign io_out_15 = state_15; // @[PRNG.scala 78:10]
  assign io_out_16 = state_16; // @[PRNG.scala 78:10]
  assign io_out_17 = state_17; // @[PRNG.scala 78:10]
  assign io_out_18 = state_18; // @[PRNG.scala 78:10]
  assign io_out_19 = state_19; // @[PRNG.scala 78:10]
  always @(posedge clock) begin
    state_0 <= reset | _T; // @[PRNG.scala 55:{49,49}]
    if (reset) begin // @[PRNG.scala 55:49]
      state_1 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_1 <= state_0;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_2 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_2 <= state_1;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_3 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_3 <= state_2;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_4 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_4 <= state_3;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_5 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_5 <= state_4;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_6 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_6 <= state_5;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_7 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_7 <= state_6;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_8 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_8 <= state_7;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_9 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_9 <= state_8;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_10 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_10 <= state_9;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_11 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_11 <= state_10;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_12 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_12 <= state_11;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_13 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_13 <= state_12;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_14 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_14 <= state_13;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_15 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_15 <= state_14;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_16 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_16 <= state_15;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_17 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_17 <= state_16;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_18 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_18 <= state_17;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_19 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_19 <= state_18;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  state_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  state_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  state_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  state_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  state_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  state_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  state_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  state_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  state_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  state_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  state_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  state_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  state_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  state_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  state_15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  state_16 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  state_17 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  state_18 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  state_19 = _RAND_19[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module InputGen(
  input         clock,
  input         reset,
  input         io_out_ready,
  output        io_out_valid,
  output        io_out_bits_head,
  output        io_out_bits_tail,
  output [63:0] io_out_bits_payload,
  output        io_out_bits_egress_id,
  input         io_rob_ready,
  input  [6:0]  io_rob_idx,
  input  [31:0] io_tsc,
  output        io_fire,
  output [3:0]  io_n_flits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  packet_remaining_prng_clock; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_reset; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_0; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_1; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_2; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_3; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_4; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_5; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_6; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_7; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_8; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_9; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_10; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_11; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_12; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_13; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_14; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_15; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_16; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_17; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_18; // @[PRNG.scala 91:22]
  wire  packet_remaining_prng_io_out_19; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_clock; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_reset; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_0; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_1; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_2; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_3; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_4; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_5; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_6; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_7; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_8; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_9; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_10; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_11; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_12; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_13; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_14; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_15; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_16; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_17; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_18; // @[PRNG.scala 91:22]
  wire  random_flit_delay_prng_io_out_19; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_clock; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_reset; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_0; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_1; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_2; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_3; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_4; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_5; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_6; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_7; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_8; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_9; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_10; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_11; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_12; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_13; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_14; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_15; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_16; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_17; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_18; // @[PRNG.scala 91:22]
  wire  random_packet_delay_prng_io_out_19; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_clock; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_reset; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_0; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_1; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_2; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_3; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_4; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_5; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_6; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_7; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_8; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_9; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_10; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_11; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_12; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_13; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_14; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_15; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_16; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_17; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_18; // @[PRNG.scala 91:22]
  wire  io_out_bits_egress_id_prng_io_out_19; // @[PRNG.scala 91:22]
  reg [3:0] flits_left; // @[TestHarness.scala 71:27]
  reg [3:0] flits_fired; // @[TestHarness.scala 72:28]
  reg  egress; // @[TestHarness.scala 73:19]
  reg [31:0] payload_tsc; // @[TestHarness.scala 74:20]
  reg [15:0] payload_rob_idx; // @[TestHarness.scala 74:20]
  wire  can_fire = flits_left == 4'h0 & io_rob_ready; // @[TestHarness.scala 76:39]
  wire [9:0] packet_remaining_lo = {packet_remaining_prng_io_out_9,packet_remaining_prng_io_out_8,
    packet_remaining_prng_io_out_7,packet_remaining_prng_io_out_6,packet_remaining_prng_io_out_5,
    packet_remaining_prng_io_out_4,packet_remaining_prng_io_out_3,packet_remaining_prng_io_out_2,
    packet_remaining_prng_io_out_1,packet_remaining_prng_io_out_0}; // @[PRNG.scala 95:17]
  wire [9:0] packet_remaining_hi = {packet_remaining_prng_io_out_19,packet_remaining_prng_io_out_18,
    packet_remaining_prng_io_out_17,packet_remaining_prng_io_out_16,packet_remaining_prng_io_out_15,
    packet_remaining_prng_io_out_14,packet_remaining_prng_io_out_13,packet_remaining_prng_io_out_12,
    packet_remaining_prng_io_out_11,packet_remaining_prng_io_out_10}; // @[PRNG.scala 95:17]
  wire [19:0] _packet_remaining_T = {packet_remaining_hi,packet_remaining_lo}; // @[PRNG.scala 95:17]
  wire [19:0] _GEN_0 = _packet_remaining_T % 20'h8; // @[TestHarness.scala 78:89]
  wire [3:0] packet_remaining = _GEN_0[3:0]; // @[TestHarness.scala 78:89]
  wire [9:0] io_out_bits_egress_id_lo = {io_out_bits_egress_id_prng_io_out_9,io_out_bits_egress_id_prng_io_out_8,
    io_out_bits_egress_id_prng_io_out_7,io_out_bits_egress_id_prng_io_out_6,io_out_bits_egress_id_prng_io_out_5,
    io_out_bits_egress_id_prng_io_out_4,io_out_bits_egress_id_prng_io_out_3,io_out_bits_egress_id_prng_io_out_2,
    io_out_bits_egress_id_prng_io_out_1,io_out_bits_egress_id_prng_io_out_0}; // @[PRNG.scala 95:17]
  wire [9:0] io_out_bits_egress_id_hi = {io_out_bits_egress_id_prng_io_out_19,io_out_bits_egress_id_prng_io_out_18,
    io_out_bits_egress_id_prng_io_out_17,io_out_bits_egress_id_prng_io_out_16,io_out_bits_egress_id_prng_io_out_15,
    io_out_bits_egress_id_prng_io_out_14,io_out_bits_egress_id_prng_io_out_13,io_out_bits_egress_id_prng_io_out_12,
    io_out_bits_egress_id_prng_io_out_11,io_out_bits_egress_id_prng_io_out_10}; // @[PRNG.scala 95:17]
  wire [19:0] _io_out_bits_egress_id_T = {io_out_bits_egress_id_hi,io_out_bits_egress_id_lo}; // @[PRNG.scala 95:17]
  wire [19:0] _GEN_1 = _io_out_bits_egress_id_T % 20'h2; // @[TestHarness.scala 84:92]
  wire [31:0] out_payload_tsc = flits_left != 4'h0 ? payload_tsc : io_tsc; // @[TestHarness.scala 100:29 105:17 87:19]
  wire [15:0] out_payload_rob_idx = flits_left != 4'h0 ? payload_rob_idx : {{9'd0}, io_rob_idx}; // @[TestHarness.scala 100:29 105:17 88:23]
  wire [47:0] io_out_bits_payload_hi = {out_payload_tsc,out_payload_rob_idx}; // @[TestHarness.scala 86:38]
  wire [3:0] _GEN_16 = flits_left != 4'h0 ? flits_fired : 4'h0; // @[TestHarness.scala 100:29 106:29 89:27]
  wire [15:0] out_payload_flits_fired = {{12'd0}, _GEN_16}; // @[TestHarness.scala 85:25]
  wire  _io_fire_T = io_out_ready & io_out_valid; // @[Decoupled.scala 51:35]
  wire [3:0] _GEN_2 = io_fire & ~io_out_bits_tail ? packet_remaining : flits_left; // @[TestHarness.scala 94:39 95:16 71:27]
  wire [3:0] _GEN_7 = io_fire & ~io_out_bits_tail ? 4'h1 : flits_fired; // @[TestHarness.scala 94:39 98:17 72:28]
  wire [3:0] _flits_fired_T_1 = flits_fired + 4'h1; // @[TestHarness.scala 109:34]
  wire [3:0] _flits_left_T_1 = flits_left - 4'h1; // @[TestHarness.scala 110:32]
  MaxPeriodFibonacciLFSR packet_remaining_prng ( // @[PRNG.scala 91:22]
    .clock(packet_remaining_prng_clock),
    .reset(packet_remaining_prng_reset),
    .io_out_0(packet_remaining_prng_io_out_0),
    .io_out_1(packet_remaining_prng_io_out_1),
    .io_out_2(packet_remaining_prng_io_out_2),
    .io_out_3(packet_remaining_prng_io_out_3),
    .io_out_4(packet_remaining_prng_io_out_4),
    .io_out_5(packet_remaining_prng_io_out_5),
    .io_out_6(packet_remaining_prng_io_out_6),
    .io_out_7(packet_remaining_prng_io_out_7),
    .io_out_8(packet_remaining_prng_io_out_8),
    .io_out_9(packet_remaining_prng_io_out_9),
    .io_out_10(packet_remaining_prng_io_out_10),
    .io_out_11(packet_remaining_prng_io_out_11),
    .io_out_12(packet_remaining_prng_io_out_12),
    .io_out_13(packet_remaining_prng_io_out_13),
    .io_out_14(packet_remaining_prng_io_out_14),
    .io_out_15(packet_remaining_prng_io_out_15),
    .io_out_16(packet_remaining_prng_io_out_16),
    .io_out_17(packet_remaining_prng_io_out_17),
    .io_out_18(packet_remaining_prng_io_out_18),
    .io_out_19(packet_remaining_prng_io_out_19)
  );
  MaxPeriodFibonacciLFSR random_flit_delay_prng ( // @[PRNG.scala 91:22]
    .clock(random_flit_delay_prng_clock),
    .reset(random_flit_delay_prng_reset),
    .io_out_0(random_flit_delay_prng_io_out_0),
    .io_out_1(random_flit_delay_prng_io_out_1),
    .io_out_2(random_flit_delay_prng_io_out_2),
    .io_out_3(random_flit_delay_prng_io_out_3),
    .io_out_4(random_flit_delay_prng_io_out_4),
    .io_out_5(random_flit_delay_prng_io_out_5),
    .io_out_6(random_flit_delay_prng_io_out_6),
    .io_out_7(random_flit_delay_prng_io_out_7),
    .io_out_8(random_flit_delay_prng_io_out_8),
    .io_out_9(random_flit_delay_prng_io_out_9),
    .io_out_10(random_flit_delay_prng_io_out_10),
    .io_out_11(random_flit_delay_prng_io_out_11),
    .io_out_12(random_flit_delay_prng_io_out_12),
    .io_out_13(random_flit_delay_prng_io_out_13),
    .io_out_14(random_flit_delay_prng_io_out_14),
    .io_out_15(random_flit_delay_prng_io_out_15),
    .io_out_16(random_flit_delay_prng_io_out_16),
    .io_out_17(random_flit_delay_prng_io_out_17),
    .io_out_18(random_flit_delay_prng_io_out_18),
    .io_out_19(random_flit_delay_prng_io_out_19)
  );
  MaxPeriodFibonacciLFSR random_packet_delay_prng ( // @[PRNG.scala 91:22]
    .clock(random_packet_delay_prng_clock),
    .reset(random_packet_delay_prng_reset),
    .io_out_0(random_packet_delay_prng_io_out_0),
    .io_out_1(random_packet_delay_prng_io_out_1),
    .io_out_2(random_packet_delay_prng_io_out_2),
    .io_out_3(random_packet_delay_prng_io_out_3),
    .io_out_4(random_packet_delay_prng_io_out_4),
    .io_out_5(random_packet_delay_prng_io_out_5),
    .io_out_6(random_packet_delay_prng_io_out_6),
    .io_out_7(random_packet_delay_prng_io_out_7),
    .io_out_8(random_packet_delay_prng_io_out_8),
    .io_out_9(random_packet_delay_prng_io_out_9),
    .io_out_10(random_packet_delay_prng_io_out_10),
    .io_out_11(random_packet_delay_prng_io_out_11),
    .io_out_12(random_packet_delay_prng_io_out_12),
    .io_out_13(random_packet_delay_prng_io_out_13),
    .io_out_14(random_packet_delay_prng_io_out_14),
    .io_out_15(random_packet_delay_prng_io_out_15),
    .io_out_16(random_packet_delay_prng_io_out_16),
    .io_out_17(random_packet_delay_prng_io_out_17),
    .io_out_18(random_packet_delay_prng_io_out_18),
    .io_out_19(random_packet_delay_prng_io_out_19)
  );
  MaxPeriodFibonacciLFSR io_out_bits_egress_id_prng ( // @[PRNG.scala 91:22]
    .clock(io_out_bits_egress_id_prng_clock),
    .reset(io_out_bits_egress_id_prng_reset),
    .io_out_0(io_out_bits_egress_id_prng_io_out_0),
    .io_out_1(io_out_bits_egress_id_prng_io_out_1),
    .io_out_2(io_out_bits_egress_id_prng_io_out_2),
    .io_out_3(io_out_bits_egress_id_prng_io_out_3),
    .io_out_4(io_out_bits_egress_id_prng_io_out_4),
    .io_out_5(io_out_bits_egress_id_prng_io_out_5),
    .io_out_6(io_out_bits_egress_id_prng_io_out_6),
    .io_out_7(io_out_bits_egress_id_prng_io_out_7),
    .io_out_8(io_out_bits_egress_id_prng_io_out_8),
    .io_out_9(io_out_bits_egress_id_prng_io_out_9),
    .io_out_10(io_out_bits_egress_id_prng_io_out_10),
    .io_out_11(io_out_bits_egress_id_prng_io_out_11),
    .io_out_12(io_out_bits_egress_id_prng_io_out_12),
    .io_out_13(io_out_bits_egress_id_prng_io_out_13),
    .io_out_14(io_out_bits_egress_id_prng_io_out_14),
    .io_out_15(io_out_bits_egress_id_prng_io_out_15),
    .io_out_16(io_out_bits_egress_id_prng_io_out_16),
    .io_out_17(io_out_bits_egress_id_prng_io_out_17),
    .io_out_18(io_out_bits_egress_id_prng_io_out_18),
    .io_out_19(io_out_bits_egress_id_prng_io_out_19)
  );
  assign io_out_valid = flits_left != 4'h0 | can_fire; // @[TestHarness.scala 100:29 101:18 81:16]
  assign io_out_bits_head = flits_left != 4'h0 ? 1'h0 : 1'h1; // @[TestHarness.scala 100:29 102:22 82:20]
  assign io_out_bits_tail = flits_left != 4'h0 ? flits_left == 4'h1 : packet_remaining == 4'h0; // @[TestHarness.scala 100:29 103:22 83:20]
  assign io_out_bits_payload = {io_out_bits_payload_hi,out_payload_flits_fired}; // @[TestHarness.scala 86:38]
  assign io_out_bits_egress_id = flits_left != 4'h0 ? egress : _GEN_1[0]; // @[TestHarness.scala 100:29 104:27 84:25]
  assign io_fire = can_fire & _io_fire_T; // @[TestHarness.scala 92:23]
  assign io_n_flits = packet_remaining + 4'h1; // @[TestHarness.scala 91:34]
  assign packet_remaining_prng_clock = clock;
  assign packet_remaining_prng_reset = reset;
  assign random_flit_delay_prng_clock = clock;
  assign random_flit_delay_prng_reset = reset;
  assign random_packet_delay_prng_clock = clock;
  assign random_packet_delay_prng_reset = reset;
  assign io_out_bits_egress_id_prng_clock = clock;
  assign io_out_bits_egress_id_prng_reset = reset;
  always @(posedge clock) begin
    if (reset) begin // @[TestHarness.scala 71:27]
      flits_left <= 4'h0; // @[TestHarness.scala 71:27]
    end else if (flits_left != 4'h0) begin // @[TestHarness.scala 100:29]
      if (_io_fire_T) begin // @[TestHarness.scala 108:26]
        flits_left <= _flits_left_T_1; // @[TestHarness.scala 110:18]
      end else begin
        flits_left <= _GEN_2;
      end
    end else begin
      flits_left <= _GEN_2;
    end
    if (reset) begin // @[TestHarness.scala 72:28]
      flits_fired <= 4'h0; // @[TestHarness.scala 72:28]
    end else if (flits_left != 4'h0) begin // @[TestHarness.scala 100:29]
      if (_io_fire_T) begin // @[TestHarness.scala 108:26]
        flits_fired <= _flits_fired_T_1; // @[TestHarness.scala 109:19]
      end else begin
        flits_fired <= _GEN_7;
      end
    end else begin
      flits_fired <= _GEN_7;
    end
    if (io_fire & ~io_out_bits_tail) begin // @[TestHarness.scala 94:39]
      egress <= io_out_bits_egress_id; // @[TestHarness.scala 97:12]
    end
    if (io_fire & ~io_out_bits_tail) begin // @[TestHarness.scala 94:39]
      if (!(flits_left != 4'h0)) begin // @[TestHarness.scala 100:29]
        payload_tsc <= io_tsc; // @[TestHarness.scala 87:19]
      end
    end
    if (io_fire & ~io_out_bits_tail) begin // @[TestHarness.scala 94:39]
      if (!(flits_left != 4'h0)) begin // @[TestHarness.scala 100:29]
        payload_rob_idx <= {{9'd0}, io_rob_idx}; // @[TestHarness.scala 88:23]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  flits_left = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  flits_fired = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  egress = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  payload_tsc = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  payload_rob_idx = _RAND_4[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_26(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_head,
  input         io_enq_bits_tail,
  input  [63:0] io_enq_bits_payload,
  input         io_enq_bits_egress_id,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_head,
  output        io_deq_bits_tail,
  output [63:0] io_deq_bits_payload,
  output        io_deq_bits_egress_id
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg  ram_head [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_head_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_head_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_head_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_head_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_tail [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_tail_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_tail_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_tail_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_tail_MPORT_en; // @[Decoupled.scala 273:95]
  reg [63:0] ram_payload [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_payload_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_payload_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [63:0] ram_payload_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [63:0] ram_payload_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_payload_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_payload_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_payload_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_egress_id [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_egress_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_egress_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_egress_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_egress_id_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_egress_id_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_egress_id_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_egress_id_MPORT_en; // @[Decoupled.scala 273:95]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 278:28]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  wire  _GEN_12 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 318:26 280:27 318:35]
  wire  do_enq = empty ? _GEN_12 : _do_enq_T; // @[Decoupled.scala 315:17 280:27]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 315:17 317:14 281:27]
  assign ram_head_io_deq_bits_MPORT_en = 1'h1;
  assign ram_head_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_head_io_deq_bits_MPORT_data = ram_head[ram_head_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_head_MPORT_data = io_enq_bits_head;
  assign ram_head_MPORT_addr = 1'h0;
  assign ram_head_MPORT_mask = 1'h1;
  assign ram_head_MPORT_en = empty ? _GEN_12 : _do_enq_T;
  assign ram_tail_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tail_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tail_io_deq_bits_MPORT_data = ram_tail[ram_tail_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_tail_MPORT_data = io_enq_bits_tail;
  assign ram_tail_MPORT_addr = 1'h0;
  assign ram_tail_MPORT_mask = 1'h1;
  assign ram_tail_MPORT_en = empty ? _GEN_12 : _do_enq_T;
  assign ram_payload_io_deq_bits_MPORT_en = 1'h1;
  assign ram_payload_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_payload_io_deq_bits_MPORT_data = ram_payload[ram_payload_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_payload_MPORT_data = io_enq_bits_payload;
  assign ram_payload_MPORT_addr = 1'h0;
  assign ram_payload_MPORT_mask = 1'h1;
  assign ram_payload_MPORT_en = empty ? _GEN_12 : _do_enq_T;
  assign ram_egress_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_egress_id_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_egress_id_io_deq_bits_MPORT_data = ram_egress_id[ram_egress_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_egress_id_MPORT_data = io_enq_bits_egress_id;
  assign ram_egress_id_MPORT_addr = 1'h0;
  assign ram_egress_id_MPORT_mask = 1'h1;
  assign ram_egress_id_MPORT_en = empty ? _GEN_12 : _do_enq_T;
  assign io_enq_ready = io_deq_ready | empty; // @[Decoupled.scala 303:16 323:{24,39}]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 302:16 314:{24,39}]
  assign io_deq_bits_head = empty ? io_enq_bits_head : ram_head_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_tail = empty ? io_enq_bits_tail : ram_tail_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_payload = empty ? io_enq_bits_payload : ram_payload_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  assign io_deq_bits_egress_id = empty ? io_enq_bits_egress_id : ram_egress_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17 315:17 316:19]
  always @(posedge clock) begin
    if (ram_head_MPORT_en & ram_head_MPORT_mask) begin
      ram_head[ram_head_MPORT_addr] <= ram_head_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_tail_MPORT_en & ram_tail_MPORT_mask) begin
      ram_tail[ram_tail_MPORT_addr] <= ram_tail_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_payload_MPORT_en & ram_payload_MPORT_mask) begin
      ram_payload[ram_payload_MPORT_addr] <= ram_payload_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_egress_id_MPORT_en & ram_egress_id_MPORT_mask) begin
      ram_egress_id[ram_egress_id_MPORT_addr] <= ram_egress_id_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      if (empty) begin // @[Decoupled.scala 315:17]
        if (io_deq_ready) begin // @[Decoupled.scala 318:26]
          maybe_full <= 1'h0; // @[Decoupled.scala 318:35]
        end else begin
          maybe_full <= _do_enq_T; // @[Decoupled.scala 280:27]
        end
      end else begin
        maybe_full <= _do_enq_T; // @[Decoupled.scala 280:27]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_head[initvar] = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tail[initvar] = _RAND_1[0:0];
  _RAND_2 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload[initvar] = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_egress_id[initvar] = _RAND_3[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  maybe_full = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module NoCTester(
  input         clock,
  input         reset,
  input         io_to_noc_1_flit_ready,
  output        io_to_noc_1_flit_valid,
  output        io_to_noc_1_flit_bits_head,
  output        io_to_noc_1_flit_bits_tail,
  output [63:0] io_to_noc_1_flit_bits_payload,
  output        io_to_noc_1_flit_bits_egress_id,
  input         io_to_noc_0_flit_ready,
  output        io_to_noc_0_flit_valid,
  output        io_to_noc_0_flit_bits_head,
  output        io_to_noc_0_flit_bits_tail,
  output [63:0] io_to_noc_0_flit_bits_payload,
  output        io_to_noc_0_flit_bits_egress_id,
  output        io_from_noc_1_flit_ready,
  input         io_from_noc_1_flit_valid,
  input         io_from_noc_1_flit_bits_head,
  input         io_from_noc_1_flit_bits_tail,
  input  [63:0] io_from_noc_1_flit_bits_payload,
  input         io_from_noc_1_flit_bits_ingress_id,
  output        io_from_noc_0_flit_ready,
  input         io_from_noc_0_flit_valid,
  input         io_from_noc_0_flit_bits_head,
  input         io_from_noc_0_flit_bits_tail,
  input  [63:0] io_from_noc_0_flit_bits_payload,
  input         io_from_noc_0_flit_bits_ingress_id,
  output        io_success
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [127:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [63:0] _RAND_901;
  reg [63:0] _RAND_902;
  reg [63:0] _RAND_903;
  reg [63:0] _RAND_904;
  reg [63:0] _RAND_905;
  reg [63:0] _RAND_906;
  reg [63:0] _RAND_907;
  reg [63:0] _RAND_908;
  reg [63:0] _RAND_909;
  reg [63:0] _RAND_910;
  reg [63:0] _RAND_911;
  reg [63:0] _RAND_912;
  reg [63:0] _RAND_913;
  reg [63:0] _RAND_914;
  reg [63:0] _RAND_915;
  reg [63:0] _RAND_916;
  reg [63:0] _RAND_917;
  reg [63:0] _RAND_918;
  reg [63:0] _RAND_919;
  reg [63:0] _RAND_920;
  reg [63:0] _RAND_921;
  reg [63:0] _RAND_922;
  reg [63:0] _RAND_923;
  reg [63:0] _RAND_924;
  reg [63:0] _RAND_925;
  reg [63:0] _RAND_926;
  reg [63:0] _RAND_927;
  reg [63:0] _RAND_928;
  reg [63:0] _RAND_929;
  reg [63:0] _RAND_930;
  reg [63:0] _RAND_931;
  reg [63:0] _RAND_932;
  reg [63:0] _RAND_933;
  reg [63:0] _RAND_934;
  reg [63:0] _RAND_935;
  reg [63:0] _RAND_936;
  reg [63:0] _RAND_937;
  reg [63:0] _RAND_938;
  reg [63:0] _RAND_939;
  reg [63:0] _RAND_940;
  reg [63:0] _RAND_941;
  reg [63:0] _RAND_942;
  reg [63:0] _RAND_943;
  reg [63:0] _RAND_944;
  reg [63:0] _RAND_945;
  reg [63:0] _RAND_946;
  reg [63:0] _RAND_947;
  reg [63:0] _RAND_948;
  reg [63:0] _RAND_949;
  reg [63:0] _RAND_950;
  reg [63:0] _RAND_951;
  reg [63:0] _RAND_952;
  reg [63:0] _RAND_953;
  reg [63:0] _RAND_954;
  reg [63:0] _RAND_955;
  reg [63:0] _RAND_956;
  reg [63:0] _RAND_957;
  reg [63:0] _RAND_958;
  reg [63:0] _RAND_959;
  reg [63:0] _RAND_960;
  reg [63:0] _RAND_961;
  reg [63:0] _RAND_962;
  reg [63:0] _RAND_963;
  reg [63:0] _RAND_964;
  reg [63:0] _RAND_965;
  reg [63:0] _RAND_966;
  reg [63:0] _RAND_967;
  reg [63:0] _RAND_968;
  reg [63:0] _RAND_969;
  reg [63:0] _RAND_970;
  reg [63:0] _RAND_971;
  reg [63:0] _RAND_972;
  reg [63:0] _RAND_973;
  reg [63:0] _RAND_974;
  reg [63:0] _RAND_975;
  reg [63:0] _RAND_976;
  reg [63:0] _RAND_977;
  reg [63:0] _RAND_978;
  reg [63:0] _RAND_979;
  reg [63:0] _RAND_980;
  reg [63:0] _RAND_981;
  reg [63:0] _RAND_982;
  reg [63:0] _RAND_983;
  reg [63:0] _RAND_984;
  reg [63:0] _RAND_985;
  reg [63:0] _RAND_986;
  reg [63:0] _RAND_987;
  reg [63:0] _RAND_988;
  reg [63:0] _RAND_989;
  reg [63:0] _RAND_990;
  reg [63:0] _RAND_991;
  reg [63:0] _RAND_992;
  reg [63:0] _RAND_993;
  reg [63:0] _RAND_994;
  reg [63:0] _RAND_995;
  reg [63:0] _RAND_996;
  reg [63:0] _RAND_997;
  reg [63:0] _RAND_998;
  reg [63:0] _RAND_999;
  reg [63:0] _RAND_1000;
  reg [63:0] _RAND_1001;
  reg [63:0] _RAND_1002;
  reg [63:0] _RAND_1003;
  reg [63:0] _RAND_1004;
  reg [63:0] _RAND_1005;
  reg [63:0] _RAND_1006;
  reg [63:0] _RAND_1007;
  reg [63:0] _RAND_1008;
  reg [63:0] _RAND_1009;
  reg [63:0] _RAND_1010;
  reg [63:0] _RAND_1011;
  reg [63:0] _RAND_1012;
  reg [63:0] _RAND_1013;
  reg [63:0] _RAND_1014;
  reg [63:0] _RAND_1015;
  reg [63:0] _RAND_1016;
  reg [63:0] _RAND_1017;
  reg [63:0] _RAND_1018;
  reg [63:0] _RAND_1019;
  reg [63:0] _RAND_1020;
  reg [63:0] _RAND_1021;
  reg [63:0] _RAND_1022;
  reg [63:0] _RAND_1023;
  reg [63:0] _RAND_1024;
  reg [63:0] _RAND_1025;
  reg [63:0] _RAND_1026;
  reg [63:0] _RAND_1027;
  reg [63:0] _RAND_1028;
  reg [31:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
`endif // RANDOMIZE_REG_INIT
  wire  igen_clock; // @[TestHarness.scala 171:22]
  wire  igen_reset; // @[TestHarness.scala 171:22]
  wire  igen_io_out_ready; // @[TestHarness.scala 171:22]
  wire  igen_io_out_valid; // @[TestHarness.scala 171:22]
  wire  igen_io_out_bits_head; // @[TestHarness.scala 171:22]
  wire  igen_io_out_bits_tail; // @[TestHarness.scala 171:22]
  wire [63:0] igen_io_out_bits_payload; // @[TestHarness.scala 171:22]
  wire  igen_io_out_bits_egress_id; // @[TestHarness.scala 171:22]
  wire  igen_io_rob_ready; // @[TestHarness.scala 171:22]
  wire [6:0] igen_io_rob_idx; // @[TestHarness.scala 171:22]
  wire [31:0] igen_io_tsc; // @[TestHarness.scala 171:22]
  wire  igen_io_fire; // @[TestHarness.scala 171:22]
  wire [3:0] igen_io_n_flits; // @[TestHarness.scala 171:22]
  wire  io_to_noc_0_flit_q_clock; // @[Decoupled.scala 375:21]
  wire  io_to_noc_0_flit_q_reset; // @[Decoupled.scala 375:21]
  wire  io_to_noc_0_flit_q_io_enq_ready; // @[Decoupled.scala 375:21]
  wire  io_to_noc_0_flit_q_io_enq_valid; // @[Decoupled.scala 375:21]
  wire  io_to_noc_0_flit_q_io_enq_bits_head; // @[Decoupled.scala 375:21]
  wire  io_to_noc_0_flit_q_io_enq_bits_tail; // @[Decoupled.scala 375:21]
  wire [63:0] io_to_noc_0_flit_q_io_enq_bits_payload; // @[Decoupled.scala 375:21]
  wire  io_to_noc_0_flit_q_io_enq_bits_egress_id; // @[Decoupled.scala 375:21]
  wire  io_to_noc_0_flit_q_io_deq_ready; // @[Decoupled.scala 375:21]
  wire  io_to_noc_0_flit_q_io_deq_valid; // @[Decoupled.scala 375:21]
  wire  io_to_noc_0_flit_q_io_deq_bits_head; // @[Decoupled.scala 375:21]
  wire  io_to_noc_0_flit_q_io_deq_bits_tail; // @[Decoupled.scala 375:21]
  wire [63:0] io_to_noc_0_flit_q_io_deq_bits_payload; // @[Decoupled.scala 375:21]
  wire  io_to_noc_0_flit_q_io_deq_bits_egress_id; // @[Decoupled.scala 375:21]
  wire  igen_1_clock; // @[TestHarness.scala 171:22]
  wire  igen_1_reset; // @[TestHarness.scala 171:22]
  wire  igen_1_io_out_ready; // @[TestHarness.scala 171:22]
  wire  igen_1_io_out_valid; // @[TestHarness.scala 171:22]
  wire  igen_1_io_out_bits_head; // @[TestHarness.scala 171:22]
  wire  igen_1_io_out_bits_tail; // @[TestHarness.scala 171:22]
  wire [63:0] igen_1_io_out_bits_payload; // @[TestHarness.scala 171:22]
  wire  igen_1_io_out_bits_egress_id; // @[TestHarness.scala 171:22]
  wire  igen_1_io_rob_ready; // @[TestHarness.scala 171:22]
  wire [6:0] igen_1_io_rob_idx; // @[TestHarness.scala 171:22]
  wire [31:0] igen_1_io_tsc; // @[TestHarness.scala 171:22]
  wire  igen_1_io_fire; // @[TestHarness.scala 171:22]
  wire [3:0] igen_1_io_n_flits; // @[TestHarness.scala 171:22]
  wire  io_to_noc_1_flit_q_clock; // @[Decoupled.scala 375:21]
  wire  io_to_noc_1_flit_q_reset; // @[Decoupled.scala 375:21]
  wire  io_to_noc_1_flit_q_io_enq_ready; // @[Decoupled.scala 375:21]
  wire  io_to_noc_1_flit_q_io_enq_valid; // @[Decoupled.scala 375:21]
  wire  io_to_noc_1_flit_q_io_enq_bits_head; // @[Decoupled.scala 375:21]
  wire  io_to_noc_1_flit_q_io_enq_bits_tail; // @[Decoupled.scala 375:21]
  wire [63:0] io_to_noc_1_flit_q_io_enq_bits_payload; // @[Decoupled.scala 375:21]
  wire  io_to_noc_1_flit_q_io_enq_bits_egress_id; // @[Decoupled.scala 375:21]
  wire  io_to_noc_1_flit_q_io_deq_ready; // @[Decoupled.scala 375:21]
  wire  io_to_noc_1_flit_q_io_deq_valid; // @[Decoupled.scala 375:21]
  wire  io_to_noc_1_flit_q_io_deq_bits_head; // @[Decoupled.scala 375:21]
  wire  io_to_noc_1_flit_q_io_deq_bits_tail; // @[Decoupled.scala 375:21]
  wire [63:0] io_to_noc_1_flit_q_io_deq_bits_payload; // @[Decoupled.scala 375:21]
  wire  io_to_noc_1_flit_q_io_deq_bits_egress_id; // @[Decoupled.scala 375:21]
  wire  plusarg_reader_out; // @[PlusArg.scala 80:11]
  wire  io_from_noc_0_flit_ready_prng_clock; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_reset; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_0; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_1; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_2; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_3; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_4; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_5; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_6; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_7; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_8; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_9; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_10; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_11; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_12; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_13; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_14; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_15; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_16; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_17; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_18; // @[PRNG.scala 91:22]
  wire  io_from_noc_0_flit_ready_prng_io_out_19; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_clock; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_reset; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_io_out_0; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_io_out_1; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_io_out_2; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_io_out_3; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_io_out_4; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_io_out_5; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_io_out_6; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_io_out_7; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_io_out_8; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_io_out_9; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_io_out_10; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_io_out_11; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_io_out_12; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_io_out_13; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_io_out_14; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_io_out_15; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_io_out_16; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_io_out_17; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_io_out_18; // @[PRNG.scala 91:22]
  wire  io_from_noc_1_flit_ready_prng_io_out_19; // @[PRNG.scala 91:22]
  reg [31:0] txs; // @[TestHarness.scala 136:20]
  reg [31:0] flits; // @[TestHarness.scala 137:22]
  reg [31:0] tsc; // @[TestHarness.scala 141:20]
  wire [31:0] _tsc_T_1 = tsc + 32'h1; // @[TestHarness.scala 142:14]
  reg [10:0] idle_counter; // @[TestHarness.scala 144:29]
  wire [10:0] _idle_counter_T_1 = idle_counter + 11'h1; // @[TestHarness.scala 146:46]
  reg [127:0] rob_valids; // @[TestHarness.scala 156:27]
  wire [127:0] _T_5 = ~rob_valids; // @[TestHarness.scala 161:59]
  wire [6:0] _sels_0_T_128 = _T_5[126] ? 7'h7e : 7'h7f; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_129 = _T_5[125] ? 7'h7d : _sels_0_T_128; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_130 = _T_5[124] ? 7'h7c : _sels_0_T_129; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_131 = _T_5[123] ? 7'h7b : _sels_0_T_130; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_132 = _T_5[122] ? 7'h7a : _sels_0_T_131; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_133 = _T_5[121] ? 7'h79 : _sels_0_T_132; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_134 = _T_5[120] ? 7'h78 : _sels_0_T_133; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_135 = _T_5[119] ? 7'h77 : _sels_0_T_134; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_136 = _T_5[118] ? 7'h76 : _sels_0_T_135; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_137 = _T_5[117] ? 7'h75 : _sels_0_T_136; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_138 = _T_5[116] ? 7'h74 : _sels_0_T_137; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_139 = _T_5[115] ? 7'h73 : _sels_0_T_138; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_140 = _T_5[114] ? 7'h72 : _sels_0_T_139; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_141 = _T_5[113] ? 7'h71 : _sels_0_T_140; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_142 = _T_5[112] ? 7'h70 : _sels_0_T_141; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_143 = _T_5[111] ? 7'h6f : _sels_0_T_142; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_144 = _T_5[110] ? 7'h6e : _sels_0_T_143; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_145 = _T_5[109] ? 7'h6d : _sels_0_T_144; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_146 = _T_5[108] ? 7'h6c : _sels_0_T_145; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_147 = _T_5[107] ? 7'h6b : _sels_0_T_146; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_148 = _T_5[106] ? 7'h6a : _sels_0_T_147; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_149 = _T_5[105] ? 7'h69 : _sels_0_T_148; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_150 = _T_5[104] ? 7'h68 : _sels_0_T_149; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_151 = _T_5[103] ? 7'h67 : _sels_0_T_150; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_152 = _T_5[102] ? 7'h66 : _sels_0_T_151; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_153 = _T_5[101] ? 7'h65 : _sels_0_T_152; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_154 = _T_5[100] ? 7'h64 : _sels_0_T_153; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_155 = _T_5[99] ? 7'h63 : _sels_0_T_154; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_156 = _T_5[98] ? 7'h62 : _sels_0_T_155; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_157 = _T_5[97] ? 7'h61 : _sels_0_T_156; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_158 = _T_5[96] ? 7'h60 : _sels_0_T_157; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_159 = _T_5[95] ? 7'h5f : _sels_0_T_158; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_160 = _T_5[94] ? 7'h5e : _sels_0_T_159; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_161 = _T_5[93] ? 7'h5d : _sels_0_T_160; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_162 = _T_5[92] ? 7'h5c : _sels_0_T_161; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_163 = _T_5[91] ? 7'h5b : _sels_0_T_162; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_164 = _T_5[90] ? 7'h5a : _sels_0_T_163; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_165 = _T_5[89] ? 7'h59 : _sels_0_T_164; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_166 = _T_5[88] ? 7'h58 : _sels_0_T_165; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_167 = _T_5[87] ? 7'h57 : _sels_0_T_166; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_168 = _T_5[86] ? 7'h56 : _sels_0_T_167; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_169 = _T_5[85] ? 7'h55 : _sels_0_T_168; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_170 = _T_5[84] ? 7'h54 : _sels_0_T_169; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_171 = _T_5[83] ? 7'h53 : _sels_0_T_170; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_172 = _T_5[82] ? 7'h52 : _sels_0_T_171; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_173 = _T_5[81] ? 7'h51 : _sels_0_T_172; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_174 = _T_5[80] ? 7'h50 : _sels_0_T_173; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_175 = _T_5[79] ? 7'h4f : _sels_0_T_174; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_176 = _T_5[78] ? 7'h4e : _sels_0_T_175; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_177 = _T_5[77] ? 7'h4d : _sels_0_T_176; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_178 = _T_5[76] ? 7'h4c : _sels_0_T_177; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_179 = _T_5[75] ? 7'h4b : _sels_0_T_178; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_180 = _T_5[74] ? 7'h4a : _sels_0_T_179; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_181 = _T_5[73] ? 7'h49 : _sels_0_T_180; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_182 = _T_5[72] ? 7'h48 : _sels_0_T_181; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_183 = _T_5[71] ? 7'h47 : _sels_0_T_182; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_184 = _T_5[70] ? 7'h46 : _sels_0_T_183; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_185 = _T_5[69] ? 7'h45 : _sels_0_T_184; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_186 = _T_5[68] ? 7'h44 : _sels_0_T_185; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_187 = _T_5[67] ? 7'h43 : _sels_0_T_186; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_188 = _T_5[66] ? 7'h42 : _sels_0_T_187; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_189 = _T_5[65] ? 7'h41 : _sels_0_T_188; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_190 = _T_5[64] ? 7'h40 : _sels_0_T_189; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_191 = _T_5[63] ? 7'h3f : _sels_0_T_190; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_192 = _T_5[62] ? 7'h3e : _sels_0_T_191; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_193 = _T_5[61] ? 7'h3d : _sels_0_T_192; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_194 = _T_5[60] ? 7'h3c : _sels_0_T_193; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_195 = _T_5[59] ? 7'h3b : _sels_0_T_194; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_196 = _T_5[58] ? 7'h3a : _sels_0_T_195; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_197 = _T_5[57] ? 7'h39 : _sels_0_T_196; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_198 = _T_5[56] ? 7'h38 : _sels_0_T_197; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_199 = _T_5[55] ? 7'h37 : _sels_0_T_198; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_200 = _T_5[54] ? 7'h36 : _sels_0_T_199; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_201 = _T_5[53] ? 7'h35 : _sels_0_T_200; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_202 = _T_5[52] ? 7'h34 : _sels_0_T_201; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_203 = _T_5[51] ? 7'h33 : _sels_0_T_202; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_204 = _T_5[50] ? 7'h32 : _sels_0_T_203; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_205 = _T_5[49] ? 7'h31 : _sels_0_T_204; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_206 = _T_5[48] ? 7'h30 : _sels_0_T_205; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_207 = _T_5[47] ? 7'h2f : _sels_0_T_206; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_208 = _T_5[46] ? 7'h2e : _sels_0_T_207; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_209 = _T_5[45] ? 7'h2d : _sels_0_T_208; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_210 = _T_5[44] ? 7'h2c : _sels_0_T_209; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_211 = _T_5[43] ? 7'h2b : _sels_0_T_210; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_212 = _T_5[42] ? 7'h2a : _sels_0_T_211; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_213 = _T_5[41] ? 7'h29 : _sels_0_T_212; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_214 = _T_5[40] ? 7'h28 : _sels_0_T_213; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_215 = _T_5[39] ? 7'h27 : _sels_0_T_214; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_216 = _T_5[38] ? 7'h26 : _sels_0_T_215; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_217 = _T_5[37] ? 7'h25 : _sels_0_T_216; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_218 = _T_5[36] ? 7'h24 : _sels_0_T_217; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_219 = _T_5[35] ? 7'h23 : _sels_0_T_218; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_220 = _T_5[34] ? 7'h22 : _sels_0_T_219; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_221 = _T_5[33] ? 7'h21 : _sels_0_T_220; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_222 = _T_5[32] ? 7'h20 : _sels_0_T_221; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_223 = _T_5[31] ? 7'h1f : _sels_0_T_222; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_224 = _T_5[30] ? 7'h1e : _sels_0_T_223; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_225 = _T_5[29] ? 7'h1d : _sels_0_T_224; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_226 = _T_5[28] ? 7'h1c : _sels_0_T_225; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_227 = _T_5[27] ? 7'h1b : _sels_0_T_226; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_228 = _T_5[26] ? 7'h1a : _sels_0_T_227; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_229 = _T_5[25] ? 7'h19 : _sels_0_T_228; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_230 = _T_5[24] ? 7'h18 : _sels_0_T_229; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_231 = _T_5[23] ? 7'h17 : _sels_0_T_230; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_232 = _T_5[22] ? 7'h16 : _sels_0_T_231; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_233 = _T_5[21] ? 7'h15 : _sels_0_T_232; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_234 = _T_5[20] ? 7'h14 : _sels_0_T_233; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_235 = _T_5[19] ? 7'h13 : _sels_0_T_234; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_236 = _T_5[18] ? 7'h12 : _sels_0_T_235; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_237 = _T_5[17] ? 7'h11 : _sels_0_T_236; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_238 = _T_5[16] ? 7'h10 : _sels_0_T_237; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_239 = _T_5[15] ? 7'hf : _sels_0_T_238; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_240 = _T_5[14] ? 7'he : _sels_0_T_239; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_241 = _T_5[13] ? 7'hd : _sels_0_T_240; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_242 = _T_5[12] ? 7'hc : _sels_0_T_241; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_243 = _T_5[11] ? 7'hb : _sels_0_T_242; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_244 = _T_5[10] ? 7'ha : _sels_0_T_243; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_245 = _T_5[9] ? 7'h9 : _sels_0_T_244; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_246 = _T_5[8] ? 7'h8 : _sels_0_T_245; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_247 = _T_5[7] ? 7'h7 : _sels_0_T_246; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_248 = _T_5[6] ? 7'h6 : _sels_0_T_247; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_249 = _T_5[5] ? 7'h5 : _sels_0_T_248; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_250 = _T_5[4] ? 7'h4 : _sels_0_T_249; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_251 = _T_5[3] ? 7'h3 : _sels_0_T_250; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_252 = _T_5[2] ? 7'h2 : _sels_0_T_251; // @[Mux.scala 47:70]
  wire [6:0] _sels_0_T_253 = _T_5[1] ? 7'h1 : _sels_0_T_252; // @[Mux.scala 47:70]
  wire [6:0] rob_alloc_ids_0 = _T_5[0] ? 7'h0 : _sels_0_T_253; // @[Mux.scala 47:70]
  wire [127:0] _GEN_3073 = {{127'd0}, igen_io_fire}; // @[TestHarness.scala 187:45]
  wire [127:0] _T_26 = _GEN_3073 << rob_alloc_ids_0; // @[TestHarness.scala 187:45]
  wire [127:0] _T_6 = 128'h1 << rob_alloc_ids_0; // @[TestHarness.scala 31:27]
  wire [127:0] _T_7 = ~_T_6; // @[TestHarness.scala 31:21]
  wire [127:0] _T_8 = _T_5 & _T_7; // @[TestHarness.scala 31:19]
  wire [6:0] _sels_1_T_128 = _T_8[126] ? 7'h7e : 7'h7f; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_129 = _T_8[125] ? 7'h7d : _sels_1_T_128; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_130 = _T_8[124] ? 7'h7c : _sels_1_T_129; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_131 = _T_8[123] ? 7'h7b : _sels_1_T_130; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_132 = _T_8[122] ? 7'h7a : _sels_1_T_131; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_133 = _T_8[121] ? 7'h79 : _sels_1_T_132; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_134 = _T_8[120] ? 7'h78 : _sels_1_T_133; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_135 = _T_8[119] ? 7'h77 : _sels_1_T_134; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_136 = _T_8[118] ? 7'h76 : _sels_1_T_135; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_137 = _T_8[117] ? 7'h75 : _sels_1_T_136; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_138 = _T_8[116] ? 7'h74 : _sels_1_T_137; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_139 = _T_8[115] ? 7'h73 : _sels_1_T_138; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_140 = _T_8[114] ? 7'h72 : _sels_1_T_139; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_141 = _T_8[113] ? 7'h71 : _sels_1_T_140; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_142 = _T_8[112] ? 7'h70 : _sels_1_T_141; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_143 = _T_8[111] ? 7'h6f : _sels_1_T_142; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_144 = _T_8[110] ? 7'h6e : _sels_1_T_143; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_145 = _T_8[109] ? 7'h6d : _sels_1_T_144; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_146 = _T_8[108] ? 7'h6c : _sels_1_T_145; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_147 = _T_8[107] ? 7'h6b : _sels_1_T_146; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_148 = _T_8[106] ? 7'h6a : _sels_1_T_147; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_149 = _T_8[105] ? 7'h69 : _sels_1_T_148; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_150 = _T_8[104] ? 7'h68 : _sels_1_T_149; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_151 = _T_8[103] ? 7'h67 : _sels_1_T_150; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_152 = _T_8[102] ? 7'h66 : _sels_1_T_151; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_153 = _T_8[101] ? 7'h65 : _sels_1_T_152; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_154 = _T_8[100] ? 7'h64 : _sels_1_T_153; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_155 = _T_8[99] ? 7'h63 : _sels_1_T_154; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_156 = _T_8[98] ? 7'h62 : _sels_1_T_155; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_157 = _T_8[97] ? 7'h61 : _sels_1_T_156; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_158 = _T_8[96] ? 7'h60 : _sels_1_T_157; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_159 = _T_8[95] ? 7'h5f : _sels_1_T_158; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_160 = _T_8[94] ? 7'h5e : _sels_1_T_159; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_161 = _T_8[93] ? 7'h5d : _sels_1_T_160; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_162 = _T_8[92] ? 7'h5c : _sels_1_T_161; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_163 = _T_8[91] ? 7'h5b : _sels_1_T_162; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_164 = _T_8[90] ? 7'h5a : _sels_1_T_163; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_165 = _T_8[89] ? 7'h59 : _sels_1_T_164; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_166 = _T_8[88] ? 7'h58 : _sels_1_T_165; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_167 = _T_8[87] ? 7'h57 : _sels_1_T_166; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_168 = _T_8[86] ? 7'h56 : _sels_1_T_167; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_169 = _T_8[85] ? 7'h55 : _sels_1_T_168; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_170 = _T_8[84] ? 7'h54 : _sels_1_T_169; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_171 = _T_8[83] ? 7'h53 : _sels_1_T_170; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_172 = _T_8[82] ? 7'h52 : _sels_1_T_171; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_173 = _T_8[81] ? 7'h51 : _sels_1_T_172; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_174 = _T_8[80] ? 7'h50 : _sels_1_T_173; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_175 = _T_8[79] ? 7'h4f : _sels_1_T_174; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_176 = _T_8[78] ? 7'h4e : _sels_1_T_175; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_177 = _T_8[77] ? 7'h4d : _sels_1_T_176; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_178 = _T_8[76] ? 7'h4c : _sels_1_T_177; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_179 = _T_8[75] ? 7'h4b : _sels_1_T_178; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_180 = _T_8[74] ? 7'h4a : _sels_1_T_179; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_181 = _T_8[73] ? 7'h49 : _sels_1_T_180; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_182 = _T_8[72] ? 7'h48 : _sels_1_T_181; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_183 = _T_8[71] ? 7'h47 : _sels_1_T_182; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_184 = _T_8[70] ? 7'h46 : _sels_1_T_183; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_185 = _T_8[69] ? 7'h45 : _sels_1_T_184; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_186 = _T_8[68] ? 7'h44 : _sels_1_T_185; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_187 = _T_8[67] ? 7'h43 : _sels_1_T_186; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_188 = _T_8[66] ? 7'h42 : _sels_1_T_187; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_189 = _T_8[65] ? 7'h41 : _sels_1_T_188; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_190 = _T_8[64] ? 7'h40 : _sels_1_T_189; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_191 = _T_8[63] ? 7'h3f : _sels_1_T_190; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_192 = _T_8[62] ? 7'h3e : _sels_1_T_191; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_193 = _T_8[61] ? 7'h3d : _sels_1_T_192; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_194 = _T_8[60] ? 7'h3c : _sels_1_T_193; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_195 = _T_8[59] ? 7'h3b : _sels_1_T_194; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_196 = _T_8[58] ? 7'h3a : _sels_1_T_195; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_197 = _T_8[57] ? 7'h39 : _sels_1_T_196; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_198 = _T_8[56] ? 7'h38 : _sels_1_T_197; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_199 = _T_8[55] ? 7'h37 : _sels_1_T_198; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_200 = _T_8[54] ? 7'h36 : _sels_1_T_199; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_201 = _T_8[53] ? 7'h35 : _sels_1_T_200; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_202 = _T_8[52] ? 7'h34 : _sels_1_T_201; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_203 = _T_8[51] ? 7'h33 : _sels_1_T_202; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_204 = _T_8[50] ? 7'h32 : _sels_1_T_203; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_205 = _T_8[49] ? 7'h31 : _sels_1_T_204; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_206 = _T_8[48] ? 7'h30 : _sels_1_T_205; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_207 = _T_8[47] ? 7'h2f : _sels_1_T_206; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_208 = _T_8[46] ? 7'h2e : _sels_1_T_207; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_209 = _T_8[45] ? 7'h2d : _sels_1_T_208; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_210 = _T_8[44] ? 7'h2c : _sels_1_T_209; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_211 = _T_8[43] ? 7'h2b : _sels_1_T_210; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_212 = _T_8[42] ? 7'h2a : _sels_1_T_211; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_213 = _T_8[41] ? 7'h29 : _sels_1_T_212; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_214 = _T_8[40] ? 7'h28 : _sels_1_T_213; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_215 = _T_8[39] ? 7'h27 : _sels_1_T_214; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_216 = _T_8[38] ? 7'h26 : _sels_1_T_215; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_217 = _T_8[37] ? 7'h25 : _sels_1_T_216; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_218 = _T_8[36] ? 7'h24 : _sels_1_T_217; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_219 = _T_8[35] ? 7'h23 : _sels_1_T_218; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_220 = _T_8[34] ? 7'h22 : _sels_1_T_219; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_221 = _T_8[33] ? 7'h21 : _sels_1_T_220; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_222 = _T_8[32] ? 7'h20 : _sels_1_T_221; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_223 = _T_8[31] ? 7'h1f : _sels_1_T_222; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_224 = _T_8[30] ? 7'h1e : _sels_1_T_223; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_225 = _T_8[29] ? 7'h1d : _sels_1_T_224; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_226 = _T_8[28] ? 7'h1c : _sels_1_T_225; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_227 = _T_8[27] ? 7'h1b : _sels_1_T_226; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_228 = _T_8[26] ? 7'h1a : _sels_1_T_227; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_229 = _T_8[25] ? 7'h19 : _sels_1_T_228; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_230 = _T_8[24] ? 7'h18 : _sels_1_T_229; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_231 = _T_8[23] ? 7'h17 : _sels_1_T_230; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_232 = _T_8[22] ? 7'h16 : _sels_1_T_231; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_233 = _T_8[21] ? 7'h15 : _sels_1_T_232; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_234 = _T_8[20] ? 7'h14 : _sels_1_T_233; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_235 = _T_8[19] ? 7'h13 : _sels_1_T_234; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_236 = _T_8[18] ? 7'h12 : _sels_1_T_235; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_237 = _T_8[17] ? 7'h11 : _sels_1_T_236; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_238 = _T_8[16] ? 7'h10 : _sels_1_T_237; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_239 = _T_8[15] ? 7'hf : _sels_1_T_238; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_240 = _T_8[14] ? 7'he : _sels_1_T_239; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_241 = _T_8[13] ? 7'hd : _sels_1_T_240; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_242 = _T_8[12] ? 7'hc : _sels_1_T_241; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_243 = _T_8[11] ? 7'hb : _sels_1_T_242; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_244 = _T_8[10] ? 7'ha : _sels_1_T_243; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_245 = _T_8[9] ? 7'h9 : _sels_1_T_244; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_246 = _T_8[8] ? 7'h8 : _sels_1_T_245; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_247 = _T_8[7] ? 7'h7 : _sels_1_T_246; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_248 = _T_8[6] ? 7'h6 : _sels_1_T_247; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_249 = _T_8[5] ? 7'h5 : _sels_1_T_248; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_250 = _T_8[4] ? 7'h4 : _sels_1_T_249; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_251 = _T_8[3] ? 7'h3 : _sels_1_T_250; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_252 = _T_8[2] ? 7'h2 : _sels_1_T_251; // @[Mux.scala 47:70]
  wire [6:0] _sels_1_T_253 = _T_8[1] ? 7'h1 : _sels_1_T_252; // @[Mux.scala 47:70]
  wire [6:0] rob_alloc_ids_1 = _T_8[0] ? 7'h0 : _sels_1_T_253; // @[Mux.scala 47:70]
  wire [127:0] _GEN_3074 = {{127'd0}, igen_1_io_fire}; // @[TestHarness.scala 187:45]
  wire [127:0] _T_40 = _GEN_3074 << rob_alloc_ids_1; // @[TestHarness.scala 187:45]
  wire [127:0] rob_allocs = _T_26 | _T_40; // @[TestHarness.scala 187:29]
  wire  _T_84 = io_from_noc_0_flit_ready & io_from_noc_0_flit_valid; // @[Decoupled.scala 51:35]
  wire  _T_85 = _T_84 & io_from_noc_0_flit_bits_tail; // @[TestHarness.scala 218:45]
  wire [15:0] out_payload_rob_idx = io_from_noc_0_flit_bits_payload[31:16]; // @[TestHarness.scala 194:51]
  wire [65535:0] _GEN_3075 = {{65535'd0}, _T_85}; // @[TestHarness.scala 218:66]
  wire [65535:0] _T_86 = _GEN_3075 << out_payload_rob_idx; // @[TestHarness.scala 218:66]
  wire  _T_131 = io_from_noc_1_flit_ready & io_from_noc_1_flit_valid; // @[Decoupled.scala 51:35]
  wire  _T_132 = _T_131 & io_from_noc_1_flit_bits_tail; // @[TestHarness.scala 218:45]
  wire [15:0] out_payload_1_rob_idx = io_from_noc_1_flit_bits_payload[31:16]; // @[TestHarness.scala 194:51]
  wire [65535:0] _GEN_3076 = {{65535'd0}, _T_132}; // @[TestHarness.scala 218:66]
  wire [65535:0] _T_133 = _GEN_3076 << out_payload_1_rob_idx; // @[TestHarness.scala 218:66]
  wire [65535:0] rob_frees = _T_86 | _T_133; // @[TestHarness.scala 218:27]
  wire  idle = rob_allocs == 128'h0 & rob_frees == 65536'h0; // @[TestHarness.scala 223:30]
  wire  _T_3 = ~reset; // @[TestHarness.scala 148:9]
  reg [31:0] rob_payload_0_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_0_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_0_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_1_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_1_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_1_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_2_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_2_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_2_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_3_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_3_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_3_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_4_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_4_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_4_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_5_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_5_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_5_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_6_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_6_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_6_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_7_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_7_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_7_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_8_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_8_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_8_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_9_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_9_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_9_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_10_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_10_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_10_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_11_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_11_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_11_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_12_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_12_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_12_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_13_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_13_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_13_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_14_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_14_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_14_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_15_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_15_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_15_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_16_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_16_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_16_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_17_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_17_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_17_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_18_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_18_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_18_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_19_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_19_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_19_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_20_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_20_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_20_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_21_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_21_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_21_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_22_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_22_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_22_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_23_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_23_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_23_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_24_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_24_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_24_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_25_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_25_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_25_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_26_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_26_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_26_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_27_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_27_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_27_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_28_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_28_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_28_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_29_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_29_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_29_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_30_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_30_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_30_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_31_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_31_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_31_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_32_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_32_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_32_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_33_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_33_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_33_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_34_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_34_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_34_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_35_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_35_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_35_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_36_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_36_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_36_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_37_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_37_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_37_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_38_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_38_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_38_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_39_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_39_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_39_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_40_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_40_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_40_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_41_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_41_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_41_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_42_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_42_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_42_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_43_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_43_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_43_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_44_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_44_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_44_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_45_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_45_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_45_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_46_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_46_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_46_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_47_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_47_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_47_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_48_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_48_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_48_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_49_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_49_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_49_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_50_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_50_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_50_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_51_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_51_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_51_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_52_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_52_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_52_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_53_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_53_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_53_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_54_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_54_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_54_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_55_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_55_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_55_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_56_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_56_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_56_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_57_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_57_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_57_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_58_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_58_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_58_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_59_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_59_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_59_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_60_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_60_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_60_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_61_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_61_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_61_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_62_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_62_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_62_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_63_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_63_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_63_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_64_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_64_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_64_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_65_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_65_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_65_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_66_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_66_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_66_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_67_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_67_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_67_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_68_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_68_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_68_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_69_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_69_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_69_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_70_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_70_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_70_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_71_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_71_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_71_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_72_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_72_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_72_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_73_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_73_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_73_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_74_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_74_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_74_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_75_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_75_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_75_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_76_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_76_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_76_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_77_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_77_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_77_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_78_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_78_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_78_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_79_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_79_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_79_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_80_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_80_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_80_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_81_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_81_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_81_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_82_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_82_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_82_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_83_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_83_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_83_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_84_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_84_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_84_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_85_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_85_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_85_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_86_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_86_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_86_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_87_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_87_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_87_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_88_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_88_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_88_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_89_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_89_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_89_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_90_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_90_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_90_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_91_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_91_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_91_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_92_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_92_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_92_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_93_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_93_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_93_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_94_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_94_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_94_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_95_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_95_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_95_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_96_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_96_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_96_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_97_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_97_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_97_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_98_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_98_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_98_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_99_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_99_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_99_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_100_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_100_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_100_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_101_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_101_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_101_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_102_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_102_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_102_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_103_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_103_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_103_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_104_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_104_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_104_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_105_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_105_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_105_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_106_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_106_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_106_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_107_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_107_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_107_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_108_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_108_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_108_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_109_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_109_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_109_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_110_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_110_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_110_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_111_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_111_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_111_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_112_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_112_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_112_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_113_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_113_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_113_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_114_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_114_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_114_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_115_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_115_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_115_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_116_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_116_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_116_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_117_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_117_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_117_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_118_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_118_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_118_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_119_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_119_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_119_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_120_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_120_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_120_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_121_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_121_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_121_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_122_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_122_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_122_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_123_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_123_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_123_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_124_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_124_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_124_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_125_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_125_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_125_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_126_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_126_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_126_flits_fired; // @[TestHarness.scala 150:24]
  reg [31:0] rob_payload_127_tsc; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_127_rob_idx; // @[TestHarness.scala 150:24]
  reg [15:0] rob_payload_127_flits_fired; // @[TestHarness.scala 150:24]
  reg  rob_egress_id_0; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_1; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_2; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_3; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_4; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_5; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_6; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_7; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_8; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_9; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_10; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_11; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_12; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_13; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_14; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_15; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_16; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_17; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_18; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_19; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_20; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_21; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_22; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_23; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_24; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_25; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_26; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_27; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_28; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_29; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_30; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_31; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_32; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_33; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_34; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_35; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_36; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_37; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_38; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_39; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_40; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_41; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_42; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_43; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_44; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_45; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_46; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_47; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_48; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_49; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_50; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_51; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_52; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_53; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_54; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_55; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_56; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_57; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_58; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_59; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_60; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_61; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_62; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_63; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_64; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_65; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_66; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_67; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_68; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_69; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_70; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_71; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_72; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_73; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_74; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_75; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_76; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_77; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_78; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_79; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_80; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_81; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_82; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_83; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_84; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_85; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_86; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_87; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_88; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_89; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_90; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_91; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_92; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_93; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_94; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_95; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_96; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_97; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_98; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_99; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_100; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_101; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_102; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_103; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_104; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_105; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_106; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_107; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_108; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_109; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_110; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_111; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_112; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_113; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_114; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_115; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_116; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_117; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_118; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_119; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_120; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_121; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_122; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_123; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_124; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_125; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_126; // @[TestHarness.scala 151:26]
  reg  rob_egress_id_127; // @[TestHarness.scala 151:26]
  reg  rob_ingress_id_0; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_1; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_2; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_3; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_4; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_5; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_6; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_7; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_8; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_9; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_10; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_11; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_12; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_13; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_14; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_15; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_16; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_17; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_18; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_19; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_20; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_21; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_22; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_23; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_24; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_25; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_26; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_27; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_28; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_29; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_30; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_31; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_32; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_33; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_34; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_35; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_36; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_37; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_38; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_39; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_40; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_41; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_42; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_43; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_44; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_45; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_46; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_47; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_48; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_49; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_50; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_51; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_52; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_53; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_54; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_55; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_56; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_57; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_58; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_59; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_60; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_61; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_62; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_63; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_64; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_65; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_66; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_67; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_68; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_69; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_70; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_71; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_72; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_73; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_74; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_75; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_76; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_77; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_78; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_79; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_80; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_81; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_82; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_83; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_84; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_85; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_86; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_87; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_88; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_89; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_90; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_91; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_92; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_93; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_94; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_95; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_96; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_97; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_98; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_99; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_100; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_101; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_102; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_103; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_104; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_105; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_106; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_107; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_108; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_109; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_110; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_111; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_112; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_113; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_114; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_115; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_116; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_117; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_118; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_119; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_120; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_121; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_122; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_123; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_124; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_125; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_126; // @[TestHarness.scala 152:27]
  reg  rob_ingress_id_127; // @[TestHarness.scala 152:27]
  reg [3:0] rob_n_flits_0; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_1; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_2; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_3; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_4; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_5; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_6; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_7; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_8; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_9; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_10; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_11; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_12; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_13; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_14; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_15; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_16; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_17; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_18; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_19; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_20; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_21; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_22; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_23; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_24; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_25; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_26; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_27; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_28; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_29; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_30; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_31; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_32; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_33; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_34; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_35; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_36; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_37; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_38; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_39; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_40; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_41; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_42; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_43; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_44; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_45; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_46; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_47; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_48; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_49; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_50; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_51; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_52; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_53; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_54; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_55; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_56; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_57; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_58; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_59; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_60; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_61; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_62; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_63; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_64; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_65; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_66; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_67; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_68; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_69; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_70; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_71; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_72; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_73; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_74; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_75; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_76; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_77; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_78; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_79; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_80; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_81; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_82; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_83; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_84; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_85; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_86; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_87; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_88; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_89; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_90; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_91; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_92; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_93; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_94; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_95; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_96; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_97; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_98; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_99; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_100; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_101; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_102; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_103; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_104; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_105; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_106; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_107; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_108; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_109; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_110; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_111; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_112; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_113; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_114; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_115; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_116; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_117; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_118; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_119; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_120; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_121; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_122; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_123; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_124; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_125; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_126; // @[TestHarness.scala 153:24]
  reg [3:0] rob_n_flits_127; // @[TestHarness.scala 153:24]
  reg [3:0] rob_flits_returned_0; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_1; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_2; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_3; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_4; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_5; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_6; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_7; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_8; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_9; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_10; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_11; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_12; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_13; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_14; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_15; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_16; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_17; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_18; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_19; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_20; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_21; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_22; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_23; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_24; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_25; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_26; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_27; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_28; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_29; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_30; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_31; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_32; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_33; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_34; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_35; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_36; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_37; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_38; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_39; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_40; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_41; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_42; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_43; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_44; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_45; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_46; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_47; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_48; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_49; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_50; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_51; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_52; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_53; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_54; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_55; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_56; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_57; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_58; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_59; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_60; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_61; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_62; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_63; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_64; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_65; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_66; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_67; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_68; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_69; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_70; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_71; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_72; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_73; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_74; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_75; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_76; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_77; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_78; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_79; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_80; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_81; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_82; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_83; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_84; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_85; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_86; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_87; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_88; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_89; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_90; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_91; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_92; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_93; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_94; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_95; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_96; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_97; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_98; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_99; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_100; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_101; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_102; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_103; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_104; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_105; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_106; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_107; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_108; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_109; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_110; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_111; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_112; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_113; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_114; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_115; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_116; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_117; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_118; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_119; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_120; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_121; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_122; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_123; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_124; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_125; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_126; // @[TestHarness.scala 154:31]
  reg [3:0] rob_flits_returned_127; // @[TestHarness.scala 154:31]
  reg [63:0] rob_tscs_0; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_1; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_2; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_3; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_4; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_5; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_6; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_7; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_8; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_9; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_10; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_11; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_12; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_13; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_14; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_15; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_16; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_17; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_18; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_19; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_20; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_21; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_22; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_23; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_24; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_25; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_26; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_27; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_28; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_29; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_30; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_31; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_32; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_33; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_34; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_35; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_36; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_37; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_38; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_39; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_40; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_41; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_42; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_43; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_44; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_45; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_46; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_47; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_48; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_49; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_50; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_51; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_52; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_53; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_54; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_55; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_56; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_57; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_58; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_59; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_60; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_61; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_62; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_63; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_64; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_65; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_66; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_67; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_68; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_69; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_70; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_71; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_72; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_73; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_74; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_75; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_76; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_77; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_78; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_79; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_80; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_81; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_82; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_83; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_84; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_85; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_86; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_87; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_88; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_89; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_90; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_91; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_92; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_93; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_94; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_95; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_96; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_97; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_98; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_99; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_100; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_101; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_102; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_103; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_104; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_105; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_106; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_107; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_108; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_109; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_110; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_111; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_112; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_113; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_114; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_115; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_116; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_117; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_118; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_119; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_120; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_121; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_122; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_123; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_124; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_125; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_126; // @[TestHarness.scala 155:21]
  reg [63:0] rob_tscs_127; // @[TestHarness.scala 155:21]
  wire  rob_alloc_fires_0 = _T_5 != 128'h0; // @[TestHarness.scala 30:24]
  wire  rob_alloc_fires_1 = _T_8 != 128'h0; // @[TestHarness.scala 30:24]
  wire [127:0] _rob_alloc_avail_T = rob_valids >> rob_alloc_ids_0; // @[TestHarness.scala 162:61]
  wire  rob_alloc_avail_0 = ~_rob_alloc_avail_T[0]; // @[TestHarness.scala 162:50]
  wire [127:0] _rob_alloc_avail_T_2 = rob_valids >> rob_alloc_ids_1; // @[TestHarness.scala 162:61]
  wire  rob_alloc_avail_1 = ~_rob_alloc_avail_T_2[0]; // @[TestHarness.scala 162:50]
  wire  success = txs >= 32'hc350 & rob_valids == 128'h0; // @[TestHarness.scala 163:35]
  reg  io_success_REG; // @[TestHarness.scala 164:24]
  wire  _igen_io_rob_ready_T_1 = tsc >= 32'ha; // @[TestHarness.scala 175:11]
  wire  _igen_io_rob_ready_T_2 = rob_alloc_avail_0 & rob_alloc_fires_0 & _igen_io_rob_ready_T_1; // @[TestHarness.scala 174:72]
  wire [63:0] _rob_payload_WIRE_1 = igen_io_out_bits_payload; // @[TestHarness.scala 179:{72,72}]
  wire [31:0] _GEN_1 = 7'h0 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_0_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_2 = 7'h1 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_1_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_3 = 7'h2 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_2_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_4 = 7'h3 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_3_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_5 = 7'h4 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_4_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_6 = 7'h5 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_5_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_7 = 7'h6 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_6_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_8 = 7'h7 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_7_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_9 = 7'h8 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_8_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_10 = 7'h9 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_9_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_11 = 7'ha == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_10_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_12 = 7'hb == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_11_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_13 = 7'hc == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_12_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_14 = 7'hd == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_13_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_15 = 7'he == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_14_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_16 = 7'hf == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_15_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_17 = 7'h10 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_16_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_18 = 7'h11 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_17_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_19 = 7'h12 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_18_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_20 = 7'h13 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_19_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_21 = 7'h14 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_20_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_22 = 7'h15 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_21_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_23 = 7'h16 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_22_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_24 = 7'h17 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_23_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_25 = 7'h18 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_24_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_26 = 7'h19 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_25_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_27 = 7'h1a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_26_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_28 = 7'h1b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_27_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_29 = 7'h1c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_28_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_30 = 7'h1d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_29_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_31 = 7'h1e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_30_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_32 = 7'h1f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_31_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_33 = 7'h20 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_32_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_34 = 7'h21 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_33_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_35 = 7'h22 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_34_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_36 = 7'h23 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_35_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_37 = 7'h24 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_36_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_38 = 7'h25 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_37_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_39 = 7'h26 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_38_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_40 = 7'h27 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_39_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_41 = 7'h28 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_40_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_42 = 7'h29 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_41_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_43 = 7'h2a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_42_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_44 = 7'h2b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_43_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_45 = 7'h2c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_44_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_46 = 7'h2d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_45_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_47 = 7'h2e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_46_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_48 = 7'h2f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_47_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_49 = 7'h30 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_48_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_50 = 7'h31 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_49_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_51 = 7'h32 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_50_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_52 = 7'h33 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_51_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_53 = 7'h34 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_52_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_54 = 7'h35 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_53_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_55 = 7'h36 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_54_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_56 = 7'h37 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_55_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_57 = 7'h38 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_56_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_58 = 7'h39 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_57_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_59 = 7'h3a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_58_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_60 = 7'h3b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_59_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_61 = 7'h3c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_60_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_62 = 7'h3d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_61_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_63 = 7'h3e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_62_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_64 = 7'h3f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_63_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_65 = 7'h40 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_64_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_66 = 7'h41 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_65_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_67 = 7'h42 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_66_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_68 = 7'h43 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_67_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_69 = 7'h44 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_68_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_70 = 7'h45 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_69_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_71 = 7'h46 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_70_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_72 = 7'h47 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_71_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_73 = 7'h48 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_72_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_74 = 7'h49 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_73_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_75 = 7'h4a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_74_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_76 = 7'h4b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_75_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_77 = 7'h4c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_76_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_78 = 7'h4d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_77_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_79 = 7'h4e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_78_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_80 = 7'h4f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_79_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_81 = 7'h50 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_80_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_82 = 7'h51 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_81_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_83 = 7'h52 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_82_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_84 = 7'h53 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_83_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_85 = 7'h54 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_84_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_86 = 7'h55 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_85_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_87 = 7'h56 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_86_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_88 = 7'h57 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_87_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_89 = 7'h58 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_88_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_90 = 7'h59 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_89_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_91 = 7'h5a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_90_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_92 = 7'h5b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_91_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_93 = 7'h5c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_92_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_94 = 7'h5d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_93_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_95 = 7'h5e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_94_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_96 = 7'h5f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_95_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_97 = 7'h60 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_96_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_98 = 7'h61 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_97_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_99 = 7'h62 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_98_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_100 = 7'h63 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_99_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_101 = 7'h64 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_100_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_102 = 7'h65 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_101_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_103 = 7'h66 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_102_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_104 = 7'h67 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_103_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_105 = 7'h68 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_104_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_106 = 7'h69 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_105_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_107 = 7'h6a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_106_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_108 = 7'h6b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_107_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_109 = 7'h6c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_108_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_110 = 7'h6d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_109_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_111 = 7'h6e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_110_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_112 = 7'h6f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_111_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_113 = 7'h70 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_112_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_114 = 7'h71 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_113_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_115 = 7'h72 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_114_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_116 = 7'h73 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_115_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_117 = 7'h74 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_116_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_118 = 7'h75 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_117_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_119 = 7'h76 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_118_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_120 = 7'h77 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_119_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_121 = 7'h78 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_120_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_122 = 7'h79 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_121_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_123 = 7'h7a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_122_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_124 = 7'h7b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_123_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_125 = 7'h7c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_124_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_126 = 7'h7d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_125_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_127 = 7'h7e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_126_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [31:0] _GEN_128 = 7'h7f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[63:32] : rob_payload_127_tsc; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_129 = 7'h0 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_0_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_130 = 7'h1 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_1_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_131 = 7'h2 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_2_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_132 = 7'h3 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_3_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_133 = 7'h4 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_4_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_134 = 7'h5 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_5_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_135 = 7'h6 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_6_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_136 = 7'h7 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_7_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_137 = 7'h8 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_8_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_138 = 7'h9 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_9_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_139 = 7'ha == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_10_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_140 = 7'hb == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_11_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_141 = 7'hc == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_12_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_142 = 7'hd == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_13_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_143 = 7'he == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_14_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_144 = 7'hf == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_15_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_145 = 7'h10 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_16_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_146 = 7'h11 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_17_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_147 = 7'h12 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_18_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_148 = 7'h13 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_19_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_149 = 7'h14 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_20_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_150 = 7'h15 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_21_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_151 = 7'h16 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_22_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_152 = 7'h17 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_23_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_153 = 7'h18 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_24_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_154 = 7'h19 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_25_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_155 = 7'h1a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_26_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_156 = 7'h1b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_27_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_157 = 7'h1c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_28_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_158 = 7'h1d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_29_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_159 = 7'h1e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_30_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_160 = 7'h1f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_31_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_161 = 7'h20 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_32_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_162 = 7'h21 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_33_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_163 = 7'h22 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_34_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_164 = 7'h23 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_35_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_165 = 7'h24 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_36_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_166 = 7'h25 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_37_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_167 = 7'h26 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_38_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_168 = 7'h27 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_39_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_169 = 7'h28 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_40_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_170 = 7'h29 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_41_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_171 = 7'h2a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_42_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_172 = 7'h2b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_43_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_173 = 7'h2c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_44_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_174 = 7'h2d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_45_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_175 = 7'h2e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_46_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_176 = 7'h2f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_47_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_177 = 7'h30 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_48_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_178 = 7'h31 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_49_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_179 = 7'h32 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_50_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_180 = 7'h33 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_51_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_181 = 7'h34 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_52_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_182 = 7'h35 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_53_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_183 = 7'h36 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_54_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_184 = 7'h37 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_55_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_185 = 7'h38 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_56_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_186 = 7'h39 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_57_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_187 = 7'h3a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_58_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_188 = 7'h3b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_59_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_189 = 7'h3c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_60_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_190 = 7'h3d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_61_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_191 = 7'h3e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_62_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_192 = 7'h3f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_63_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_193 = 7'h40 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_64_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_194 = 7'h41 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_65_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_195 = 7'h42 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_66_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_196 = 7'h43 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_67_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_197 = 7'h44 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_68_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_198 = 7'h45 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_69_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_199 = 7'h46 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_70_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_200 = 7'h47 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_71_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_201 = 7'h48 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_72_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_202 = 7'h49 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_73_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_203 = 7'h4a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_74_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_204 = 7'h4b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_75_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_205 = 7'h4c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_76_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_206 = 7'h4d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_77_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_207 = 7'h4e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_78_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_208 = 7'h4f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_79_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_209 = 7'h50 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_80_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_210 = 7'h51 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_81_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_211 = 7'h52 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_82_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_212 = 7'h53 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_83_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_213 = 7'h54 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_84_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_214 = 7'h55 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_85_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_215 = 7'h56 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_86_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_216 = 7'h57 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_87_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_217 = 7'h58 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_88_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_218 = 7'h59 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_89_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_219 = 7'h5a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_90_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_220 = 7'h5b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_91_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_221 = 7'h5c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_92_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_222 = 7'h5d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_93_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_223 = 7'h5e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_94_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_224 = 7'h5f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_95_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_225 = 7'h60 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_96_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_226 = 7'h61 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_97_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_227 = 7'h62 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_98_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_228 = 7'h63 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_99_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_229 = 7'h64 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_100_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_230 = 7'h65 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_101_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_231 = 7'h66 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_102_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_232 = 7'h67 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_103_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_233 = 7'h68 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_104_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_234 = 7'h69 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_105_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_235 = 7'h6a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_106_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_236 = 7'h6b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_107_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_237 = 7'h6c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_108_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_238 = 7'h6d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_109_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_239 = 7'h6e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_110_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_240 = 7'h6f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_111_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_241 = 7'h70 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_112_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_242 = 7'h71 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_113_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_243 = 7'h72 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_114_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_244 = 7'h73 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_115_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_245 = 7'h74 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_116_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_246 = 7'h75 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_117_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_247 = 7'h76 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_118_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_248 = 7'h77 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_119_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_249 = 7'h78 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_120_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_250 = 7'h79 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_121_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_251 = 7'h7a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_122_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_252 = 7'h7b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_123_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_253 = 7'h7c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_124_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_254 = 7'h7d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_125_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_255 = 7'h7e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_126_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_256 = 7'h7f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[31:16] : rob_payload_127_rob_idx; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_257 = 7'h0 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_0_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_258 = 7'h1 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_1_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_259 = 7'h2 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_2_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_260 = 7'h3 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_3_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_261 = 7'h4 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_4_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_262 = 7'h5 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_5_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_263 = 7'h6 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_6_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_264 = 7'h7 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_7_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_265 = 7'h8 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_8_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_266 = 7'h9 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_9_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_267 = 7'ha == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_10_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_268 = 7'hb == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_11_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_269 = 7'hc == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_12_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_270 = 7'hd == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_13_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_271 = 7'he == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_14_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_272 = 7'hf == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_15_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_273 = 7'h10 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_16_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_274 = 7'h11 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_17_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_275 = 7'h12 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_18_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_276 = 7'h13 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_19_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_277 = 7'h14 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_20_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_278 = 7'h15 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_21_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_279 = 7'h16 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_22_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_280 = 7'h17 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_23_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_281 = 7'h18 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_24_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_282 = 7'h19 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_25_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_283 = 7'h1a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_26_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_284 = 7'h1b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_27_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_285 = 7'h1c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_28_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_286 = 7'h1d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_29_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_287 = 7'h1e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_30_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_288 = 7'h1f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_31_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_289 = 7'h20 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_32_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_290 = 7'h21 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_33_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_291 = 7'h22 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_34_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_292 = 7'h23 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_35_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_293 = 7'h24 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_36_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_294 = 7'h25 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_37_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_295 = 7'h26 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_38_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_296 = 7'h27 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_39_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_297 = 7'h28 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_40_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_298 = 7'h29 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_41_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_299 = 7'h2a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_42_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_300 = 7'h2b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_43_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_301 = 7'h2c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_44_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_302 = 7'h2d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_45_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_303 = 7'h2e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_46_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_304 = 7'h2f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_47_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_305 = 7'h30 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_48_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_306 = 7'h31 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_49_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_307 = 7'h32 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_50_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_308 = 7'h33 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_51_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_309 = 7'h34 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_52_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_310 = 7'h35 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_53_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_311 = 7'h36 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_54_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_312 = 7'h37 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_55_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_313 = 7'h38 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_56_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_314 = 7'h39 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_57_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_315 = 7'h3a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_58_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_316 = 7'h3b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_59_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_317 = 7'h3c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_60_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_318 = 7'h3d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_61_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_319 = 7'h3e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_62_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_320 = 7'h3f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_63_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_321 = 7'h40 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_64_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_322 = 7'h41 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_65_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_323 = 7'h42 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_66_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_324 = 7'h43 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_67_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_325 = 7'h44 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_68_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_326 = 7'h45 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_69_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_327 = 7'h46 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_70_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_328 = 7'h47 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_71_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_329 = 7'h48 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_72_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_330 = 7'h49 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_73_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_331 = 7'h4a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_74_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_332 = 7'h4b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_75_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_333 = 7'h4c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_76_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_334 = 7'h4d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_77_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_335 = 7'h4e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_78_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_336 = 7'h4f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_79_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_337 = 7'h50 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_80_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_338 = 7'h51 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_81_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_339 = 7'h52 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_82_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_340 = 7'h53 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_83_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_341 = 7'h54 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_84_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_342 = 7'h55 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_85_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_343 = 7'h56 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_86_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_344 = 7'h57 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_87_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_345 = 7'h58 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_88_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_346 = 7'h59 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_89_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_347 = 7'h5a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_90_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_348 = 7'h5b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_91_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_349 = 7'h5c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_92_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_350 = 7'h5d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_93_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_351 = 7'h5e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_94_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_352 = 7'h5f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_95_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_353 = 7'h60 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_96_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_354 = 7'h61 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_97_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_355 = 7'h62 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_98_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_356 = 7'h63 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_99_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_357 = 7'h64 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_100_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_358 = 7'h65 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_101_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_359 = 7'h66 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_102_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_360 = 7'h67 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_103_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_361 = 7'h68 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_104_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_362 = 7'h69 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_105_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_363 = 7'h6a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_106_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_364 = 7'h6b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_107_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_365 = 7'h6c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_108_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_366 = 7'h6d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_109_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_367 = 7'h6e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_110_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_368 = 7'h6f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_111_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_369 = 7'h70 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_112_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_370 = 7'h71 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_113_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_371 = 7'h72 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_114_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_372 = 7'h73 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_115_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_373 = 7'h74 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_116_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_374 = 7'h75 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_117_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_375 = 7'h76 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_118_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_376 = 7'h77 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_119_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_377 = 7'h78 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_120_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_378 = 7'h79 == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_121_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_379 = 7'h7a == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_122_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_380 = 7'h7b == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_123_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_381 = 7'h7c == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_124_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_382 = 7'h7d == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_125_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_383 = 7'h7e == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_126_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire [15:0] _GEN_384 = 7'h7f == rob_alloc_ids_0 ? _rob_payload_WIRE_1[15:0] : rob_payload_127_flits_fired; // @[TestHarness.scala 150:24 179:{36,36}]
  wire  _GEN_385 = 7'h0 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_0; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_386 = 7'h1 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_1; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_387 = 7'h2 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_2; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_388 = 7'h3 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_3; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_389 = 7'h4 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_4; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_390 = 7'h5 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_5; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_391 = 7'h6 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_6; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_392 = 7'h7 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_7; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_393 = 7'h8 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_8; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_394 = 7'h9 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_9; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_395 = 7'ha == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_10; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_396 = 7'hb == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_11; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_397 = 7'hc == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_12; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_398 = 7'hd == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_13; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_399 = 7'he == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_14; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_400 = 7'hf == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_15; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_401 = 7'h10 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_16; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_402 = 7'h11 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_17; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_403 = 7'h12 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_18; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_404 = 7'h13 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_19; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_405 = 7'h14 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_20; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_406 = 7'h15 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_21; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_407 = 7'h16 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_22; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_408 = 7'h17 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_23; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_409 = 7'h18 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_24; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_410 = 7'h19 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_25; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_411 = 7'h1a == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_26; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_412 = 7'h1b == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_27; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_413 = 7'h1c == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_28; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_414 = 7'h1d == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_29; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_415 = 7'h1e == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_30; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_416 = 7'h1f == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_31; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_417 = 7'h20 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_32; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_418 = 7'h21 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_33; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_419 = 7'h22 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_34; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_420 = 7'h23 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_35; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_421 = 7'h24 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_36; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_422 = 7'h25 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_37; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_423 = 7'h26 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_38; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_424 = 7'h27 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_39; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_425 = 7'h28 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_40; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_426 = 7'h29 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_41; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_427 = 7'h2a == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_42; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_428 = 7'h2b == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_43; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_429 = 7'h2c == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_44; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_430 = 7'h2d == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_45; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_431 = 7'h2e == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_46; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_432 = 7'h2f == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_47; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_433 = 7'h30 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_48; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_434 = 7'h31 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_49; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_435 = 7'h32 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_50; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_436 = 7'h33 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_51; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_437 = 7'h34 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_52; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_438 = 7'h35 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_53; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_439 = 7'h36 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_54; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_440 = 7'h37 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_55; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_441 = 7'h38 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_56; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_442 = 7'h39 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_57; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_443 = 7'h3a == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_58; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_444 = 7'h3b == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_59; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_445 = 7'h3c == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_60; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_446 = 7'h3d == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_61; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_447 = 7'h3e == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_62; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_448 = 7'h3f == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_63; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_449 = 7'h40 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_64; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_450 = 7'h41 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_65; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_451 = 7'h42 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_66; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_452 = 7'h43 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_67; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_453 = 7'h44 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_68; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_454 = 7'h45 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_69; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_455 = 7'h46 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_70; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_456 = 7'h47 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_71; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_457 = 7'h48 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_72; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_458 = 7'h49 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_73; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_459 = 7'h4a == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_74; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_460 = 7'h4b == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_75; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_461 = 7'h4c == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_76; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_462 = 7'h4d == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_77; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_463 = 7'h4e == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_78; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_464 = 7'h4f == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_79; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_465 = 7'h50 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_80; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_466 = 7'h51 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_81; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_467 = 7'h52 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_82; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_468 = 7'h53 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_83; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_469 = 7'h54 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_84; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_470 = 7'h55 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_85; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_471 = 7'h56 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_86; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_472 = 7'h57 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_87; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_473 = 7'h58 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_88; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_474 = 7'h59 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_89; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_475 = 7'h5a == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_90; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_476 = 7'h5b == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_91; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_477 = 7'h5c == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_92; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_478 = 7'h5d == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_93; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_479 = 7'h5e == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_94; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_480 = 7'h5f == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_95; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_481 = 7'h60 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_96; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_482 = 7'h61 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_97; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_483 = 7'h62 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_98; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_484 = 7'h63 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_99; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_485 = 7'h64 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_100; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_486 = 7'h65 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_101; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_487 = 7'h66 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_102; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_488 = 7'h67 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_103; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_489 = 7'h68 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_104; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_490 = 7'h69 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_105; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_491 = 7'h6a == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_106; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_492 = 7'h6b == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_107; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_493 = 7'h6c == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_108; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_494 = 7'h6d == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_109; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_495 = 7'h6e == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_110; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_496 = 7'h6f == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_111; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_497 = 7'h70 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_112; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_498 = 7'h71 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_113; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_499 = 7'h72 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_114; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_500 = 7'h73 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_115; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_501 = 7'h74 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_116; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_502 = 7'h75 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_117; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_503 = 7'h76 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_118; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_504 = 7'h77 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_119; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_505 = 7'h78 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_120; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_506 = 7'h79 == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_121; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_507 = 7'h7a == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_122; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_508 = 7'h7b == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_123; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_509 = 7'h7c == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_124; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_510 = 7'h7d == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_125; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_511 = 7'h7e == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_126; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_512 = 7'h7f == rob_alloc_ids_0 ? igen_io_out_bits_egress_id : rob_egress_id_127; // @[TestHarness.scala 151:26 180:{36,36}]
  wire  _GEN_513 = 7'h0 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_0; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_514 = 7'h1 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_1; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_515 = 7'h2 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_2; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_516 = 7'h3 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_3; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_517 = 7'h4 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_4; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_518 = 7'h5 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_5; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_519 = 7'h6 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_6; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_520 = 7'h7 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_7; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_521 = 7'h8 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_8; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_522 = 7'h9 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_9; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_523 = 7'ha == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_10; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_524 = 7'hb == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_11; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_525 = 7'hc == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_12; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_526 = 7'hd == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_13; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_527 = 7'he == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_14; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_528 = 7'hf == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_15; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_529 = 7'h10 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_16; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_530 = 7'h11 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_17; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_531 = 7'h12 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_18; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_532 = 7'h13 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_19; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_533 = 7'h14 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_20; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_534 = 7'h15 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_21; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_535 = 7'h16 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_22; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_536 = 7'h17 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_23; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_537 = 7'h18 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_24; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_538 = 7'h19 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_25; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_539 = 7'h1a == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_26; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_540 = 7'h1b == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_27; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_541 = 7'h1c == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_28; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_542 = 7'h1d == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_29; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_543 = 7'h1e == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_30; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_544 = 7'h1f == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_31; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_545 = 7'h20 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_32; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_546 = 7'h21 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_33; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_547 = 7'h22 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_34; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_548 = 7'h23 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_35; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_549 = 7'h24 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_36; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_550 = 7'h25 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_37; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_551 = 7'h26 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_38; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_552 = 7'h27 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_39; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_553 = 7'h28 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_40; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_554 = 7'h29 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_41; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_555 = 7'h2a == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_42; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_556 = 7'h2b == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_43; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_557 = 7'h2c == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_44; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_558 = 7'h2d == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_45; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_559 = 7'h2e == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_46; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_560 = 7'h2f == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_47; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_561 = 7'h30 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_48; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_562 = 7'h31 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_49; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_563 = 7'h32 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_50; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_564 = 7'h33 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_51; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_565 = 7'h34 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_52; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_566 = 7'h35 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_53; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_567 = 7'h36 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_54; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_568 = 7'h37 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_55; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_569 = 7'h38 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_56; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_570 = 7'h39 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_57; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_571 = 7'h3a == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_58; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_572 = 7'h3b == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_59; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_573 = 7'h3c == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_60; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_574 = 7'h3d == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_61; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_575 = 7'h3e == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_62; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_576 = 7'h3f == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_63; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_577 = 7'h40 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_64; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_578 = 7'h41 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_65; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_579 = 7'h42 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_66; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_580 = 7'h43 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_67; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_581 = 7'h44 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_68; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_582 = 7'h45 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_69; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_583 = 7'h46 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_70; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_584 = 7'h47 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_71; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_585 = 7'h48 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_72; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_586 = 7'h49 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_73; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_587 = 7'h4a == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_74; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_588 = 7'h4b == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_75; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_589 = 7'h4c == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_76; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_590 = 7'h4d == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_77; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_591 = 7'h4e == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_78; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_592 = 7'h4f == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_79; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_593 = 7'h50 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_80; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_594 = 7'h51 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_81; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_595 = 7'h52 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_82; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_596 = 7'h53 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_83; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_597 = 7'h54 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_84; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_598 = 7'h55 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_85; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_599 = 7'h56 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_86; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_600 = 7'h57 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_87; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_601 = 7'h58 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_88; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_602 = 7'h59 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_89; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_603 = 7'h5a == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_90; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_604 = 7'h5b == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_91; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_605 = 7'h5c == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_92; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_606 = 7'h5d == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_93; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_607 = 7'h5e == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_94; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_608 = 7'h5f == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_95; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_609 = 7'h60 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_96; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_610 = 7'h61 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_97; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_611 = 7'h62 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_98; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_612 = 7'h63 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_99; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_613 = 7'h64 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_100; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_614 = 7'h65 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_101; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_615 = 7'h66 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_102; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_616 = 7'h67 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_103; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_617 = 7'h68 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_104; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_618 = 7'h69 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_105; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_619 = 7'h6a == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_106; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_620 = 7'h6b == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_107; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_621 = 7'h6c == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_108; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_622 = 7'h6d == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_109; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_623 = 7'h6e == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_110; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_624 = 7'h6f == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_111; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_625 = 7'h70 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_112; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_626 = 7'h71 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_113; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_627 = 7'h72 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_114; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_628 = 7'h73 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_115; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_629 = 7'h74 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_116; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_630 = 7'h75 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_117; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_631 = 7'h76 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_118; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_632 = 7'h77 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_119; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_633 = 7'h78 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_120; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_634 = 7'h79 == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_121; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_635 = 7'h7a == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_122; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_636 = 7'h7b == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_123; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_637 = 7'h7c == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_124; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_638 = 7'h7d == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_125; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_639 = 7'h7e == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_126; // @[TestHarness.scala 152:27 181:{36,36}]
  wire  _GEN_640 = 7'h7f == rob_alloc_ids_0 ? 1'h0 : rob_ingress_id_127; // @[TestHarness.scala 152:27 181:{36,36}]
  wire [3:0] _rob_n_flits_T_21 = igen_io_n_flits; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_641 = 7'h0 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_0; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_642 = 7'h1 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_1; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_643 = 7'h2 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_2; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_644 = 7'h3 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_3; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_645 = 7'h4 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_4; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_646 = 7'h5 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_5; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_647 = 7'h6 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_6; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_648 = 7'h7 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_7; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_649 = 7'h8 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_8; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_650 = 7'h9 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_9; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_651 = 7'ha == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_10; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_652 = 7'hb == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_11; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_653 = 7'hc == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_12; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_654 = 7'hd == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_13; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_655 = 7'he == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_14; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_656 = 7'hf == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_15; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_657 = 7'h10 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_16; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_658 = 7'h11 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_17; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_659 = 7'h12 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_18; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_660 = 7'h13 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_19; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_661 = 7'h14 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_20; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_662 = 7'h15 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_21; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_663 = 7'h16 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_22; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_664 = 7'h17 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_23; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_665 = 7'h18 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_24; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_666 = 7'h19 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_25; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_667 = 7'h1a == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_26; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_668 = 7'h1b == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_27; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_669 = 7'h1c == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_28; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_670 = 7'h1d == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_29; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_671 = 7'h1e == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_30; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_672 = 7'h1f == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_31; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_673 = 7'h20 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_32; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_674 = 7'h21 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_33; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_675 = 7'h22 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_34; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_676 = 7'h23 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_35; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_677 = 7'h24 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_36; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_678 = 7'h25 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_37; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_679 = 7'h26 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_38; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_680 = 7'h27 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_39; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_681 = 7'h28 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_40; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_682 = 7'h29 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_41; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_683 = 7'h2a == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_42; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_684 = 7'h2b == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_43; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_685 = 7'h2c == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_44; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_686 = 7'h2d == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_45; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_687 = 7'h2e == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_46; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_688 = 7'h2f == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_47; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_689 = 7'h30 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_48; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_690 = 7'h31 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_49; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_691 = 7'h32 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_50; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_692 = 7'h33 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_51; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_693 = 7'h34 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_52; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_694 = 7'h35 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_53; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_695 = 7'h36 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_54; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_696 = 7'h37 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_55; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_697 = 7'h38 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_56; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_698 = 7'h39 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_57; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_699 = 7'h3a == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_58; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_700 = 7'h3b == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_59; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_701 = 7'h3c == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_60; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_702 = 7'h3d == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_61; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_703 = 7'h3e == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_62; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_704 = 7'h3f == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_63; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_705 = 7'h40 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_64; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_706 = 7'h41 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_65; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_707 = 7'h42 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_66; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_708 = 7'h43 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_67; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_709 = 7'h44 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_68; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_710 = 7'h45 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_69; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_711 = 7'h46 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_70; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_712 = 7'h47 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_71; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_713 = 7'h48 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_72; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_714 = 7'h49 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_73; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_715 = 7'h4a == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_74; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_716 = 7'h4b == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_75; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_717 = 7'h4c == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_76; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_718 = 7'h4d == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_77; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_719 = 7'h4e == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_78; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_720 = 7'h4f == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_79; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_721 = 7'h50 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_80; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_722 = 7'h51 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_81; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_723 = 7'h52 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_82; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_724 = 7'h53 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_83; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_725 = 7'h54 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_84; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_726 = 7'h55 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_85; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_727 = 7'h56 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_86; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_728 = 7'h57 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_87; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_729 = 7'h58 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_88; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_730 = 7'h59 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_89; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_731 = 7'h5a == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_90; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_732 = 7'h5b == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_91; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_733 = 7'h5c == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_92; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_734 = 7'h5d == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_93; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_735 = 7'h5e == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_94; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_736 = 7'h5f == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_95; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_737 = 7'h60 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_96; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_738 = 7'h61 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_97; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_739 = 7'h62 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_98; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_740 = 7'h63 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_99; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_741 = 7'h64 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_100; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_742 = 7'h65 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_101; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_743 = 7'h66 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_102; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_744 = 7'h67 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_103; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_745 = 7'h68 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_104; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_746 = 7'h69 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_105; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_747 = 7'h6a == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_106; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_748 = 7'h6b == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_107; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_749 = 7'h6c == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_108; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_750 = 7'h6d == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_109; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_751 = 7'h6e == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_110; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_752 = 7'h6f == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_111; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_753 = 7'h70 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_112; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_754 = 7'h71 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_113; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_755 = 7'h72 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_114; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_756 = 7'h73 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_115; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_757 = 7'h74 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_116; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_758 = 7'h75 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_117; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_759 = 7'h76 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_118; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_760 = 7'h77 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_119; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_761 = 7'h78 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_120; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_762 = 7'h79 == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_121; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_763 = 7'h7a == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_122; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_764 = 7'h7b == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_123; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_765 = 7'h7c == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_124; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_766 = 7'h7d == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_125; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_767 = 7'h7e == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_126; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_768 = 7'h7f == rob_alloc_ids_0 ? _rob_n_flits_T_21 : rob_n_flits_127; // @[TestHarness.scala 153:24 182:{36,36}]
  wire [3:0] _GEN_769 = 7'h0 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_0; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_770 = 7'h1 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_1; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_771 = 7'h2 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_2; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_772 = 7'h3 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_3; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_773 = 7'h4 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_4; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_774 = 7'h5 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_5; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_775 = 7'h6 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_6; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_776 = 7'h7 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_7; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_777 = 7'h8 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_8; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_778 = 7'h9 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_9; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_779 = 7'ha == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_10; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_780 = 7'hb == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_11; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_781 = 7'hc == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_12; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_782 = 7'hd == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_13; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_783 = 7'he == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_14; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_784 = 7'hf == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_15; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_785 = 7'h10 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_16; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_786 = 7'h11 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_17; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_787 = 7'h12 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_18; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_788 = 7'h13 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_19; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_789 = 7'h14 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_20; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_790 = 7'h15 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_21; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_791 = 7'h16 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_22; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_792 = 7'h17 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_23; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_793 = 7'h18 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_24; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_794 = 7'h19 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_25; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_795 = 7'h1a == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_26; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_796 = 7'h1b == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_27; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_797 = 7'h1c == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_28; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_798 = 7'h1d == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_29; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_799 = 7'h1e == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_30; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_800 = 7'h1f == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_31; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_801 = 7'h20 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_32; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_802 = 7'h21 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_33; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_803 = 7'h22 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_34; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_804 = 7'h23 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_35; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_805 = 7'h24 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_36; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_806 = 7'h25 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_37; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_807 = 7'h26 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_38; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_808 = 7'h27 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_39; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_809 = 7'h28 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_40; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_810 = 7'h29 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_41; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_811 = 7'h2a == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_42; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_812 = 7'h2b == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_43; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_813 = 7'h2c == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_44; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_814 = 7'h2d == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_45; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_815 = 7'h2e == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_46; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_816 = 7'h2f == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_47; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_817 = 7'h30 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_48; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_818 = 7'h31 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_49; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_819 = 7'h32 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_50; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_820 = 7'h33 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_51; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_821 = 7'h34 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_52; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_822 = 7'h35 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_53; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_823 = 7'h36 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_54; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_824 = 7'h37 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_55; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_825 = 7'h38 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_56; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_826 = 7'h39 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_57; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_827 = 7'h3a == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_58; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_828 = 7'h3b == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_59; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_829 = 7'h3c == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_60; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_830 = 7'h3d == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_61; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_831 = 7'h3e == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_62; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_832 = 7'h3f == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_63; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_833 = 7'h40 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_64; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_834 = 7'h41 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_65; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_835 = 7'h42 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_66; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_836 = 7'h43 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_67; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_837 = 7'h44 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_68; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_838 = 7'h45 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_69; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_839 = 7'h46 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_70; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_840 = 7'h47 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_71; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_841 = 7'h48 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_72; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_842 = 7'h49 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_73; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_843 = 7'h4a == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_74; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_844 = 7'h4b == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_75; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_845 = 7'h4c == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_76; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_846 = 7'h4d == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_77; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_847 = 7'h4e == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_78; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_848 = 7'h4f == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_79; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_849 = 7'h50 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_80; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_850 = 7'h51 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_81; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_851 = 7'h52 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_82; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_852 = 7'h53 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_83; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_853 = 7'h54 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_84; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_854 = 7'h55 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_85; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_855 = 7'h56 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_86; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_856 = 7'h57 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_87; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_857 = 7'h58 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_88; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_858 = 7'h59 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_89; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_859 = 7'h5a == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_90; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_860 = 7'h5b == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_91; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_861 = 7'h5c == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_92; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_862 = 7'h5d == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_93; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_863 = 7'h5e == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_94; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_864 = 7'h5f == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_95; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_865 = 7'h60 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_96; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_866 = 7'h61 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_97; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_867 = 7'h62 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_98; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_868 = 7'h63 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_99; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_869 = 7'h64 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_100; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_870 = 7'h65 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_101; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_871 = 7'h66 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_102; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_872 = 7'h67 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_103; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_873 = 7'h68 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_104; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_874 = 7'h69 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_105; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_875 = 7'h6a == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_106; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_876 = 7'h6b == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_107; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_877 = 7'h6c == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_108; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_878 = 7'h6d == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_109; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_879 = 7'h6e == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_110; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_880 = 7'h6f == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_111; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_881 = 7'h70 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_112; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_882 = 7'h71 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_113; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_883 = 7'h72 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_114; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_884 = 7'h73 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_115; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_885 = 7'h74 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_116; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_886 = 7'h75 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_117; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_887 = 7'h76 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_118; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_888 = 7'h77 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_119; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_889 = 7'h78 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_120; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_890 = 7'h79 == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_121; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_891 = 7'h7a == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_122; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_892 = 7'h7b == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_123; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_893 = 7'h7c == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_124; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_894 = 7'h7d == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_125; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_895 = 7'h7e == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_126; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [3:0] _GEN_896 = 7'h7f == rob_alloc_ids_0 ? 4'h0 : rob_flits_returned_127; // @[TestHarness.scala 154:31 183:{36,36}]
  wire [63:0] _rob_tscs_T_25 = {{32'd0}, tsc}; // @[TestHarness.scala 184:{36,36}]
  wire [63:0] _GEN_897 = 7'h0 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_0; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_898 = 7'h1 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_1; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_899 = 7'h2 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_2; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_900 = 7'h3 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_3; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_901 = 7'h4 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_4; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_902 = 7'h5 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_5; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_903 = 7'h6 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_6; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_904 = 7'h7 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_7; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_905 = 7'h8 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_8; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_906 = 7'h9 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_9; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_907 = 7'ha == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_10; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_908 = 7'hb == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_11; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_909 = 7'hc == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_12; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_910 = 7'hd == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_13; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_911 = 7'he == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_14; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_912 = 7'hf == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_15; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_913 = 7'h10 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_16; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_914 = 7'h11 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_17; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_915 = 7'h12 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_18; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_916 = 7'h13 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_19; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_917 = 7'h14 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_20; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_918 = 7'h15 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_21; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_919 = 7'h16 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_22; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_920 = 7'h17 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_23; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_921 = 7'h18 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_24; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_922 = 7'h19 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_25; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_923 = 7'h1a == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_26; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_924 = 7'h1b == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_27; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_925 = 7'h1c == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_28; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_926 = 7'h1d == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_29; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_927 = 7'h1e == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_30; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_928 = 7'h1f == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_31; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_929 = 7'h20 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_32; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_930 = 7'h21 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_33; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_931 = 7'h22 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_34; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_932 = 7'h23 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_35; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_933 = 7'h24 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_36; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_934 = 7'h25 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_37; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_935 = 7'h26 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_38; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_936 = 7'h27 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_39; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_937 = 7'h28 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_40; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_938 = 7'h29 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_41; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_939 = 7'h2a == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_42; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_940 = 7'h2b == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_43; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_941 = 7'h2c == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_44; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_942 = 7'h2d == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_45; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_943 = 7'h2e == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_46; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_944 = 7'h2f == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_47; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_945 = 7'h30 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_48; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_946 = 7'h31 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_49; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_947 = 7'h32 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_50; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_948 = 7'h33 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_51; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_949 = 7'h34 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_52; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_950 = 7'h35 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_53; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_951 = 7'h36 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_54; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_952 = 7'h37 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_55; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_953 = 7'h38 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_56; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_954 = 7'h39 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_57; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_955 = 7'h3a == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_58; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_956 = 7'h3b == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_59; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_957 = 7'h3c == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_60; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_958 = 7'h3d == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_61; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_959 = 7'h3e == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_62; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_960 = 7'h3f == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_63; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_961 = 7'h40 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_64; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_962 = 7'h41 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_65; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_963 = 7'h42 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_66; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_964 = 7'h43 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_67; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_965 = 7'h44 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_68; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_966 = 7'h45 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_69; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_967 = 7'h46 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_70; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_968 = 7'h47 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_71; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_969 = 7'h48 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_72; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_970 = 7'h49 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_73; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_971 = 7'h4a == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_74; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_972 = 7'h4b == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_75; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_973 = 7'h4c == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_76; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_974 = 7'h4d == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_77; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_975 = 7'h4e == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_78; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_976 = 7'h4f == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_79; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_977 = 7'h50 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_80; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_978 = 7'h51 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_81; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_979 = 7'h52 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_82; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_980 = 7'h53 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_83; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_981 = 7'h54 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_84; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_982 = 7'h55 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_85; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_983 = 7'h56 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_86; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_984 = 7'h57 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_87; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_985 = 7'h58 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_88; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_986 = 7'h59 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_89; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_987 = 7'h5a == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_90; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_988 = 7'h5b == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_91; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_989 = 7'h5c == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_92; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_990 = 7'h5d == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_93; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_991 = 7'h5e == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_94; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_992 = 7'h5f == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_95; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_993 = 7'h60 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_96; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_994 = 7'h61 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_97; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_995 = 7'h62 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_98; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_996 = 7'h63 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_99; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_997 = 7'h64 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_100; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_998 = 7'h65 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_101; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_999 = 7'h66 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_102; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1000 = 7'h67 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_103; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1001 = 7'h68 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_104; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1002 = 7'h69 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_105; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1003 = 7'h6a == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_106; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1004 = 7'h6b == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_107; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1005 = 7'h6c == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_108; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1006 = 7'h6d == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_109; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1007 = 7'h6e == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_110; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1008 = 7'h6f == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_111; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1009 = 7'h70 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_112; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1010 = 7'h71 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_113; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1011 = 7'h72 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_114; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1012 = 7'h73 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_115; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1013 = 7'h74 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_116; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1014 = 7'h75 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_117; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1015 = 7'h76 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_118; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1016 = 7'h77 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_119; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1017 = 7'h78 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_120; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1018 = 7'h79 == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_121; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1019 = 7'h7a == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_122; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1020 = 7'h7b == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_123; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1021 = 7'h7c == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_124; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1022 = 7'h7d == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_125; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1023 = 7'h7e == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_126; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [63:0] _GEN_1024 = 7'h7f == rob_alloc_ids_0 ? _rob_tscs_T_25 : rob_tscs_127; // @[TestHarness.scala 155:21 184:{36,36}]
  wire [31:0] _GEN_1025 = igen_io_fire ? _GEN_1 : rob_payload_0_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1026 = igen_io_fire ? _GEN_2 : rob_payload_1_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1027 = igen_io_fire ? _GEN_3 : rob_payload_2_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1028 = igen_io_fire ? _GEN_4 : rob_payload_3_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1029 = igen_io_fire ? _GEN_5 : rob_payload_4_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1030 = igen_io_fire ? _GEN_6 : rob_payload_5_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1031 = igen_io_fire ? _GEN_7 : rob_payload_6_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1032 = igen_io_fire ? _GEN_8 : rob_payload_7_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1033 = igen_io_fire ? _GEN_9 : rob_payload_8_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1034 = igen_io_fire ? _GEN_10 : rob_payload_9_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1035 = igen_io_fire ? _GEN_11 : rob_payload_10_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1036 = igen_io_fire ? _GEN_12 : rob_payload_11_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1037 = igen_io_fire ? _GEN_13 : rob_payload_12_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1038 = igen_io_fire ? _GEN_14 : rob_payload_13_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1039 = igen_io_fire ? _GEN_15 : rob_payload_14_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1040 = igen_io_fire ? _GEN_16 : rob_payload_15_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1041 = igen_io_fire ? _GEN_17 : rob_payload_16_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1042 = igen_io_fire ? _GEN_18 : rob_payload_17_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1043 = igen_io_fire ? _GEN_19 : rob_payload_18_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1044 = igen_io_fire ? _GEN_20 : rob_payload_19_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1045 = igen_io_fire ? _GEN_21 : rob_payload_20_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1046 = igen_io_fire ? _GEN_22 : rob_payload_21_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1047 = igen_io_fire ? _GEN_23 : rob_payload_22_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1048 = igen_io_fire ? _GEN_24 : rob_payload_23_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1049 = igen_io_fire ? _GEN_25 : rob_payload_24_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1050 = igen_io_fire ? _GEN_26 : rob_payload_25_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1051 = igen_io_fire ? _GEN_27 : rob_payload_26_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1052 = igen_io_fire ? _GEN_28 : rob_payload_27_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1053 = igen_io_fire ? _GEN_29 : rob_payload_28_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1054 = igen_io_fire ? _GEN_30 : rob_payload_29_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1055 = igen_io_fire ? _GEN_31 : rob_payload_30_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1056 = igen_io_fire ? _GEN_32 : rob_payload_31_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1057 = igen_io_fire ? _GEN_33 : rob_payload_32_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1058 = igen_io_fire ? _GEN_34 : rob_payload_33_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1059 = igen_io_fire ? _GEN_35 : rob_payload_34_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1060 = igen_io_fire ? _GEN_36 : rob_payload_35_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1061 = igen_io_fire ? _GEN_37 : rob_payload_36_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1062 = igen_io_fire ? _GEN_38 : rob_payload_37_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1063 = igen_io_fire ? _GEN_39 : rob_payload_38_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1064 = igen_io_fire ? _GEN_40 : rob_payload_39_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1065 = igen_io_fire ? _GEN_41 : rob_payload_40_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1066 = igen_io_fire ? _GEN_42 : rob_payload_41_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1067 = igen_io_fire ? _GEN_43 : rob_payload_42_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1068 = igen_io_fire ? _GEN_44 : rob_payload_43_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1069 = igen_io_fire ? _GEN_45 : rob_payload_44_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1070 = igen_io_fire ? _GEN_46 : rob_payload_45_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1071 = igen_io_fire ? _GEN_47 : rob_payload_46_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1072 = igen_io_fire ? _GEN_48 : rob_payload_47_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1073 = igen_io_fire ? _GEN_49 : rob_payload_48_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1074 = igen_io_fire ? _GEN_50 : rob_payload_49_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1075 = igen_io_fire ? _GEN_51 : rob_payload_50_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1076 = igen_io_fire ? _GEN_52 : rob_payload_51_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1077 = igen_io_fire ? _GEN_53 : rob_payload_52_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1078 = igen_io_fire ? _GEN_54 : rob_payload_53_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1079 = igen_io_fire ? _GEN_55 : rob_payload_54_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1080 = igen_io_fire ? _GEN_56 : rob_payload_55_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1081 = igen_io_fire ? _GEN_57 : rob_payload_56_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1082 = igen_io_fire ? _GEN_58 : rob_payload_57_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1083 = igen_io_fire ? _GEN_59 : rob_payload_58_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1084 = igen_io_fire ? _GEN_60 : rob_payload_59_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1085 = igen_io_fire ? _GEN_61 : rob_payload_60_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1086 = igen_io_fire ? _GEN_62 : rob_payload_61_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1087 = igen_io_fire ? _GEN_63 : rob_payload_62_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1088 = igen_io_fire ? _GEN_64 : rob_payload_63_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1089 = igen_io_fire ? _GEN_65 : rob_payload_64_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1090 = igen_io_fire ? _GEN_66 : rob_payload_65_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1091 = igen_io_fire ? _GEN_67 : rob_payload_66_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1092 = igen_io_fire ? _GEN_68 : rob_payload_67_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1093 = igen_io_fire ? _GEN_69 : rob_payload_68_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1094 = igen_io_fire ? _GEN_70 : rob_payload_69_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1095 = igen_io_fire ? _GEN_71 : rob_payload_70_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1096 = igen_io_fire ? _GEN_72 : rob_payload_71_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1097 = igen_io_fire ? _GEN_73 : rob_payload_72_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1098 = igen_io_fire ? _GEN_74 : rob_payload_73_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1099 = igen_io_fire ? _GEN_75 : rob_payload_74_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1100 = igen_io_fire ? _GEN_76 : rob_payload_75_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1101 = igen_io_fire ? _GEN_77 : rob_payload_76_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1102 = igen_io_fire ? _GEN_78 : rob_payload_77_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1103 = igen_io_fire ? _GEN_79 : rob_payload_78_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1104 = igen_io_fire ? _GEN_80 : rob_payload_79_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1105 = igen_io_fire ? _GEN_81 : rob_payload_80_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1106 = igen_io_fire ? _GEN_82 : rob_payload_81_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1107 = igen_io_fire ? _GEN_83 : rob_payload_82_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1108 = igen_io_fire ? _GEN_84 : rob_payload_83_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1109 = igen_io_fire ? _GEN_85 : rob_payload_84_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1110 = igen_io_fire ? _GEN_86 : rob_payload_85_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1111 = igen_io_fire ? _GEN_87 : rob_payload_86_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1112 = igen_io_fire ? _GEN_88 : rob_payload_87_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1113 = igen_io_fire ? _GEN_89 : rob_payload_88_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1114 = igen_io_fire ? _GEN_90 : rob_payload_89_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1115 = igen_io_fire ? _GEN_91 : rob_payload_90_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1116 = igen_io_fire ? _GEN_92 : rob_payload_91_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1117 = igen_io_fire ? _GEN_93 : rob_payload_92_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1118 = igen_io_fire ? _GEN_94 : rob_payload_93_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1119 = igen_io_fire ? _GEN_95 : rob_payload_94_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1120 = igen_io_fire ? _GEN_96 : rob_payload_95_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1121 = igen_io_fire ? _GEN_97 : rob_payload_96_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1122 = igen_io_fire ? _GEN_98 : rob_payload_97_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1123 = igen_io_fire ? _GEN_99 : rob_payload_98_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1124 = igen_io_fire ? _GEN_100 : rob_payload_99_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1125 = igen_io_fire ? _GEN_101 : rob_payload_100_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1126 = igen_io_fire ? _GEN_102 : rob_payload_101_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1127 = igen_io_fire ? _GEN_103 : rob_payload_102_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1128 = igen_io_fire ? _GEN_104 : rob_payload_103_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1129 = igen_io_fire ? _GEN_105 : rob_payload_104_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1130 = igen_io_fire ? _GEN_106 : rob_payload_105_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1131 = igen_io_fire ? _GEN_107 : rob_payload_106_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1132 = igen_io_fire ? _GEN_108 : rob_payload_107_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1133 = igen_io_fire ? _GEN_109 : rob_payload_108_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1134 = igen_io_fire ? _GEN_110 : rob_payload_109_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1135 = igen_io_fire ? _GEN_111 : rob_payload_110_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1136 = igen_io_fire ? _GEN_112 : rob_payload_111_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1137 = igen_io_fire ? _GEN_113 : rob_payload_112_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1138 = igen_io_fire ? _GEN_114 : rob_payload_113_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1139 = igen_io_fire ? _GEN_115 : rob_payload_114_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1140 = igen_io_fire ? _GEN_116 : rob_payload_115_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1141 = igen_io_fire ? _GEN_117 : rob_payload_116_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1142 = igen_io_fire ? _GEN_118 : rob_payload_117_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1143 = igen_io_fire ? _GEN_119 : rob_payload_118_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1144 = igen_io_fire ? _GEN_120 : rob_payload_119_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1145 = igen_io_fire ? _GEN_121 : rob_payload_120_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1146 = igen_io_fire ? _GEN_122 : rob_payload_121_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1147 = igen_io_fire ? _GEN_123 : rob_payload_122_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1148 = igen_io_fire ? _GEN_124 : rob_payload_123_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1149 = igen_io_fire ? _GEN_125 : rob_payload_124_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1150 = igen_io_fire ? _GEN_126 : rob_payload_125_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1151 = igen_io_fire ? _GEN_127 : rob_payload_126_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [31:0] _GEN_1152 = igen_io_fire ? _GEN_128 : rob_payload_127_tsc; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1153 = igen_io_fire ? _GEN_129 : rob_payload_0_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1154 = igen_io_fire ? _GEN_130 : rob_payload_1_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1155 = igen_io_fire ? _GEN_131 : rob_payload_2_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1156 = igen_io_fire ? _GEN_132 : rob_payload_3_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1157 = igen_io_fire ? _GEN_133 : rob_payload_4_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1158 = igen_io_fire ? _GEN_134 : rob_payload_5_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1159 = igen_io_fire ? _GEN_135 : rob_payload_6_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1160 = igen_io_fire ? _GEN_136 : rob_payload_7_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1161 = igen_io_fire ? _GEN_137 : rob_payload_8_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1162 = igen_io_fire ? _GEN_138 : rob_payload_9_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1163 = igen_io_fire ? _GEN_139 : rob_payload_10_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1164 = igen_io_fire ? _GEN_140 : rob_payload_11_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1165 = igen_io_fire ? _GEN_141 : rob_payload_12_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1166 = igen_io_fire ? _GEN_142 : rob_payload_13_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1167 = igen_io_fire ? _GEN_143 : rob_payload_14_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1168 = igen_io_fire ? _GEN_144 : rob_payload_15_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1169 = igen_io_fire ? _GEN_145 : rob_payload_16_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1170 = igen_io_fire ? _GEN_146 : rob_payload_17_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1171 = igen_io_fire ? _GEN_147 : rob_payload_18_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1172 = igen_io_fire ? _GEN_148 : rob_payload_19_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1173 = igen_io_fire ? _GEN_149 : rob_payload_20_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1174 = igen_io_fire ? _GEN_150 : rob_payload_21_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1175 = igen_io_fire ? _GEN_151 : rob_payload_22_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1176 = igen_io_fire ? _GEN_152 : rob_payload_23_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1177 = igen_io_fire ? _GEN_153 : rob_payload_24_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1178 = igen_io_fire ? _GEN_154 : rob_payload_25_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1179 = igen_io_fire ? _GEN_155 : rob_payload_26_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1180 = igen_io_fire ? _GEN_156 : rob_payload_27_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1181 = igen_io_fire ? _GEN_157 : rob_payload_28_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1182 = igen_io_fire ? _GEN_158 : rob_payload_29_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1183 = igen_io_fire ? _GEN_159 : rob_payload_30_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1184 = igen_io_fire ? _GEN_160 : rob_payload_31_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1185 = igen_io_fire ? _GEN_161 : rob_payload_32_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1186 = igen_io_fire ? _GEN_162 : rob_payload_33_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1187 = igen_io_fire ? _GEN_163 : rob_payload_34_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1188 = igen_io_fire ? _GEN_164 : rob_payload_35_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1189 = igen_io_fire ? _GEN_165 : rob_payload_36_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1190 = igen_io_fire ? _GEN_166 : rob_payload_37_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1191 = igen_io_fire ? _GEN_167 : rob_payload_38_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1192 = igen_io_fire ? _GEN_168 : rob_payload_39_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1193 = igen_io_fire ? _GEN_169 : rob_payload_40_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1194 = igen_io_fire ? _GEN_170 : rob_payload_41_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1195 = igen_io_fire ? _GEN_171 : rob_payload_42_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1196 = igen_io_fire ? _GEN_172 : rob_payload_43_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1197 = igen_io_fire ? _GEN_173 : rob_payload_44_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1198 = igen_io_fire ? _GEN_174 : rob_payload_45_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1199 = igen_io_fire ? _GEN_175 : rob_payload_46_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1200 = igen_io_fire ? _GEN_176 : rob_payload_47_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1201 = igen_io_fire ? _GEN_177 : rob_payload_48_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1202 = igen_io_fire ? _GEN_178 : rob_payload_49_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1203 = igen_io_fire ? _GEN_179 : rob_payload_50_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1204 = igen_io_fire ? _GEN_180 : rob_payload_51_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1205 = igen_io_fire ? _GEN_181 : rob_payload_52_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1206 = igen_io_fire ? _GEN_182 : rob_payload_53_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1207 = igen_io_fire ? _GEN_183 : rob_payload_54_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1208 = igen_io_fire ? _GEN_184 : rob_payload_55_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1209 = igen_io_fire ? _GEN_185 : rob_payload_56_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1210 = igen_io_fire ? _GEN_186 : rob_payload_57_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1211 = igen_io_fire ? _GEN_187 : rob_payload_58_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1212 = igen_io_fire ? _GEN_188 : rob_payload_59_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1213 = igen_io_fire ? _GEN_189 : rob_payload_60_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1214 = igen_io_fire ? _GEN_190 : rob_payload_61_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1215 = igen_io_fire ? _GEN_191 : rob_payload_62_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1216 = igen_io_fire ? _GEN_192 : rob_payload_63_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1217 = igen_io_fire ? _GEN_193 : rob_payload_64_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1218 = igen_io_fire ? _GEN_194 : rob_payload_65_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1219 = igen_io_fire ? _GEN_195 : rob_payload_66_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1220 = igen_io_fire ? _GEN_196 : rob_payload_67_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1221 = igen_io_fire ? _GEN_197 : rob_payload_68_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1222 = igen_io_fire ? _GEN_198 : rob_payload_69_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1223 = igen_io_fire ? _GEN_199 : rob_payload_70_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1224 = igen_io_fire ? _GEN_200 : rob_payload_71_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1225 = igen_io_fire ? _GEN_201 : rob_payload_72_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1226 = igen_io_fire ? _GEN_202 : rob_payload_73_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1227 = igen_io_fire ? _GEN_203 : rob_payload_74_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1228 = igen_io_fire ? _GEN_204 : rob_payload_75_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1229 = igen_io_fire ? _GEN_205 : rob_payload_76_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1230 = igen_io_fire ? _GEN_206 : rob_payload_77_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1231 = igen_io_fire ? _GEN_207 : rob_payload_78_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1232 = igen_io_fire ? _GEN_208 : rob_payload_79_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1233 = igen_io_fire ? _GEN_209 : rob_payload_80_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1234 = igen_io_fire ? _GEN_210 : rob_payload_81_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1235 = igen_io_fire ? _GEN_211 : rob_payload_82_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1236 = igen_io_fire ? _GEN_212 : rob_payload_83_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1237 = igen_io_fire ? _GEN_213 : rob_payload_84_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1238 = igen_io_fire ? _GEN_214 : rob_payload_85_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1239 = igen_io_fire ? _GEN_215 : rob_payload_86_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1240 = igen_io_fire ? _GEN_216 : rob_payload_87_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1241 = igen_io_fire ? _GEN_217 : rob_payload_88_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1242 = igen_io_fire ? _GEN_218 : rob_payload_89_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1243 = igen_io_fire ? _GEN_219 : rob_payload_90_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1244 = igen_io_fire ? _GEN_220 : rob_payload_91_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1245 = igen_io_fire ? _GEN_221 : rob_payload_92_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1246 = igen_io_fire ? _GEN_222 : rob_payload_93_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1247 = igen_io_fire ? _GEN_223 : rob_payload_94_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1248 = igen_io_fire ? _GEN_224 : rob_payload_95_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1249 = igen_io_fire ? _GEN_225 : rob_payload_96_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1250 = igen_io_fire ? _GEN_226 : rob_payload_97_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1251 = igen_io_fire ? _GEN_227 : rob_payload_98_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1252 = igen_io_fire ? _GEN_228 : rob_payload_99_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1253 = igen_io_fire ? _GEN_229 : rob_payload_100_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1254 = igen_io_fire ? _GEN_230 : rob_payload_101_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1255 = igen_io_fire ? _GEN_231 : rob_payload_102_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1256 = igen_io_fire ? _GEN_232 : rob_payload_103_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1257 = igen_io_fire ? _GEN_233 : rob_payload_104_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1258 = igen_io_fire ? _GEN_234 : rob_payload_105_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1259 = igen_io_fire ? _GEN_235 : rob_payload_106_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1260 = igen_io_fire ? _GEN_236 : rob_payload_107_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1261 = igen_io_fire ? _GEN_237 : rob_payload_108_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1262 = igen_io_fire ? _GEN_238 : rob_payload_109_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1263 = igen_io_fire ? _GEN_239 : rob_payload_110_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1264 = igen_io_fire ? _GEN_240 : rob_payload_111_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1265 = igen_io_fire ? _GEN_241 : rob_payload_112_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1266 = igen_io_fire ? _GEN_242 : rob_payload_113_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1267 = igen_io_fire ? _GEN_243 : rob_payload_114_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1268 = igen_io_fire ? _GEN_244 : rob_payload_115_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1269 = igen_io_fire ? _GEN_245 : rob_payload_116_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1270 = igen_io_fire ? _GEN_246 : rob_payload_117_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1271 = igen_io_fire ? _GEN_247 : rob_payload_118_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1272 = igen_io_fire ? _GEN_248 : rob_payload_119_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1273 = igen_io_fire ? _GEN_249 : rob_payload_120_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1274 = igen_io_fire ? _GEN_250 : rob_payload_121_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1275 = igen_io_fire ? _GEN_251 : rob_payload_122_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1276 = igen_io_fire ? _GEN_252 : rob_payload_123_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1277 = igen_io_fire ? _GEN_253 : rob_payload_124_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1278 = igen_io_fire ? _GEN_254 : rob_payload_125_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1279 = igen_io_fire ? _GEN_255 : rob_payload_126_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1280 = igen_io_fire ? _GEN_256 : rob_payload_127_rob_idx; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1281 = igen_io_fire ? _GEN_257 : rob_payload_0_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1282 = igen_io_fire ? _GEN_258 : rob_payload_1_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1283 = igen_io_fire ? _GEN_259 : rob_payload_2_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1284 = igen_io_fire ? _GEN_260 : rob_payload_3_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1285 = igen_io_fire ? _GEN_261 : rob_payload_4_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1286 = igen_io_fire ? _GEN_262 : rob_payload_5_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1287 = igen_io_fire ? _GEN_263 : rob_payload_6_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1288 = igen_io_fire ? _GEN_264 : rob_payload_7_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1289 = igen_io_fire ? _GEN_265 : rob_payload_8_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1290 = igen_io_fire ? _GEN_266 : rob_payload_9_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1291 = igen_io_fire ? _GEN_267 : rob_payload_10_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1292 = igen_io_fire ? _GEN_268 : rob_payload_11_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1293 = igen_io_fire ? _GEN_269 : rob_payload_12_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1294 = igen_io_fire ? _GEN_270 : rob_payload_13_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1295 = igen_io_fire ? _GEN_271 : rob_payload_14_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1296 = igen_io_fire ? _GEN_272 : rob_payload_15_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1297 = igen_io_fire ? _GEN_273 : rob_payload_16_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1298 = igen_io_fire ? _GEN_274 : rob_payload_17_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1299 = igen_io_fire ? _GEN_275 : rob_payload_18_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1300 = igen_io_fire ? _GEN_276 : rob_payload_19_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1301 = igen_io_fire ? _GEN_277 : rob_payload_20_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1302 = igen_io_fire ? _GEN_278 : rob_payload_21_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1303 = igen_io_fire ? _GEN_279 : rob_payload_22_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1304 = igen_io_fire ? _GEN_280 : rob_payload_23_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1305 = igen_io_fire ? _GEN_281 : rob_payload_24_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1306 = igen_io_fire ? _GEN_282 : rob_payload_25_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1307 = igen_io_fire ? _GEN_283 : rob_payload_26_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1308 = igen_io_fire ? _GEN_284 : rob_payload_27_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1309 = igen_io_fire ? _GEN_285 : rob_payload_28_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1310 = igen_io_fire ? _GEN_286 : rob_payload_29_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1311 = igen_io_fire ? _GEN_287 : rob_payload_30_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1312 = igen_io_fire ? _GEN_288 : rob_payload_31_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1313 = igen_io_fire ? _GEN_289 : rob_payload_32_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1314 = igen_io_fire ? _GEN_290 : rob_payload_33_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1315 = igen_io_fire ? _GEN_291 : rob_payload_34_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1316 = igen_io_fire ? _GEN_292 : rob_payload_35_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1317 = igen_io_fire ? _GEN_293 : rob_payload_36_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1318 = igen_io_fire ? _GEN_294 : rob_payload_37_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1319 = igen_io_fire ? _GEN_295 : rob_payload_38_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1320 = igen_io_fire ? _GEN_296 : rob_payload_39_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1321 = igen_io_fire ? _GEN_297 : rob_payload_40_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1322 = igen_io_fire ? _GEN_298 : rob_payload_41_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1323 = igen_io_fire ? _GEN_299 : rob_payload_42_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1324 = igen_io_fire ? _GEN_300 : rob_payload_43_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1325 = igen_io_fire ? _GEN_301 : rob_payload_44_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1326 = igen_io_fire ? _GEN_302 : rob_payload_45_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1327 = igen_io_fire ? _GEN_303 : rob_payload_46_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1328 = igen_io_fire ? _GEN_304 : rob_payload_47_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1329 = igen_io_fire ? _GEN_305 : rob_payload_48_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1330 = igen_io_fire ? _GEN_306 : rob_payload_49_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1331 = igen_io_fire ? _GEN_307 : rob_payload_50_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1332 = igen_io_fire ? _GEN_308 : rob_payload_51_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1333 = igen_io_fire ? _GEN_309 : rob_payload_52_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1334 = igen_io_fire ? _GEN_310 : rob_payload_53_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1335 = igen_io_fire ? _GEN_311 : rob_payload_54_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1336 = igen_io_fire ? _GEN_312 : rob_payload_55_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1337 = igen_io_fire ? _GEN_313 : rob_payload_56_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1338 = igen_io_fire ? _GEN_314 : rob_payload_57_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1339 = igen_io_fire ? _GEN_315 : rob_payload_58_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1340 = igen_io_fire ? _GEN_316 : rob_payload_59_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1341 = igen_io_fire ? _GEN_317 : rob_payload_60_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1342 = igen_io_fire ? _GEN_318 : rob_payload_61_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1343 = igen_io_fire ? _GEN_319 : rob_payload_62_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1344 = igen_io_fire ? _GEN_320 : rob_payload_63_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1345 = igen_io_fire ? _GEN_321 : rob_payload_64_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1346 = igen_io_fire ? _GEN_322 : rob_payload_65_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1347 = igen_io_fire ? _GEN_323 : rob_payload_66_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1348 = igen_io_fire ? _GEN_324 : rob_payload_67_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1349 = igen_io_fire ? _GEN_325 : rob_payload_68_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1350 = igen_io_fire ? _GEN_326 : rob_payload_69_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1351 = igen_io_fire ? _GEN_327 : rob_payload_70_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1352 = igen_io_fire ? _GEN_328 : rob_payload_71_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1353 = igen_io_fire ? _GEN_329 : rob_payload_72_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1354 = igen_io_fire ? _GEN_330 : rob_payload_73_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1355 = igen_io_fire ? _GEN_331 : rob_payload_74_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1356 = igen_io_fire ? _GEN_332 : rob_payload_75_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1357 = igen_io_fire ? _GEN_333 : rob_payload_76_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1358 = igen_io_fire ? _GEN_334 : rob_payload_77_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1359 = igen_io_fire ? _GEN_335 : rob_payload_78_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1360 = igen_io_fire ? _GEN_336 : rob_payload_79_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1361 = igen_io_fire ? _GEN_337 : rob_payload_80_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1362 = igen_io_fire ? _GEN_338 : rob_payload_81_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1363 = igen_io_fire ? _GEN_339 : rob_payload_82_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1364 = igen_io_fire ? _GEN_340 : rob_payload_83_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1365 = igen_io_fire ? _GEN_341 : rob_payload_84_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1366 = igen_io_fire ? _GEN_342 : rob_payload_85_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1367 = igen_io_fire ? _GEN_343 : rob_payload_86_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1368 = igen_io_fire ? _GEN_344 : rob_payload_87_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1369 = igen_io_fire ? _GEN_345 : rob_payload_88_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1370 = igen_io_fire ? _GEN_346 : rob_payload_89_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1371 = igen_io_fire ? _GEN_347 : rob_payload_90_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1372 = igen_io_fire ? _GEN_348 : rob_payload_91_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1373 = igen_io_fire ? _GEN_349 : rob_payload_92_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1374 = igen_io_fire ? _GEN_350 : rob_payload_93_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1375 = igen_io_fire ? _GEN_351 : rob_payload_94_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1376 = igen_io_fire ? _GEN_352 : rob_payload_95_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1377 = igen_io_fire ? _GEN_353 : rob_payload_96_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1378 = igen_io_fire ? _GEN_354 : rob_payload_97_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1379 = igen_io_fire ? _GEN_355 : rob_payload_98_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1380 = igen_io_fire ? _GEN_356 : rob_payload_99_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1381 = igen_io_fire ? _GEN_357 : rob_payload_100_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1382 = igen_io_fire ? _GEN_358 : rob_payload_101_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1383 = igen_io_fire ? _GEN_359 : rob_payload_102_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1384 = igen_io_fire ? _GEN_360 : rob_payload_103_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1385 = igen_io_fire ? _GEN_361 : rob_payload_104_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1386 = igen_io_fire ? _GEN_362 : rob_payload_105_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1387 = igen_io_fire ? _GEN_363 : rob_payload_106_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1388 = igen_io_fire ? _GEN_364 : rob_payload_107_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1389 = igen_io_fire ? _GEN_365 : rob_payload_108_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1390 = igen_io_fire ? _GEN_366 : rob_payload_109_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1391 = igen_io_fire ? _GEN_367 : rob_payload_110_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1392 = igen_io_fire ? _GEN_368 : rob_payload_111_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1393 = igen_io_fire ? _GEN_369 : rob_payload_112_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1394 = igen_io_fire ? _GEN_370 : rob_payload_113_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1395 = igen_io_fire ? _GEN_371 : rob_payload_114_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1396 = igen_io_fire ? _GEN_372 : rob_payload_115_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1397 = igen_io_fire ? _GEN_373 : rob_payload_116_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1398 = igen_io_fire ? _GEN_374 : rob_payload_117_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1399 = igen_io_fire ? _GEN_375 : rob_payload_118_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1400 = igen_io_fire ? _GEN_376 : rob_payload_119_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1401 = igen_io_fire ? _GEN_377 : rob_payload_120_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1402 = igen_io_fire ? _GEN_378 : rob_payload_121_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1403 = igen_io_fire ? _GEN_379 : rob_payload_122_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1404 = igen_io_fire ? _GEN_380 : rob_payload_123_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1405 = igen_io_fire ? _GEN_381 : rob_payload_124_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1406 = igen_io_fire ? _GEN_382 : rob_payload_125_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1407 = igen_io_fire ? _GEN_383 : rob_payload_126_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire [15:0] _GEN_1408 = igen_io_fire ? _GEN_384 : rob_payload_127_flits_fired; // @[TestHarness.scala 150:24 178:25]
  wire  _GEN_1409 = igen_io_fire ? _GEN_385 : rob_egress_id_0; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1410 = igen_io_fire ? _GEN_386 : rob_egress_id_1; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1411 = igen_io_fire ? _GEN_387 : rob_egress_id_2; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1412 = igen_io_fire ? _GEN_388 : rob_egress_id_3; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1413 = igen_io_fire ? _GEN_389 : rob_egress_id_4; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1414 = igen_io_fire ? _GEN_390 : rob_egress_id_5; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1415 = igen_io_fire ? _GEN_391 : rob_egress_id_6; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1416 = igen_io_fire ? _GEN_392 : rob_egress_id_7; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1417 = igen_io_fire ? _GEN_393 : rob_egress_id_8; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1418 = igen_io_fire ? _GEN_394 : rob_egress_id_9; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1419 = igen_io_fire ? _GEN_395 : rob_egress_id_10; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1420 = igen_io_fire ? _GEN_396 : rob_egress_id_11; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1421 = igen_io_fire ? _GEN_397 : rob_egress_id_12; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1422 = igen_io_fire ? _GEN_398 : rob_egress_id_13; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1423 = igen_io_fire ? _GEN_399 : rob_egress_id_14; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1424 = igen_io_fire ? _GEN_400 : rob_egress_id_15; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1425 = igen_io_fire ? _GEN_401 : rob_egress_id_16; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1426 = igen_io_fire ? _GEN_402 : rob_egress_id_17; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1427 = igen_io_fire ? _GEN_403 : rob_egress_id_18; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1428 = igen_io_fire ? _GEN_404 : rob_egress_id_19; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1429 = igen_io_fire ? _GEN_405 : rob_egress_id_20; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1430 = igen_io_fire ? _GEN_406 : rob_egress_id_21; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1431 = igen_io_fire ? _GEN_407 : rob_egress_id_22; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1432 = igen_io_fire ? _GEN_408 : rob_egress_id_23; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1433 = igen_io_fire ? _GEN_409 : rob_egress_id_24; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1434 = igen_io_fire ? _GEN_410 : rob_egress_id_25; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1435 = igen_io_fire ? _GEN_411 : rob_egress_id_26; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1436 = igen_io_fire ? _GEN_412 : rob_egress_id_27; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1437 = igen_io_fire ? _GEN_413 : rob_egress_id_28; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1438 = igen_io_fire ? _GEN_414 : rob_egress_id_29; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1439 = igen_io_fire ? _GEN_415 : rob_egress_id_30; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1440 = igen_io_fire ? _GEN_416 : rob_egress_id_31; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1441 = igen_io_fire ? _GEN_417 : rob_egress_id_32; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1442 = igen_io_fire ? _GEN_418 : rob_egress_id_33; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1443 = igen_io_fire ? _GEN_419 : rob_egress_id_34; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1444 = igen_io_fire ? _GEN_420 : rob_egress_id_35; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1445 = igen_io_fire ? _GEN_421 : rob_egress_id_36; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1446 = igen_io_fire ? _GEN_422 : rob_egress_id_37; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1447 = igen_io_fire ? _GEN_423 : rob_egress_id_38; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1448 = igen_io_fire ? _GEN_424 : rob_egress_id_39; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1449 = igen_io_fire ? _GEN_425 : rob_egress_id_40; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1450 = igen_io_fire ? _GEN_426 : rob_egress_id_41; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1451 = igen_io_fire ? _GEN_427 : rob_egress_id_42; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1452 = igen_io_fire ? _GEN_428 : rob_egress_id_43; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1453 = igen_io_fire ? _GEN_429 : rob_egress_id_44; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1454 = igen_io_fire ? _GEN_430 : rob_egress_id_45; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1455 = igen_io_fire ? _GEN_431 : rob_egress_id_46; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1456 = igen_io_fire ? _GEN_432 : rob_egress_id_47; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1457 = igen_io_fire ? _GEN_433 : rob_egress_id_48; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1458 = igen_io_fire ? _GEN_434 : rob_egress_id_49; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1459 = igen_io_fire ? _GEN_435 : rob_egress_id_50; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1460 = igen_io_fire ? _GEN_436 : rob_egress_id_51; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1461 = igen_io_fire ? _GEN_437 : rob_egress_id_52; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1462 = igen_io_fire ? _GEN_438 : rob_egress_id_53; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1463 = igen_io_fire ? _GEN_439 : rob_egress_id_54; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1464 = igen_io_fire ? _GEN_440 : rob_egress_id_55; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1465 = igen_io_fire ? _GEN_441 : rob_egress_id_56; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1466 = igen_io_fire ? _GEN_442 : rob_egress_id_57; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1467 = igen_io_fire ? _GEN_443 : rob_egress_id_58; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1468 = igen_io_fire ? _GEN_444 : rob_egress_id_59; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1469 = igen_io_fire ? _GEN_445 : rob_egress_id_60; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1470 = igen_io_fire ? _GEN_446 : rob_egress_id_61; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1471 = igen_io_fire ? _GEN_447 : rob_egress_id_62; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1472 = igen_io_fire ? _GEN_448 : rob_egress_id_63; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1473 = igen_io_fire ? _GEN_449 : rob_egress_id_64; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1474 = igen_io_fire ? _GEN_450 : rob_egress_id_65; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1475 = igen_io_fire ? _GEN_451 : rob_egress_id_66; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1476 = igen_io_fire ? _GEN_452 : rob_egress_id_67; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1477 = igen_io_fire ? _GEN_453 : rob_egress_id_68; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1478 = igen_io_fire ? _GEN_454 : rob_egress_id_69; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1479 = igen_io_fire ? _GEN_455 : rob_egress_id_70; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1480 = igen_io_fire ? _GEN_456 : rob_egress_id_71; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1481 = igen_io_fire ? _GEN_457 : rob_egress_id_72; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1482 = igen_io_fire ? _GEN_458 : rob_egress_id_73; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1483 = igen_io_fire ? _GEN_459 : rob_egress_id_74; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1484 = igen_io_fire ? _GEN_460 : rob_egress_id_75; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1485 = igen_io_fire ? _GEN_461 : rob_egress_id_76; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1486 = igen_io_fire ? _GEN_462 : rob_egress_id_77; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1487 = igen_io_fire ? _GEN_463 : rob_egress_id_78; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1488 = igen_io_fire ? _GEN_464 : rob_egress_id_79; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1489 = igen_io_fire ? _GEN_465 : rob_egress_id_80; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1490 = igen_io_fire ? _GEN_466 : rob_egress_id_81; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1491 = igen_io_fire ? _GEN_467 : rob_egress_id_82; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1492 = igen_io_fire ? _GEN_468 : rob_egress_id_83; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1493 = igen_io_fire ? _GEN_469 : rob_egress_id_84; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1494 = igen_io_fire ? _GEN_470 : rob_egress_id_85; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1495 = igen_io_fire ? _GEN_471 : rob_egress_id_86; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1496 = igen_io_fire ? _GEN_472 : rob_egress_id_87; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1497 = igen_io_fire ? _GEN_473 : rob_egress_id_88; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1498 = igen_io_fire ? _GEN_474 : rob_egress_id_89; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1499 = igen_io_fire ? _GEN_475 : rob_egress_id_90; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1500 = igen_io_fire ? _GEN_476 : rob_egress_id_91; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1501 = igen_io_fire ? _GEN_477 : rob_egress_id_92; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1502 = igen_io_fire ? _GEN_478 : rob_egress_id_93; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1503 = igen_io_fire ? _GEN_479 : rob_egress_id_94; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1504 = igen_io_fire ? _GEN_480 : rob_egress_id_95; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1505 = igen_io_fire ? _GEN_481 : rob_egress_id_96; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1506 = igen_io_fire ? _GEN_482 : rob_egress_id_97; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1507 = igen_io_fire ? _GEN_483 : rob_egress_id_98; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1508 = igen_io_fire ? _GEN_484 : rob_egress_id_99; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1509 = igen_io_fire ? _GEN_485 : rob_egress_id_100; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1510 = igen_io_fire ? _GEN_486 : rob_egress_id_101; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1511 = igen_io_fire ? _GEN_487 : rob_egress_id_102; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1512 = igen_io_fire ? _GEN_488 : rob_egress_id_103; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1513 = igen_io_fire ? _GEN_489 : rob_egress_id_104; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1514 = igen_io_fire ? _GEN_490 : rob_egress_id_105; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1515 = igen_io_fire ? _GEN_491 : rob_egress_id_106; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1516 = igen_io_fire ? _GEN_492 : rob_egress_id_107; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1517 = igen_io_fire ? _GEN_493 : rob_egress_id_108; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1518 = igen_io_fire ? _GEN_494 : rob_egress_id_109; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1519 = igen_io_fire ? _GEN_495 : rob_egress_id_110; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1520 = igen_io_fire ? _GEN_496 : rob_egress_id_111; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1521 = igen_io_fire ? _GEN_497 : rob_egress_id_112; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1522 = igen_io_fire ? _GEN_498 : rob_egress_id_113; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1523 = igen_io_fire ? _GEN_499 : rob_egress_id_114; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1524 = igen_io_fire ? _GEN_500 : rob_egress_id_115; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1525 = igen_io_fire ? _GEN_501 : rob_egress_id_116; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1526 = igen_io_fire ? _GEN_502 : rob_egress_id_117; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1527 = igen_io_fire ? _GEN_503 : rob_egress_id_118; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1528 = igen_io_fire ? _GEN_504 : rob_egress_id_119; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1529 = igen_io_fire ? _GEN_505 : rob_egress_id_120; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1530 = igen_io_fire ? _GEN_506 : rob_egress_id_121; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1531 = igen_io_fire ? _GEN_507 : rob_egress_id_122; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1532 = igen_io_fire ? _GEN_508 : rob_egress_id_123; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1533 = igen_io_fire ? _GEN_509 : rob_egress_id_124; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1534 = igen_io_fire ? _GEN_510 : rob_egress_id_125; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1535 = igen_io_fire ? _GEN_511 : rob_egress_id_126; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1536 = igen_io_fire ? _GEN_512 : rob_egress_id_127; // @[TestHarness.scala 178:25 151:26]
  wire  _GEN_1537 = igen_io_fire ? _GEN_513 : rob_ingress_id_0; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1538 = igen_io_fire ? _GEN_514 : rob_ingress_id_1; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1539 = igen_io_fire ? _GEN_515 : rob_ingress_id_2; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1540 = igen_io_fire ? _GEN_516 : rob_ingress_id_3; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1541 = igen_io_fire ? _GEN_517 : rob_ingress_id_4; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1542 = igen_io_fire ? _GEN_518 : rob_ingress_id_5; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1543 = igen_io_fire ? _GEN_519 : rob_ingress_id_6; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1544 = igen_io_fire ? _GEN_520 : rob_ingress_id_7; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1545 = igen_io_fire ? _GEN_521 : rob_ingress_id_8; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1546 = igen_io_fire ? _GEN_522 : rob_ingress_id_9; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1547 = igen_io_fire ? _GEN_523 : rob_ingress_id_10; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1548 = igen_io_fire ? _GEN_524 : rob_ingress_id_11; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1549 = igen_io_fire ? _GEN_525 : rob_ingress_id_12; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1550 = igen_io_fire ? _GEN_526 : rob_ingress_id_13; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1551 = igen_io_fire ? _GEN_527 : rob_ingress_id_14; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1552 = igen_io_fire ? _GEN_528 : rob_ingress_id_15; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1553 = igen_io_fire ? _GEN_529 : rob_ingress_id_16; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1554 = igen_io_fire ? _GEN_530 : rob_ingress_id_17; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1555 = igen_io_fire ? _GEN_531 : rob_ingress_id_18; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1556 = igen_io_fire ? _GEN_532 : rob_ingress_id_19; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1557 = igen_io_fire ? _GEN_533 : rob_ingress_id_20; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1558 = igen_io_fire ? _GEN_534 : rob_ingress_id_21; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1559 = igen_io_fire ? _GEN_535 : rob_ingress_id_22; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1560 = igen_io_fire ? _GEN_536 : rob_ingress_id_23; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1561 = igen_io_fire ? _GEN_537 : rob_ingress_id_24; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1562 = igen_io_fire ? _GEN_538 : rob_ingress_id_25; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1563 = igen_io_fire ? _GEN_539 : rob_ingress_id_26; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1564 = igen_io_fire ? _GEN_540 : rob_ingress_id_27; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1565 = igen_io_fire ? _GEN_541 : rob_ingress_id_28; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1566 = igen_io_fire ? _GEN_542 : rob_ingress_id_29; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1567 = igen_io_fire ? _GEN_543 : rob_ingress_id_30; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1568 = igen_io_fire ? _GEN_544 : rob_ingress_id_31; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1569 = igen_io_fire ? _GEN_545 : rob_ingress_id_32; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1570 = igen_io_fire ? _GEN_546 : rob_ingress_id_33; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1571 = igen_io_fire ? _GEN_547 : rob_ingress_id_34; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1572 = igen_io_fire ? _GEN_548 : rob_ingress_id_35; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1573 = igen_io_fire ? _GEN_549 : rob_ingress_id_36; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1574 = igen_io_fire ? _GEN_550 : rob_ingress_id_37; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1575 = igen_io_fire ? _GEN_551 : rob_ingress_id_38; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1576 = igen_io_fire ? _GEN_552 : rob_ingress_id_39; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1577 = igen_io_fire ? _GEN_553 : rob_ingress_id_40; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1578 = igen_io_fire ? _GEN_554 : rob_ingress_id_41; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1579 = igen_io_fire ? _GEN_555 : rob_ingress_id_42; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1580 = igen_io_fire ? _GEN_556 : rob_ingress_id_43; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1581 = igen_io_fire ? _GEN_557 : rob_ingress_id_44; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1582 = igen_io_fire ? _GEN_558 : rob_ingress_id_45; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1583 = igen_io_fire ? _GEN_559 : rob_ingress_id_46; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1584 = igen_io_fire ? _GEN_560 : rob_ingress_id_47; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1585 = igen_io_fire ? _GEN_561 : rob_ingress_id_48; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1586 = igen_io_fire ? _GEN_562 : rob_ingress_id_49; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1587 = igen_io_fire ? _GEN_563 : rob_ingress_id_50; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1588 = igen_io_fire ? _GEN_564 : rob_ingress_id_51; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1589 = igen_io_fire ? _GEN_565 : rob_ingress_id_52; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1590 = igen_io_fire ? _GEN_566 : rob_ingress_id_53; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1591 = igen_io_fire ? _GEN_567 : rob_ingress_id_54; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1592 = igen_io_fire ? _GEN_568 : rob_ingress_id_55; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1593 = igen_io_fire ? _GEN_569 : rob_ingress_id_56; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1594 = igen_io_fire ? _GEN_570 : rob_ingress_id_57; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1595 = igen_io_fire ? _GEN_571 : rob_ingress_id_58; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1596 = igen_io_fire ? _GEN_572 : rob_ingress_id_59; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1597 = igen_io_fire ? _GEN_573 : rob_ingress_id_60; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1598 = igen_io_fire ? _GEN_574 : rob_ingress_id_61; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1599 = igen_io_fire ? _GEN_575 : rob_ingress_id_62; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1600 = igen_io_fire ? _GEN_576 : rob_ingress_id_63; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1601 = igen_io_fire ? _GEN_577 : rob_ingress_id_64; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1602 = igen_io_fire ? _GEN_578 : rob_ingress_id_65; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1603 = igen_io_fire ? _GEN_579 : rob_ingress_id_66; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1604 = igen_io_fire ? _GEN_580 : rob_ingress_id_67; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1605 = igen_io_fire ? _GEN_581 : rob_ingress_id_68; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1606 = igen_io_fire ? _GEN_582 : rob_ingress_id_69; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1607 = igen_io_fire ? _GEN_583 : rob_ingress_id_70; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1608 = igen_io_fire ? _GEN_584 : rob_ingress_id_71; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1609 = igen_io_fire ? _GEN_585 : rob_ingress_id_72; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1610 = igen_io_fire ? _GEN_586 : rob_ingress_id_73; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1611 = igen_io_fire ? _GEN_587 : rob_ingress_id_74; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1612 = igen_io_fire ? _GEN_588 : rob_ingress_id_75; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1613 = igen_io_fire ? _GEN_589 : rob_ingress_id_76; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1614 = igen_io_fire ? _GEN_590 : rob_ingress_id_77; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1615 = igen_io_fire ? _GEN_591 : rob_ingress_id_78; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1616 = igen_io_fire ? _GEN_592 : rob_ingress_id_79; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1617 = igen_io_fire ? _GEN_593 : rob_ingress_id_80; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1618 = igen_io_fire ? _GEN_594 : rob_ingress_id_81; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1619 = igen_io_fire ? _GEN_595 : rob_ingress_id_82; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1620 = igen_io_fire ? _GEN_596 : rob_ingress_id_83; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1621 = igen_io_fire ? _GEN_597 : rob_ingress_id_84; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1622 = igen_io_fire ? _GEN_598 : rob_ingress_id_85; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1623 = igen_io_fire ? _GEN_599 : rob_ingress_id_86; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1624 = igen_io_fire ? _GEN_600 : rob_ingress_id_87; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1625 = igen_io_fire ? _GEN_601 : rob_ingress_id_88; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1626 = igen_io_fire ? _GEN_602 : rob_ingress_id_89; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1627 = igen_io_fire ? _GEN_603 : rob_ingress_id_90; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1628 = igen_io_fire ? _GEN_604 : rob_ingress_id_91; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1629 = igen_io_fire ? _GEN_605 : rob_ingress_id_92; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1630 = igen_io_fire ? _GEN_606 : rob_ingress_id_93; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1631 = igen_io_fire ? _GEN_607 : rob_ingress_id_94; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1632 = igen_io_fire ? _GEN_608 : rob_ingress_id_95; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1633 = igen_io_fire ? _GEN_609 : rob_ingress_id_96; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1634 = igen_io_fire ? _GEN_610 : rob_ingress_id_97; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1635 = igen_io_fire ? _GEN_611 : rob_ingress_id_98; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1636 = igen_io_fire ? _GEN_612 : rob_ingress_id_99; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1637 = igen_io_fire ? _GEN_613 : rob_ingress_id_100; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1638 = igen_io_fire ? _GEN_614 : rob_ingress_id_101; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1639 = igen_io_fire ? _GEN_615 : rob_ingress_id_102; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1640 = igen_io_fire ? _GEN_616 : rob_ingress_id_103; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1641 = igen_io_fire ? _GEN_617 : rob_ingress_id_104; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1642 = igen_io_fire ? _GEN_618 : rob_ingress_id_105; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1643 = igen_io_fire ? _GEN_619 : rob_ingress_id_106; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1644 = igen_io_fire ? _GEN_620 : rob_ingress_id_107; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1645 = igen_io_fire ? _GEN_621 : rob_ingress_id_108; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1646 = igen_io_fire ? _GEN_622 : rob_ingress_id_109; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1647 = igen_io_fire ? _GEN_623 : rob_ingress_id_110; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1648 = igen_io_fire ? _GEN_624 : rob_ingress_id_111; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1649 = igen_io_fire ? _GEN_625 : rob_ingress_id_112; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1650 = igen_io_fire ? _GEN_626 : rob_ingress_id_113; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1651 = igen_io_fire ? _GEN_627 : rob_ingress_id_114; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1652 = igen_io_fire ? _GEN_628 : rob_ingress_id_115; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1653 = igen_io_fire ? _GEN_629 : rob_ingress_id_116; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1654 = igen_io_fire ? _GEN_630 : rob_ingress_id_117; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1655 = igen_io_fire ? _GEN_631 : rob_ingress_id_118; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1656 = igen_io_fire ? _GEN_632 : rob_ingress_id_119; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1657 = igen_io_fire ? _GEN_633 : rob_ingress_id_120; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1658 = igen_io_fire ? _GEN_634 : rob_ingress_id_121; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1659 = igen_io_fire ? _GEN_635 : rob_ingress_id_122; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1660 = igen_io_fire ? _GEN_636 : rob_ingress_id_123; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1661 = igen_io_fire ? _GEN_637 : rob_ingress_id_124; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1662 = igen_io_fire ? _GEN_638 : rob_ingress_id_125; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1663 = igen_io_fire ? _GEN_639 : rob_ingress_id_126; // @[TestHarness.scala 178:25 152:27]
  wire  _GEN_1664 = igen_io_fire ? _GEN_640 : rob_ingress_id_127; // @[TestHarness.scala 178:25 152:27]
  wire [3:0] _GEN_1665 = igen_io_fire ? _GEN_641 : rob_n_flits_0; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1666 = igen_io_fire ? _GEN_642 : rob_n_flits_1; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1667 = igen_io_fire ? _GEN_643 : rob_n_flits_2; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1668 = igen_io_fire ? _GEN_644 : rob_n_flits_3; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1669 = igen_io_fire ? _GEN_645 : rob_n_flits_4; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1670 = igen_io_fire ? _GEN_646 : rob_n_flits_5; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1671 = igen_io_fire ? _GEN_647 : rob_n_flits_6; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1672 = igen_io_fire ? _GEN_648 : rob_n_flits_7; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1673 = igen_io_fire ? _GEN_649 : rob_n_flits_8; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1674 = igen_io_fire ? _GEN_650 : rob_n_flits_9; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1675 = igen_io_fire ? _GEN_651 : rob_n_flits_10; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1676 = igen_io_fire ? _GEN_652 : rob_n_flits_11; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1677 = igen_io_fire ? _GEN_653 : rob_n_flits_12; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1678 = igen_io_fire ? _GEN_654 : rob_n_flits_13; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1679 = igen_io_fire ? _GEN_655 : rob_n_flits_14; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1680 = igen_io_fire ? _GEN_656 : rob_n_flits_15; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1681 = igen_io_fire ? _GEN_657 : rob_n_flits_16; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1682 = igen_io_fire ? _GEN_658 : rob_n_flits_17; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1683 = igen_io_fire ? _GEN_659 : rob_n_flits_18; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1684 = igen_io_fire ? _GEN_660 : rob_n_flits_19; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1685 = igen_io_fire ? _GEN_661 : rob_n_flits_20; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1686 = igen_io_fire ? _GEN_662 : rob_n_flits_21; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1687 = igen_io_fire ? _GEN_663 : rob_n_flits_22; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1688 = igen_io_fire ? _GEN_664 : rob_n_flits_23; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1689 = igen_io_fire ? _GEN_665 : rob_n_flits_24; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1690 = igen_io_fire ? _GEN_666 : rob_n_flits_25; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1691 = igen_io_fire ? _GEN_667 : rob_n_flits_26; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1692 = igen_io_fire ? _GEN_668 : rob_n_flits_27; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1693 = igen_io_fire ? _GEN_669 : rob_n_flits_28; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1694 = igen_io_fire ? _GEN_670 : rob_n_flits_29; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1695 = igen_io_fire ? _GEN_671 : rob_n_flits_30; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1696 = igen_io_fire ? _GEN_672 : rob_n_flits_31; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1697 = igen_io_fire ? _GEN_673 : rob_n_flits_32; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1698 = igen_io_fire ? _GEN_674 : rob_n_flits_33; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1699 = igen_io_fire ? _GEN_675 : rob_n_flits_34; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1700 = igen_io_fire ? _GEN_676 : rob_n_flits_35; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1701 = igen_io_fire ? _GEN_677 : rob_n_flits_36; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1702 = igen_io_fire ? _GEN_678 : rob_n_flits_37; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1703 = igen_io_fire ? _GEN_679 : rob_n_flits_38; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1704 = igen_io_fire ? _GEN_680 : rob_n_flits_39; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1705 = igen_io_fire ? _GEN_681 : rob_n_flits_40; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1706 = igen_io_fire ? _GEN_682 : rob_n_flits_41; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1707 = igen_io_fire ? _GEN_683 : rob_n_flits_42; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1708 = igen_io_fire ? _GEN_684 : rob_n_flits_43; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1709 = igen_io_fire ? _GEN_685 : rob_n_flits_44; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1710 = igen_io_fire ? _GEN_686 : rob_n_flits_45; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1711 = igen_io_fire ? _GEN_687 : rob_n_flits_46; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1712 = igen_io_fire ? _GEN_688 : rob_n_flits_47; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1713 = igen_io_fire ? _GEN_689 : rob_n_flits_48; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1714 = igen_io_fire ? _GEN_690 : rob_n_flits_49; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1715 = igen_io_fire ? _GEN_691 : rob_n_flits_50; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1716 = igen_io_fire ? _GEN_692 : rob_n_flits_51; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1717 = igen_io_fire ? _GEN_693 : rob_n_flits_52; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1718 = igen_io_fire ? _GEN_694 : rob_n_flits_53; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1719 = igen_io_fire ? _GEN_695 : rob_n_flits_54; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1720 = igen_io_fire ? _GEN_696 : rob_n_flits_55; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1721 = igen_io_fire ? _GEN_697 : rob_n_flits_56; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1722 = igen_io_fire ? _GEN_698 : rob_n_flits_57; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1723 = igen_io_fire ? _GEN_699 : rob_n_flits_58; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1724 = igen_io_fire ? _GEN_700 : rob_n_flits_59; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1725 = igen_io_fire ? _GEN_701 : rob_n_flits_60; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1726 = igen_io_fire ? _GEN_702 : rob_n_flits_61; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1727 = igen_io_fire ? _GEN_703 : rob_n_flits_62; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1728 = igen_io_fire ? _GEN_704 : rob_n_flits_63; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1729 = igen_io_fire ? _GEN_705 : rob_n_flits_64; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1730 = igen_io_fire ? _GEN_706 : rob_n_flits_65; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1731 = igen_io_fire ? _GEN_707 : rob_n_flits_66; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1732 = igen_io_fire ? _GEN_708 : rob_n_flits_67; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1733 = igen_io_fire ? _GEN_709 : rob_n_flits_68; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1734 = igen_io_fire ? _GEN_710 : rob_n_flits_69; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1735 = igen_io_fire ? _GEN_711 : rob_n_flits_70; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1736 = igen_io_fire ? _GEN_712 : rob_n_flits_71; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1737 = igen_io_fire ? _GEN_713 : rob_n_flits_72; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1738 = igen_io_fire ? _GEN_714 : rob_n_flits_73; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1739 = igen_io_fire ? _GEN_715 : rob_n_flits_74; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1740 = igen_io_fire ? _GEN_716 : rob_n_flits_75; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1741 = igen_io_fire ? _GEN_717 : rob_n_flits_76; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1742 = igen_io_fire ? _GEN_718 : rob_n_flits_77; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1743 = igen_io_fire ? _GEN_719 : rob_n_flits_78; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1744 = igen_io_fire ? _GEN_720 : rob_n_flits_79; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1745 = igen_io_fire ? _GEN_721 : rob_n_flits_80; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1746 = igen_io_fire ? _GEN_722 : rob_n_flits_81; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1747 = igen_io_fire ? _GEN_723 : rob_n_flits_82; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1748 = igen_io_fire ? _GEN_724 : rob_n_flits_83; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1749 = igen_io_fire ? _GEN_725 : rob_n_flits_84; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1750 = igen_io_fire ? _GEN_726 : rob_n_flits_85; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1751 = igen_io_fire ? _GEN_727 : rob_n_flits_86; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1752 = igen_io_fire ? _GEN_728 : rob_n_flits_87; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1753 = igen_io_fire ? _GEN_729 : rob_n_flits_88; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1754 = igen_io_fire ? _GEN_730 : rob_n_flits_89; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1755 = igen_io_fire ? _GEN_731 : rob_n_flits_90; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1756 = igen_io_fire ? _GEN_732 : rob_n_flits_91; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1757 = igen_io_fire ? _GEN_733 : rob_n_flits_92; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1758 = igen_io_fire ? _GEN_734 : rob_n_flits_93; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1759 = igen_io_fire ? _GEN_735 : rob_n_flits_94; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1760 = igen_io_fire ? _GEN_736 : rob_n_flits_95; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1761 = igen_io_fire ? _GEN_737 : rob_n_flits_96; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1762 = igen_io_fire ? _GEN_738 : rob_n_flits_97; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1763 = igen_io_fire ? _GEN_739 : rob_n_flits_98; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1764 = igen_io_fire ? _GEN_740 : rob_n_flits_99; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1765 = igen_io_fire ? _GEN_741 : rob_n_flits_100; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1766 = igen_io_fire ? _GEN_742 : rob_n_flits_101; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1767 = igen_io_fire ? _GEN_743 : rob_n_flits_102; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1768 = igen_io_fire ? _GEN_744 : rob_n_flits_103; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1769 = igen_io_fire ? _GEN_745 : rob_n_flits_104; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1770 = igen_io_fire ? _GEN_746 : rob_n_flits_105; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1771 = igen_io_fire ? _GEN_747 : rob_n_flits_106; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1772 = igen_io_fire ? _GEN_748 : rob_n_flits_107; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1773 = igen_io_fire ? _GEN_749 : rob_n_flits_108; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1774 = igen_io_fire ? _GEN_750 : rob_n_flits_109; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1775 = igen_io_fire ? _GEN_751 : rob_n_flits_110; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1776 = igen_io_fire ? _GEN_752 : rob_n_flits_111; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1777 = igen_io_fire ? _GEN_753 : rob_n_flits_112; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1778 = igen_io_fire ? _GEN_754 : rob_n_flits_113; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1779 = igen_io_fire ? _GEN_755 : rob_n_flits_114; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1780 = igen_io_fire ? _GEN_756 : rob_n_flits_115; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1781 = igen_io_fire ? _GEN_757 : rob_n_flits_116; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1782 = igen_io_fire ? _GEN_758 : rob_n_flits_117; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1783 = igen_io_fire ? _GEN_759 : rob_n_flits_118; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1784 = igen_io_fire ? _GEN_760 : rob_n_flits_119; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1785 = igen_io_fire ? _GEN_761 : rob_n_flits_120; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1786 = igen_io_fire ? _GEN_762 : rob_n_flits_121; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1787 = igen_io_fire ? _GEN_763 : rob_n_flits_122; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1788 = igen_io_fire ? _GEN_764 : rob_n_flits_123; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1789 = igen_io_fire ? _GEN_765 : rob_n_flits_124; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1790 = igen_io_fire ? _GEN_766 : rob_n_flits_125; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1791 = igen_io_fire ? _GEN_767 : rob_n_flits_126; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1792 = igen_io_fire ? _GEN_768 : rob_n_flits_127; // @[TestHarness.scala 153:24 178:25]
  wire [3:0] _GEN_1793 = igen_io_fire ? _GEN_769 : rob_flits_returned_0; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1794 = igen_io_fire ? _GEN_770 : rob_flits_returned_1; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1795 = igen_io_fire ? _GEN_771 : rob_flits_returned_2; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1796 = igen_io_fire ? _GEN_772 : rob_flits_returned_3; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1797 = igen_io_fire ? _GEN_773 : rob_flits_returned_4; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1798 = igen_io_fire ? _GEN_774 : rob_flits_returned_5; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1799 = igen_io_fire ? _GEN_775 : rob_flits_returned_6; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1800 = igen_io_fire ? _GEN_776 : rob_flits_returned_7; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1801 = igen_io_fire ? _GEN_777 : rob_flits_returned_8; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1802 = igen_io_fire ? _GEN_778 : rob_flits_returned_9; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1803 = igen_io_fire ? _GEN_779 : rob_flits_returned_10; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1804 = igen_io_fire ? _GEN_780 : rob_flits_returned_11; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1805 = igen_io_fire ? _GEN_781 : rob_flits_returned_12; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1806 = igen_io_fire ? _GEN_782 : rob_flits_returned_13; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1807 = igen_io_fire ? _GEN_783 : rob_flits_returned_14; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1808 = igen_io_fire ? _GEN_784 : rob_flits_returned_15; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1809 = igen_io_fire ? _GEN_785 : rob_flits_returned_16; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1810 = igen_io_fire ? _GEN_786 : rob_flits_returned_17; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1811 = igen_io_fire ? _GEN_787 : rob_flits_returned_18; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1812 = igen_io_fire ? _GEN_788 : rob_flits_returned_19; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1813 = igen_io_fire ? _GEN_789 : rob_flits_returned_20; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1814 = igen_io_fire ? _GEN_790 : rob_flits_returned_21; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1815 = igen_io_fire ? _GEN_791 : rob_flits_returned_22; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1816 = igen_io_fire ? _GEN_792 : rob_flits_returned_23; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1817 = igen_io_fire ? _GEN_793 : rob_flits_returned_24; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1818 = igen_io_fire ? _GEN_794 : rob_flits_returned_25; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1819 = igen_io_fire ? _GEN_795 : rob_flits_returned_26; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1820 = igen_io_fire ? _GEN_796 : rob_flits_returned_27; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1821 = igen_io_fire ? _GEN_797 : rob_flits_returned_28; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1822 = igen_io_fire ? _GEN_798 : rob_flits_returned_29; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1823 = igen_io_fire ? _GEN_799 : rob_flits_returned_30; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1824 = igen_io_fire ? _GEN_800 : rob_flits_returned_31; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1825 = igen_io_fire ? _GEN_801 : rob_flits_returned_32; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1826 = igen_io_fire ? _GEN_802 : rob_flits_returned_33; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1827 = igen_io_fire ? _GEN_803 : rob_flits_returned_34; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1828 = igen_io_fire ? _GEN_804 : rob_flits_returned_35; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1829 = igen_io_fire ? _GEN_805 : rob_flits_returned_36; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1830 = igen_io_fire ? _GEN_806 : rob_flits_returned_37; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1831 = igen_io_fire ? _GEN_807 : rob_flits_returned_38; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1832 = igen_io_fire ? _GEN_808 : rob_flits_returned_39; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1833 = igen_io_fire ? _GEN_809 : rob_flits_returned_40; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1834 = igen_io_fire ? _GEN_810 : rob_flits_returned_41; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1835 = igen_io_fire ? _GEN_811 : rob_flits_returned_42; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1836 = igen_io_fire ? _GEN_812 : rob_flits_returned_43; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1837 = igen_io_fire ? _GEN_813 : rob_flits_returned_44; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1838 = igen_io_fire ? _GEN_814 : rob_flits_returned_45; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1839 = igen_io_fire ? _GEN_815 : rob_flits_returned_46; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1840 = igen_io_fire ? _GEN_816 : rob_flits_returned_47; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1841 = igen_io_fire ? _GEN_817 : rob_flits_returned_48; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1842 = igen_io_fire ? _GEN_818 : rob_flits_returned_49; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1843 = igen_io_fire ? _GEN_819 : rob_flits_returned_50; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1844 = igen_io_fire ? _GEN_820 : rob_flits_returned_51; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1845 = igen_io_fire ? _GEN_821 : rob_flits_returned_52; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1846 = igen_io_fire ? _GEN_822 : rob_flits_returned_53; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1847 = igen_io_fire ? _GEN_823 : rob_flits_returned_54; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1848 = igen_io_fire ? _GEN_824 : rob_flits_returned_55; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1849 = igen_io_fire ? _GEN_825 : rob_flits_returned_56; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1850 = igen_io_fire ? _GEN_826 : rob_flits_returned_57; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1851 = igen_io_fire ? _GEN_827 : rob_flits_returned_58; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1852 = igen_io_fire ? _GEN_828 : rob_flits_returned_59; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1853 = igen_io_fire ? _GEN_829 : rob_flits_returned_60; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1854 = igen_io_fire ? _GEN_830 : rob_flits_returned_61; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1855 = igen_io_fire ? _GEN_831 : rob_flits_returned_62; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1856 = igen_io_fire ? _GEN_832 : rob_flits_returned_63; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1857 = igen_io_fire ? _GEN_833 : rob_flits_returned_64; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1858 = igen_io_fire ? _GEN_834 : rob_flits_returned_65; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1859 = igen_io_fire ? _GEN_835 : rob_flits_returned_66; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1860 = igen_io_fire ? _GEN_836 : rob_flits_returned_67; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1861 = igen_io_fire ? _GEN_837 : rob_flits_returned_68; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1862 = igen_io_fire ? _GEN_838 : rob_flits_returned_69; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1863 = igen_io_fire ? _GEN_839 : rob_flits_returned_70; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1864 = igen_io_fire ? _GEN_840 : rob_flits_returned_71; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1865 = igen_io_fire ? _GEN_841 : rob_flits_returned_72; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1866 = igen_io_fire ? _GEN_842 : rob_flits_returned_73; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1867 = igen_io_fire ? _GEN_843 : rob_flits_returned_74; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1868 = igen_io_fire ? _GEN_844 : rob_flits_returned_75; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1869 = igen_io_fire ? _GEN_845 : rob_flits_returned_76; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1870 = igen_io_fire ? _GEN_846 : rob_flits_returned_77; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1871 = igen_io_fire ? _GEN_847 : rob_flits_returned_78; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1872 = igen_io_fire ? _GEN_848 : rob_flits_returned_79; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1873 = igen_io_fire ? _GEN_849 : rob_flits_returned_80; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1874 = igen_io_fire ? _GEN_850 : rob_flits_returned_81; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1875 = igen_io_fire ? _GEN_851 : rob_flits_returned_82; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1876 = igen_io_fire ? _GEN_852 : rob_flits_returned_83; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1877 = igen_io_fire ? _GEN_853 : rob_flits_returned_84; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1878 = igen_io_fire ? _GEN_854 : rob_flits_returned_85; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1879 = igen_io_fire ? _GEN_855 : rob_flits_returned_86; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1880 = igen_io_fire ? _GEN_856 : rob_flits_returned_87; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1881 = igen_io_fire ? _GEN_857 : rob_flits_returned_88; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1882 = igen_io_fire ? _GEN_858 : rob_flits_returned_89; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1883 = igen_io_fire ? _GEN_859 : rob_flits_returned_90; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1884 = igen_io_fire ? _GEN_860 : rob_flits_returned_91; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1885 = igen_io_fire ? _GEN_861 : rob_flits_returned_92; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1886 = igen_io_fire ? _GEN_862 : rob_flits_returned_93; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1887 = igen_io_fire ? _GEN_863 : rob_flits_returned_94; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1888 = igen_io_fire ? _GEN_864 : rob_flits_returned_95; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1889 = igen_io_fire ? _GEN_865 : rob_flits_returned_96; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1890 = igen_io_fire ? _GEN_866 : rob_flits_returned_97; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1891 = igen_io_fire ? _GEN_867 : rob_flits_returned_98; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1892 = igen_io_fire ? _GEN_868 : rob_flits_returned_99; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1893 = igen_io_fire ? _GEN_869 : rob_flits_returned_100; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1894 = igen_io_fire ? _GEN_870 : rob_flits_returned_101; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1895 = igen_io_fire ? _GEN_871 : rob_flits_returned_102; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1896 = igen_io_fire ? _GEN_872 : rob_flits_returned_103; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1897 = igen_io_fire ? _GEN_873 : rob_flits_returned_104; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1898 = igen_io_fire ? _GEN_874 : rob_flits_returned_105; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1899 = igen_io_fire ? _GEN_875 : rob_flits_returned_106; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1900 = igen_io_fire ? _GEN_876 : rob_flits_returned_107; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1901 = igen_io_fire ? _GEN_877 : rob_flits_returned_108; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1902 = igen_io_fire ? _GEN_878 : rob_flits_returned_109; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1903 = igen_io_fire ? _GEN_879 : rob_flits_returned_110; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1904 = igen_io_fire ? _GEN_880 : rob_flits_returned_111; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1905 = igen_io_fire ? _GEN_881 : rob_flits_returned_112; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1906 = igen_io_fire ? _GEN_882 : rob_flits_returned_113; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1907 = igen_io_fire ? _GEN_883 : rob_flits_returned_114; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1908 = igen_io_fire ? _GEN_884 : rob_flits_returned_115; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1909 = igen_io_fire ? _GEN_885 : rob_flits_returned_116; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1910 = igen_io_fire ? _GEN_886 : rob_flits_returned_117; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1911 = igen_io_fire ? _GEN_887 : rob_flits_returned_118; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1912 = igen_io_fire ? _GEN_888 : rob_flits_returned_119; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1913 = igen_io_fire ? _GEN_889 : rob_flits_returned_120; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1914 = igen_io_fire ? _GEN_890 : rob_flits_returned_121; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1915 = igen_io_fire ? _GEN_891 : rob_flits_returned_122; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1916 = igen_io_fire ? _GEN_892 : rob_flits_returned_123; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1917 = igen_io_fire ? _GEN_893 : rob_flits_returned_124; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1918 = igen_io_fire ? _GEN_894 : rob_flits_returned_125; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1919 = igen_io_fire ? _GEN_895 : rob_flits_returned_126; // @[TestHarness.scala 178:25 154:31]
  wire [3:0] _GEN_1920 = igen_io_fire ? _GEN_896 : rob_flits_returned_127; // @[TestHarness.scala 178:25 154:31]
  wire [63:0] _GEN_1921 = igen_io_fire ? _GEN_897 : rob_tscs_0; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1922 = igen_io_fire ? _GEN_898 : rob_tscs_1; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1923 = igen_io_fire ? _GEN_899 : rob_tscs_2; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1924 = igen_io_fire ? _GEN_900 : rob_tscs_3; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1925 = igen_io_fire ? _GEN_901 : rob_tscs_4; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1926 = igen_io_fire ? _GEN_902 : rob_tscs_5; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1927 = igen_io_fire ? _GEN_903 : rob_tscs_6; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1928 = igen_io_fire ? _GEN_904 : rob_tscs_7; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1929 = igen_io_fire ? _GEN_905 : rob_tscs_8; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1930 = igen_io_fire ? _GEN_906 : rob_tscs_9; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1931 = igen_io_fire ? _GEN_907 : rob_tscs_10; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1932 = igen_io_fire ? _GEN_908 : rob_tscs_11; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1933 = igen_io_fire ? _GEN_909 : rob_tscs_12; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1934 = igen_io_fire ? _GEN_910 : rob_tscs_13; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1935 = igen_io_fire ? _GEN_911 : rob_tscs_14; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1936 = igen_io_fire ? _GEN_912 : rob_tscs_15; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1937 = igen_io_fire ? _GEN_913 : rob_tscs_16; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1938 = igen_io_fire ? _GEN_914 : rob_tscs_17; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1939 = igen_io_fire ? _GEN_915 : rob_tscs_18; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1940 = igen_io_fire ? _GEN_916 : rob_tscs_19; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1941 = igen_io_fire ? _GEN_917 : rob_tscs_20; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1942 = igen_io_fire ? _GEN_918 : rob_tscs_21; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1943 = igen_io_fire ? _GEN_919 : rob_tscs_22; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1944 = igen_io_fire ? _GEN_920 : rob_tscs_23; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1945 = igen_io_fire ? _GEN_921 : rob_tscs_24; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1946 = igen_io_fire ? _GEN_922 : rob_tscs_25; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1947 = igen_io_fire ? _GEN_923 : rob_tscs_26; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1948 = igen_io_fire ? _GEN_924 : rob_tscs_27; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1949 = igen_io_fire ? _GEN_925 : rob_tscs_28; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1950 = igen_io_fire ? _GEN_926 : rob_tscs_29; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1951 = igen_io_fire ? _GEN_927 : rob_tscs_30; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1952 = igen_io_fire ? _GEN_928 : rob_tscs_31; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1953 = igen_io_fire ? _GEN_929 : rob_tscs_32; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1954 = igen_io_fire ? _GEN_930 : rob_tscs_33; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1955 = igen_io_fire ? _GEN_931 : rob_tscs_34; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1956 = igen_io_fire ? _GEN_932 : rob_tscs_35; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1957 = igen_io_fire ? _GEN_933 : rob_tscs_36; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1958 = igen_io_fire ? _GEN_934 : rob_tscs_37; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1959 = igen_io_fire ? _GEN_935 : rob_tscs_38; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1960 = igen_io_fire ? _GEN_936 : rob_tscs_39; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1961 = igen_io_fire ? _GEN_937 : rob_tscs_40; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1962 = igen_io_fire ? _GEN_938 : rob_tscs_41; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1963 = igen_io_fire ? _GEN_939 : rob_tscs_42; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1964 = igen_io_fire ? _GEN_940 : rob_tscs_43; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1965 = igen_io_fire ? _GEN_941 : rob_tscs_44; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1966 = igen_io_fire ? _GEN_942 : rob_tscs_45; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1967 = igen_io_fire ? _GEN_943 : rob_tscs_46; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1968 = igen_io_fire ? _GEN_944 : rob_tscs_47; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1969 = igen_io_fire ? _GEN_945 : rob_tscs_48; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1970 = igen_io_fire ? _GEN_946 : rob_tscs_49; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1971 = igen_io_fire ? _GEN_947 : rob_tscs_50; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1972 = igen_io_fire ? _GEN_948 : rob_tscs_51; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1973 = igen_io_fire ? _GEN_949 : rob_tscs_52; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1974 = igen_io_fire ? _GEN_950 : rob_tscs_53; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1975 = igen_io_fire ? _GEN_951 : rob_tscs_54; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1976 = igen_io_fire ? _GEN_952 : rob_tscs_55; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1977 = igen_io_fire ? _GEN_953 : rob_tscs_56; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1978 = igen_io_fire ? _GEN_954 : rob_tscs_57; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1979 = igen_io_fire ? _GEN_955 : rob_tscs_58; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1980 = igen_io_fire ? _GEN_956 : rob_tscs_59; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1981 = igen_io_fire ? _GEN_957 : rob_tscs_60; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1982 = igen_io_fire ? _GEN_958 : rob_tscs_61; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1983 = igen_io_fire ? _GEN_959 : rob_tscs_62; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1984 = igen_io_fire ? _GEN_960 : rob_tscs_63; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1985 = igen_io_fire ? _GEN_961 : rob_tscs_64; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1986 = igen_io_fire ? _GEN_962 : rob_tscs_65; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1987 = igen_io_fire ? _GEN_963 : rob_tscs_66; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1988 = igen_io_fire ? _GEN_964 : rob_tscs_67; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1989 = igen_io_fire ? _GEN_965 : rob_tscs_68; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1990 = igen_io_fire ? _GEN_966 : rob_tscs_69; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1991 = igen_io_fire ? _GEN_967 : rob_tscs_70; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1992 = igen_io_fire ? _GEN_968 : rob_tscs_71; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1993 = igen_io_fire ? _GEN_969 : rob_tscs_72; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1994 = igen_io_fire ? _GEN_970 : rob_tscs_73; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1995 = igen_io_fire ? _GEN_971 : rob_tscs_74; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1996 = igen_io_fire ? _GEN_972 : rob_tscs_75; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1997 = igen_io_fire ? _GEN_973 : rob_tscs_76; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1998 = igen_io_fire ? _GEN_974 : rob_tscs_77; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_1999 = igen_io_fire ? _GEN_975 : rob_tscs_78; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2000 = igen_io_fire ? _GEN_976 : rob_tscs_79; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2001 = igen_io_fire ? _GEN_977 : rob_tscs_80; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2002 = igen_io_fire ? _GEN_978 : rob_tscs_81; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2003 = igen_io_fire ? _GEN_979 : rob_tscs_82; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2004 = igen_io_fire ? _GEN_980 : rob_tscs_83; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2005 = igen_io_fire ? _GEN_981 : rob_tscs_84; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2006 = igen_io_fire ? _GEN_982 : rob_tscs_85; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2007 = igen_io_fire ? _GEN_983 : rob_tscs_86; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2008 = igen_io_fire ? _GEN_984 : rob_tscs_87; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2009 = igen_io_fire ? _GEN_985 : rob_tscs_88; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2010 = igen_io_fire ? _GEN_986 : rob_tscs_89; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2011 = igen_io_fire ? _GEN_987 : rob_tscs_90; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2012 = igen_io_fire ? _GEN_988 : rob_tscs_91; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2013 = igen_io_fire ? _GEN_989 : rob_tscs_92; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2014 = igen_io_fire ? _GEN_990 : rob_tscs_93; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2015 = igen_io_fire ? _GEN_991 : rob_tscs_94; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2016 = igen_io_fire ? _GEN_992 : rob_tscs_95; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2017 = igen_io_fire ? _GEN_993 : rob_tscs_96; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2018 = igen_io_fire ? _GEN_994 : rob_tscs_97; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2019 = igen_io_fire ? _GEN_995 : rob_tscs_98; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2020 = igen_io_fire ? _GEN_996 : rob_tscs_99; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2021 = igen_io_fire ? _GEN_997 : rob_tscs_100; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2022 = igen_io_fire ? _GEN_998 : rob_tscs_101; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2023 = igen_io_fire ? _GEN_999 : rob_tscs_102; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2024 = igen_io_fire ? _GEN_1000 : rob_tscs_103; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2025 = igen_io_fire ? _GEN_1001 : rob_tscs_104; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2026 = igen_io_fire ? _GEN_1002 : rob_tscs_105; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2027 = igen_io_fire ? _GEN_1003 : rob_tscs_106; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2028 = igen_io_fire ? _GEN_1004 : rob_tscs_107; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2029 = igen_io_fire ? _GEN_1005 : rob_tscs_108; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2030 = igen_io_fire ? _GEN_1006 : rob_tscs_109; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2031 = igen_io_fire ? _GEN_1007 : rob_tscs_110; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2032 = igen_io_fire ? _GEN_1008 : rob_tscs_111; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2033 = igen_io_fire ? _GEN_1009 : rob_tscs_112; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2034 = igen_io_fire ? _GEN_1010 : rob_tscs_113; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2035 = igen_io_fire ? _GEN_1011 : rob_tscs_114; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2036 = igen_io_fire ? _GEN_1012 : rob_tscs_115; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2037 = igen_io_fire ? _GEN_1013 : rob_tscs_116; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2038 = igen_io_fire ? _GEN_1014 : rob_tscs_117; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2039 = igen_io_fire ? _GEN_1015 : rob_tscs_118; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2040 = igen_io_fire ? _GEN_1016 : rob_tscs_119; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2041 = igen_io_fire ? _GEN_1017 : rob_tscs_120; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2042 = igen_io_fire ? _GEN_1018 : rob_tscs_121; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2043 = igen_io_fire ? _GEN_1019 : rob_tscs_122; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2044 = igen_io_fire ? _GEN_1020 : rob_tscs_123; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2045 = igen_io_fire ? _GEN_1021 : rob_tscs_124; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2046 = igen_io_fire ? _GEN_1022 : rob_tscs_125; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2047 = igen_io_fire ? _GEN_1023 : rob_tscs_126; // @[TestHarness.scala 155:21 178:25]
  wire [63:0] _GEN_2048 = igen_io_fire ? _GEN_1024 : rob_tscs_127; // @[TestHarness.scala 155:21 178:25]
  wire  _igen_io_rob_ready_T_7 = rob_alloc_avail_1 & rob_alloc_fires_1 & _igen_io_rob_ready_T_1; // @[TestHarness.scala 174:72]
  wire [63:0] _rob_payload_WIRE_3 = igen_1_io_out_bits_payload; // @[TestHarness.scala 179:{72,72}]
  wire [15:0] _GEN_2305 = 7'h0 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1281; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2306 = 7'h1 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1282; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2307 = 7'h2 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1283; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2308 = 7'h3 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1284; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2309 = 7'h4 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1285; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2310 = 7'h5 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1286; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2311 = 7'h6 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1287; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2312 = 7'h7 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1288; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2313 = 7'h8 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1289; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2314 = 7'h9 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1290; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2315 = 7'ha == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1291; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2316 = 7'hb == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1292; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2317 = 7'hc == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1293; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2318 = 7'hd == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1294; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2319 = 7'he == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1295; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2320 = 7'hf == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1296; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2321 = 7'h10 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1297; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2322 = 7'h11 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1298; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2323 = 7'h12 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1299; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2324 = 7'h13 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1300; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2325 = 7'h14 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1301; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2326 = 7'h15 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1302; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2327 = 7'h16 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1303; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2328 = 7'h17 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1304; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2329 = 7'h18 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1305; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2330 = 7'h19 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1306; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2331 = 7'h1a == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1307; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2332 = 7'h1b == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1308; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2333 = 7'h1c == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1309; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2334 = 7'h1d == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1310; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2335 = 7'h1e == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1311; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2336 = 7'h1f == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1312; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2337 = 7'h20 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1313; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2338 = 7'h21 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1314; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2339 = 7'h22 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1315; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2340 = 7'h23 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1316; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2341 = 7'h24 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1317; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2342 = 7'h25 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1318; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2343 = 7'h26 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1319; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2344 = 7'h27 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1320; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2345 = 7'h28 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1321; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2346 = 7'h29 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1322; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2347 = 7'h2a == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1323; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2348 = 7'h2b == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1324; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2349 = 7'h2c == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1325; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2350 = 7'h2d == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1326; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2351 = 7'h2e == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1327; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2352 = 7'h2f == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1328; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2353 = 7'h30 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1329; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2354 = 7'h31 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1330; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2355 = 7'h32 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1331; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2356 = 7'h33 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1332; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2357 = 7'h34 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1333; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2358 = 7'h35 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1334; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2359 = 7'h36 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1335; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2360 = 7'h37 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1336; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2361 = 7'h38 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1337; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2362 = 7'h39 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1338; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2363 = 7'h3a == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1339; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2364 = 7'h3b == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1340; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2365 = 7'h3c == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1341; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2366 = 7'h3d == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1342; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2367 = 7'h3e == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1343; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2368 = 7'h3f == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1344; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2369 = 7'h40 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1345; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2370 = 7'h41 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1346; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2371 = 7'h42 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1347; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2372 = 7'h43 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1348; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2373 = 7'h44 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1349; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2374 = 7'h45 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1350; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2375 = 7'h46 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1351; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2376 = 7'h47 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1352; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2377 = 7'h48 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1353; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2378 = 7'h49 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1354; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2379 = 7'h4a == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1355; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2380 = 7'h4b == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1356; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2381 = 7'h4c == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1357; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2382 = 7'h4d == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1358; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2383 = 7'h4e == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1359; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2384 = 7'h4f == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1360; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2385 = 7'h50 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1361; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2386 = 7'h51 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1362; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2387 = 7'h52 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1363; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2388 = 7'h53 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1364; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2389 = 7'h54 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1365; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2390 = 7'h55 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1366; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2391 = 7'h56 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1367; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2392 = 7'h57 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1368; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2393 = 7'h58 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1369; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2394 = 7'h59 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1370; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2395 = 7'h5a == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1371; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2396 = 7'h5b == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1372; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2397 = 7'h5c == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1373; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2398 = 7'h5d == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1374; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2399 = 7'h5e == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1375; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2400 = 7'h5f == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1376; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2401 = 7'h60 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1377; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2402 = 7'h61 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1378; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2403 = 7'h62 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1379; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2404 = 7'h63 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1380; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2405 = 7'h64 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1381; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2406 = 7'h65 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1382; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2407 = 7'h66 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1383; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2408 = 7'h67 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1384; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2409 = 7'h68 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1385; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2410 = 7'h69 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1386; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2411 = 7'h6a == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1387; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2412 = 7'h6b == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1388; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2413 = 7'h6c == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1389; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2414 = 7'h6d == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1390; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2415 = 7'h6e == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1391; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2416 = 7'h6f == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1392; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2417 = 7'h70 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1393; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2418 = 7'h71 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1394; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2419 = 7'h72 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1395; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2420 = 7'h73 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1396; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2421 = 7'h74 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1397; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2422 = 7'h75 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1398; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2423 = 7'h76 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1399; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2424 = 7'h77 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1400; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2425 = 7'h78 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1401; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2426 = 7'h79 == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1402; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2427 = 7'h7a == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1403; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2428 = 7'h7b == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1404; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2429 = 7'h7c == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1405; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2430 = 7'h7d == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1406; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2431 = 7'h7e == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1407; // @[TestHarness.scala 179:{36,36}]
  wire [15:0] _GEN_2432 = 7'h7f == rob_alloc_ids_1 ? _rob_payload_WIRE_3[15:0] : _GEN_1408; // @[TestHarness.scala 179:{36,36}]
  wire  _GEN_2561 = 7'h0 == rob_alloc_ids_1 | _GEN_1537; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2562 = 7'h1 == rob_alloc_ids_1 | _GEN_1538; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2563 = 7'h2 == rob_alloc_ids_1 | _GEN_1539; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2564 = 7'h3 == rob_alloc_ids_1 | _GEN_1540; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2565 = 7'h4 == rob_alloc_ids_1 | _GEN_1541; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2566 = 7'h5 == rob_alloc_ids_1 | _GEN_1542; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2567 = 7'h6 == rob_alloc_ids_1 | _GEN_1543; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2568 = 7'h7 == rob_alloc_ids_1 | _GEN_1544; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2569 = 7'h8 == rob_alloc_ids_1 | _GEN_1545; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2570 = 7'h9 == rob_alloc_ids_1 | _GEN_1546; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2571 = 7'ha == rob_alloc_ids_1 | _GEN_1547; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2572 = 7'hb == rob_alloc_ids_1 | _GEN_1548; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2573 = 7'hc == rob_alloc_ids_1 | _GEN_1549; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2574 = 7'hd == rob_alloc_ids_1 | _GEN_1550; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2575 = 7'he == rob_alloc_ids_1 | _GEN_1551; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2576 = 7'hf == rob_alloc_ids_1 | _GEN_1552; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2577 = 7'h10 == rob_alloc_ids_1 | _GEN_1553; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2578 = 7'h11 == rob_alloc_ids_1 | _GEN_1554; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2579 = 7'h12 == rob_alloc_ids_1 | _GEN_1555; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2580 = 7'h13 == rob_alloc_ids_1 | _GEN_1556; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2581 = 7'h14 == rob_alloc_ids_1 | _GEN_1557; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2582 = 7'h15 == rob_alloc_ids_1 | _GEN_1558; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2583 = 7'h16 == rob_alloc_ids_1 | _GEN_1559; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2584 = 7'h17 == rob_alloc_ids_1 | _GEN_1560; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2585 = 7'h18 == rob_alloc_ids_1 | _GEN_1561; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2586 = 7'h19 == rob_alloc_ids_1 | _GEN_1562; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2587 = 7'h1a == rob_alloc_ids_1 | _GEN_1563; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2588 = 7'h1b == rob_alloc_ids_1 | _GEN_1564; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2589 = 7'h1c == rob_alloc_ids_1 | _GEN_1565; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2590 = 7'h1d == rob_alloc_ids_1 | _GEN_1566; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2591 = 7'h1e == rob_alloc_ids_1 | _GEN_1567; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2592 = 7'h1f == rob_alloc_ids_1 | _GEN_1568; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2593 = 7'h20 == rob_alloc_ids_1 | _GEN_1569; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2594 = 7'h21 == rob_alloc_ids_1 | _GEN_1570; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2595 = 7'h22 == rob_alloc_ids_1 | _GEN_1571; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2596 = 7'h23 == rob_alloc_ids_1 | _GEN_1572; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2597 = 7'h24 == rob_alloc_ids_1 | _GEN_1573; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2598 = 7'h25 == rob_alloc_ids_1 | _GEN_1574; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2599 = 7'h26 == rob_alloc_ids_1 | _GEN_1575; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2600 = 7'h27 == rob_alloc_ids_1 | _GEN_1576; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2601 = 7'h28 == rob_alloc_ids_1 | _GEN_1577; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2602 = 7'h29 == rob_alloc_ids_1 | _GEN_1578; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2603 = 7'h2a == rob_alloc_ids_1 | _GEN_1579; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2604 = 7'h2b == rob_alloc_ids_1 | _GEN_1580; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2605 = 7'h2c == rob_alloc_ids_1 | _GEN_1581; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2606 = 7'h2d == rob_alloc_ids_1 | _GEN_1582; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2607 = 7'h2e == rob_alloc_ids_1 | _GEN_1583; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2608 = 7'h2f == rob_alloc_ids_1 | _GEN_1584; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2609 = 7'h30 == rob_alloc_ids_1 | _GEN_1585; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2610 = 7'h31 == rob_alloc_ids_1 | _GEN_1586; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2611 = 7'h32 == rob_alloc_ids_1 | _GEN_1587; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2612 = 7'h33 == rob_alloc_ids_1 | _GEN_1588; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2613 = 7'h34 == rob_alloc_ids_1 | _GEN_1589; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2614 = 7'h35 == rob_alloc_ids_1 | _GEN_1590; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2615 = 7'h36 == rob_alloc_ids_1 | _GEN_1591; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2616 = 7'h37 == rob_alloc_ids_1 | _GEN_1592; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2617 = 7'h38 == rob_alloc_ids_1 | _GEN_1593; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2618 = 7'h39 == rob_alloc_ids_1 | _GEN_1594; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2619 = 7'h3a == rob_alloc_ids_1 | _GEN_1595; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2620 = 7'h3b == rob_alloc_ids_1 | _GEN_1596; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2621 = 7'h3c == rob_alloc_ids_1 | _GEN_1597; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2622 = 7'h3d == rob_alloc_ids_1 | _GEN_1598; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2623 = 7'h3e == rob_alloc_ids_1 | _GEN_1599; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2624 = 7'h3f == rob_alloc_ids_1 | _GEN_1600; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2625 = 7'h40 == rob_alloc_ids_1 | _GEN_1601; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2626 = 7'h41 == rob_alloc_ids_1 | _GEN_1602; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2627 = 7'h42 == rob_alloc_ids_1 | _GEN_1603; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2628 = 7'h43 == rob_alloc_ids_1 | _GEN_1604; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2629 = 7'h44 == rob_alloc_ids_1 | _GEN_1605; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2630 = 7'h45 == rob_alloc_ids_1 | _GEN_1606; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2631 = 7'h46 == rob_alloc_ids_1 | _GEN_1607; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2632 = 7'h47 == rob_alloc_ids_1 | _GEN_1608; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2633 = 7'h48 == rob_alloc_ids_1 | _GEN_1609; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2634 = 7'h49 == rob_alloc_ids_1 | _GEN_1610; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2635 = 7'h4a == rob_alloc_ids_1 | _GEN_1611; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2636 = 7'h4b == rob_alloc_ids_1 | _GEN_1612; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2637 = 7'h4c == rob_alloc_ids_1 | _GEN_1613; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2638 = 7'h4d == rob_alloc_ids_1 | _GEN_1614; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2639 = 7'h4e == rob_alloc_ids_1 | _GEN_1615; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2640 = 7'h4f == rob_alloc_ids_1 | _GEN_1616; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2641 = 7'h50 == rob_alloc_ids_1 | _GEN_1617; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2642 = 7'h51 == rob_alloc_ids_1 | _GEN_1618; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2643 = 7'h52 == rob_alloc_ids_1 | _GEN_1619; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2644 = 7'h53 == rob_alloc_ids_1 | _GEN_1620; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2645 = 7'h54 == rob_alloc_ids_1 | _GEN_1621; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2646 = 7'h55 == rob_alloc_ids_1 | _GEN_1622; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2647 = 7'h56 == rob_alloc_ids_1 | _GEN_1623; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2648 = 7'h57 == rob_alloc_ids_1 | _GEN_1624; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2649 = 7'h58 == rob_alloc_ids_1 | _GEN_1625; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2650 = 7'h59 == rob_alloc_ids_1 | _GEN_1626; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2651 = 7'h5a == rob_alloc_ids_1 | _GEN_1627; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2652 = 7'h5b == rob_alloc_ids_1 | _GEN_1628; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2653 = 7'h5c == rob_alloc_ids_1 | _GEN_1629; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2654 = 7'h5d == rob_alloc_ids_1 | _GEN_1630; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2655 = 7'h5e == rob_alloc_ids_1 | _GEN_1631; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2656 = 7'h5f == rob_alloc_ids_1 | _GEN_1632; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2657 = 7'h60 == rob_alloc_ids_1 | _GEN_1633; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2658 = 7'h61 == rob_alloc_ids_1 | _GEN_1634; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2659 = 7'h62 == rob_alloc_ids_1 | _GEN_1635; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2660 = 7'h63 == rob_alloc_ids_1 | _GEN_1636; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2661 = 7'h64 == rob_alloc_ids_1 | _GEN_1637; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2662 = 7'h65 == rob_alloc_ids_1 | _GEN_1638; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2663 = 7'h66 == rob_alloc_ids_1 | _GEN_1639; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2664 = 7'h67 == rob_alloc_ids_1 | _GEN_1640; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2665 = 7'h68 == rob_alloc_ids_1 | _GEN_1641; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2666 = 7'h69 == rob_alloc_ids_1 | _GEN_1642; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2667 = 7'h6a == rob_alloc_ids_1 | _GEN_1643; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2668 = 7'h6b == rob_alloc_ids_1 | _GEN_1644; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2669 = 7'h6c == rob_alloc_ids_1 | _GEN_1645; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2670 = 7'h6d == rob_alloc_ids_1 | _GEN_1646; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2671 = 7'h6e == rob_alloc_ids_1 | _GEN_1647; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2672 = 7'h6f == rob_alloc_ids_1 | _GEN_1648; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2673 = 7'h70 == rob_alloc_ids_1 | _GEN_1649; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2674 = 7'h71 == rob_alloc_ids_1 | _GEN_1650; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2675 = 7'h72 == rob_alloc_ids_1 | _GEN_1651; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2676 = 7'h73 == rob_alloc_ids_1 | _GEN_1652; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2677 = 7'h74 == rob_alloc_ids_1 | _GEN_1653; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2678 = 7'h75 == rob_alloc_ids_1 | _GEN_1654; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2679 = 7'h76 == rob_alloc_ids_1 | _GEN_1655; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2680 = 7'h77 == rob_alloc_ids_1 | _GEN_1656; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2681 = 7'h78 == rob_alloc_ids_1 | _GEN_1657; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2682 = 7'h79 == rob_alloc_ids_1 | _GEN_1658; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2683 = 7'h7a == rob_alloc_ids_1 | _GEN_1659; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2684 = 7'h7b == rob_alloc_ids_1 | _GEN_1660; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2685 = 7'h7c == rob_alloc_ids_1 | _GEN_1661; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2686 = 7'h7d == rob_alloc_ids_1 | _GEN_1662; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2687 = 7'h7e == rob_alloc_ids_1 | _GEN_1663; // @[TestHarness.scala 181:{36,36}]
  wire  _GEN_2688 = 7'h7f == rob_alloc_ids_1 | _GEN_1664; // @[TestHarness.scala 181:{36,36}]
  wire [3:0] _rob_n_flits_T_35 = igen_1_io_n_flits; // @[TestHarness.scala 182:{36,36}]
  wire [3:0] _GEN_2817 = 7'h0 == rob_alloc_ids_1 ? 4'h0 : _GEN_1793; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2818 = 7'h1 == rob_alloc_ids_1 ? 4'h0 : _GEN_1794; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2819 = 7'h2 == rob_alloc_ids_1 ? 4'h0 : _GEN_1795; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2820 = 7'h3 == rob_alloc_ids_1 ? 4'h0 : _GEN_1796; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2821 = 7'h4 == rob_alloc_ids_1 ? 4'h0 : _GEN_1797; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2822 = 7'h5 == rob_alloc_ids_1 ? 4'h0 : _GEN_1798; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2823 = 7'h6 == rob_alloc_ids_1 ? 4'h0 : _GEN_1799; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2824 = 7'h7 == rob_alloc_ids_1 ? 4'h0 : _GEN_1800; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2825 = 7'h8 == rob_alloc_ids_1 ? 4'h0 : _GEN_1801; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2826 = 7'h9 == rob_alloc_ids_1 ? 4'h0 : _GEN_1802; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2827 = 7'ha == rob_alloc_ids_1 ? 4'h0 : _GEN_1803; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2828 = 7'hb == rob_alloc_ids_1 ? 4'h0 : _GEN_1804; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2829 = 7'hc == rob_alloc_ids_1 ? 4'h0 : _GEN_1805; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2830 = 7'hd == rob_alloc_ids_1 ? 4'h0 : _GEN_1806; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2831 = 7'he == rob_alloc_ids_1 ? 4'h0 : _GEN_1807; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2832 = 7'hf == rob_alloc_ids_1 ? 4'h0 : _GEN_1808; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2833 = 7'h10 == rob_alloc_ids_1 ? 4'h0 : _GEN_1809; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2834 = 7'h11 == rob_alloc_ids_1 ? 4'h0 : _GEN_1810; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2835 = 7'h12 == rob_alloc_ids_1 ? 4'h0 : _GEN_1811; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2836 = 7'h13 == rob_alloc_ids_1 ? 4'h0 : _GEN_1812; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2837 = 7'h14 == rob_alloc_ids_1 ? 4'h0 : _GEN_1813; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2838 = 7'h15 == rob_alloc_ids_1 ? 4'h0 : _GEN_1814; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2839 = 7'h16 == rob_alloc_ids_1 ? 4'h0 : _GEN_1815; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2840 = 7'h17 == rob_alloc_ids_1 ? 4'h0 : _GEN_1816; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2841 = 7'h18 == rob_alloc_ids_1 ? 4'h0 : _GEN_1817; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2842 = 7'h19 == rob_alloc_ids_1 ? 4'h0 : _GEN_1818; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2843 = 7'h1a == rob_alloc_ids_1 ? 4'h0 : _GEN_1819; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2844 = 7'h1b == rob_alloc_ids_1 ? 4'h0 : _GEN_1820; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2845 = 7'h1c == rob_alloc_ids_1 ? 4'h0 : _GEN_1821; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2846 = 7'h1d == rob_alloc_ids_1 ? 4'h0 : _GEN_1822; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2847 = 7'h1e == rob_alloc_ids_1 ? 4'h0 : _GEN_1823; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2848 = 7'h1f == rob_alloc_ids_1 ? 4'h0 : _GEN_1824; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2849 = 7'h20 == rob_alloc_ids_1 ? 4'h0 : _GEN_1825; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2850 = 7'h21 == rob_alloc_ids_1 ? 4'h0 : _GEN_1826; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2851 = 7'h22 == rob_alloc_ids_1 ? 4'h0 : _GEN_1827; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2852 = 7'h23 == rob_alloc_ids_1 ? 4'h0 : _GEN_1828; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2853 = 7'h24 == rob_alloc_ids_1 ? 4'h0 : _GEN_1829; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2854 = 7'h25 == rob_alloc_ids_1 ? 4'h0 : _GEN_1830; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2855 = 7'h26 == rob_alloc_ids_1 ? 4'h0 : _GEN_1831; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2856 = 7'h27 == rob_alloc_ids_1 ? 4'h0 : _GEN_1832; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2857 = 7'h28 == rob_alloc_ids_1 ? 4'h0 : _GEN_1833; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2858 = 7'h29 == rob_alloc_ids_1 ? 4'h0 : _GEN_1834; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2859 = 7'h2a == rob_alloc_ids_1 ? 4'h0 : _GEN_1835; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2860 = 7'h2b == rob_alloc_ids_1 ? 4'h0 : _GEN_1836; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2861 = 7'h2c == rob_alloc_ids_1 ? 4'h0 : _GEN_1837; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2862 = 7'h2d == rob_alloc_ids_1 ? 4'h0 : _GEN_1838; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2863 = 7'h2e == rob_alloc_ids_1 ? 4'h0 : _GEN_1839; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2864 = 7'h2f == rob_alloc_ids_1 ? 4'h0 : _GEN_1840; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2865 = 7'h30 == rob_alloc_ids_1 ? 4'h0 : _GEN_1841; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2866 = 7'h31 == rob_alloc_ids_1 ? 4'h0 : _GEN_1842; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2867 = 7'h32 == rob_alloc_ids_1 ? 4'h0 : _GEN_1843; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2868 = 7'h33 == rob_alloc_ids_1 ? 4'h0 : _GEN_1844; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2869 = 7'h34 == rob_alloc_ids_1 ? 4'h0 : _GEN_1845; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2870 = 7'h35 == rob_alloc_ids_1 ? 4'h0 : _GEN_1846; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2871 = 7'h36 == rob_alloc_ids_1 ? 4'h0 : _GEN_1847; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2872 = 7'h37 == rob_alloc_ids_1 ? 4'h0 : _GEN_1848; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2873 = 7'h38 == rob_alloc_ids_1 ? 4'h0 : _GEN_1849; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2874 = 7'h39 == rob_alloc_ids_1 ? 4'h0 : _GEN_1850; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2875 = 7'h3a == rob_alloc_ids_1 ? 4'h0 : _GEN_1851; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2876 = 7'h3b == rob_alloc_ids_1 ? 4'h0 : _GEN_1852; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2877 = 7'h3c == rob_alloc_ids_1 ? 4'h0 : _GEN_1853; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2878 = 7'h3d == rob_alloc_ids_1 ? 4'h0 : _GEN_1854; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2879 = 7'h3e == rob_alloc_ids_1 ? 4'h0 : _GEN_1855; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2880 = 7'h3f == rob_alloc_ids_1 ? 4'h0 : _GEN_1856; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2881 = 7'h40 == rob_alloc_ids_1 ? 4'h0 : _GEN_1857; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2882 = 7'h41 == rob_alloc_ids_1 ? 4'h0 : _GEN_1858; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2883 = 7'h42 == rob_alloc_ids_1 ? 4'h0 : _GEN_1859; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2884 = 7'h43 == rob_alloc_ids_1 ? 4'h0 : _GEN_1860; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2885 = 7'h44 == rob_alloc_ids_1 ? 4'h0 : _GEN_1861; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2886 = 7'h45 == rob_alloc_ids_1 ? 4'h0 : _GEN_1862; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2887 = 7'h46 == rob_alloc_ids_1 ? 4'h0 : _GEN_1863; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2888 = 7'h47 == rob_alloc_ids_1 ? 4'h0 : _GEN_1864; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2889 = 7'h48 == rob_alloc_ids_1 ? 4'h0 : _GEN_1865; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2890 = 7'h49 == rob_alloc_ids_1 ? 4'h0 : _GEN_1866; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2891 = 7'h4a == rob_alloc_ids_1 ? 4'h0 : _GEN_1867; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2892 = 7'h4b == rob_alloc_ids_1 ? 4'h0 : _GEN_1868; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2893 = 7'h4c == rob_alloc_ids_1 ? 4'h0 : _GEN_1869; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2894 = 7'h4d == rob_alloc_ids_1 ? 4'h0 : _GEN_1870; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2895 = 7'h4e == rob_alloc_ids_1 ? 4'h0 : _GEN_1871; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2896 = 7'h4f == rob_alloc_ids_1 ? 4'h0 : _GEN_1872; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2897 = 7'h50 == rob_alloc_ids_1 ? 4'h0 : _GEN_1873; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2898 = 7'h51 == rob_alloc_ids_1 ? 4'h0 : _GEN_1874; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2899 = 7'h52 == rob_alloc_ids_1 ? 4'h0 : _GEN_1875; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2900 = 7'h53 == rob_alloc_ids_1 ? 4'h0 : _GEN_1876; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2901 = 7'h54 == rob_alloc_ids_1 ? 4'h0 : _GEN_1877; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2902 = 7'h55 == rob_alloc_ids_1 ? 4'h0 : _GEN_1878; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2903 = 7'h56 == rob_alloc_ids_1 ? 4'h0 : _GEN_1879; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2904 = 7'h57 == rob_alloc_ids_1 ? 4'h0 : _GEN_1880; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2905 = 7'h58 == rob_alloc_ids_1 ? 4'h0 : _GEN_1881; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2906 = 7'h59 == rob_alloc_ids_1 ? 4'h0 : _GEN_1882; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2907 = 7'h5a == rob_alloc_ids_1 ? 4'h0 : _GEN_1883; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2908 = 7'h5b == rob_alloc_ids_1 ? 4'h0 : _GEN_1884; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2909 = 7'h5c == rob_alloc_ids_1 ? 4'h0 : _GEN_1885; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2910 = 7'h5d == rob_alloc_ids_1 ? 4'h0 : _GEN_1886; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2911 = 7'h5e == rob_alloc_ids_1 ? 4'h0 : _GEN_1887; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2912 = 7'h5f == rob_alloc_ids_1 ? 4'h0 : _GEN_1888; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2913 = 7'h60 == rob_alloc_ids_1 ? 4'h0 : _GEN_1889; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2914 = 7'h61 == rob_alloc_ids_1 ? 4'h0 : _GEN_1890; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2915 = 7'h62 == rob_alloc_ids_1 ? 4'h0 : _GEN_1891; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2916 = 7'h63 == rob_alloc_ids_1 ? 4'h0 : _GEN_1892; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2917 = 7'h64 == rob_alloc_ids_1 ? 4'h0 : _GEN_1893; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2918 = 7'h65 == rob_alloc_ids_1 ? 4'h0 : _GEN_1894; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2919 = 7'h66 == rob_alloc_ids_1 ? 4'h0 : _GEN_1895; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2920 = 7'h67 == rob_alloc_ids_1 ? 4'h0 : _GEN_1896; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2921 = 7'h68 == rob_alloc_ids_1 ? 4'h0 : _GEN_1897; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2922 = 7'h69 == rob_alloc_ids_1 ? 4'h0 : _GEN_1898; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2923 = 7'h6a == rob_alloc_ids_1 ? 4'h0 : _GEN_1899; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2924 = 7'h6b == rob_alloc_ids_1 ? 4'h0 : _GEN_1900; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2925 = 7'h6c == rob_alloc_ids_1 ? 4'h0 : _GEN_1901; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2926 = 7'h6d == rob_alloc_ids_1 ? 4'h0 : _GEN_1902; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2927 = 7'h6e == rob_alloc_ids_1 ? 4'h0 : _GEN_1903; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2928 = 7'h6f == rob_alloc_ids_1 ? 4'h0 : _GEN_1904; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2929 = 7'h70 == rob_alloc_ids_1 ? 4'h0 : _GEN_1905; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2930 = 7'h71 == rob_alloc_ids_1 ? 4'h0 : _GEN_1906; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2931 = 7'h72 == rob_alloc_ids_1 ? 4'h0 : _GEN_1907; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2932 = 7'h73 == rob_alloc_ids_1 ? 4'h0 : _GEN_1908; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2933 = 7'h74 == rob_alloc_ids_1 ? 4'h0 : _GEN_1909; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2934 = 7'h75 == rob_alloc_ids_1 ? 4'h0 : _GEN_1910; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2935 = 7'h76 == rob_alloc_ids_1 ? 4'h0 : _GEN_1911; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2936 = 7'h77 == rob_alloc_ids_1 ? 4'h0 : _GEN_1912; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2937 = 7'h78 == rob_alloc_ids_1 ? 4'h0 : _GEN_1913; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2938 = 7'h79 == rob_alloc_ids_1 ? 4'h0 : _GEN_1914; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2939 = 7'h7a == rob_alloc_ids_1 ? 4'h0 : _GEN_1915; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2940 = 7'h7b == rob_alloc_ids_1 ? 4'h0 : _GEN_1916; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2941 = 7'h7c == rob_alloc_ids_1 ? 4'h0 : _GEN_1917; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2942 = 7'h7d == rob_alloc_ids_1 ? 4'h0 : _GEN_1918; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2943 = 7'h7e == rob_alloc_ids_1 ? 4'h0 : _GEN_1919; // @[TestHarness.scala 183:{36,36}]
  wire [3:0] _GEN_2944 = 7'h7f == rob_alloc_ids_1 ? 4'h0 : _GEN_1920; // @[TestHarness.scala 183:{36,36}]
  wire [15:0] _GEN_3329 = igen_1_io_fire ? _GEN_2305 : _GEN_1281; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3330 = igen_1_io_fire ? _GEN_2306 : _GEN_1282; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3331 = igen_1_io_fire ? _GEN_2307 : _GEN_1283; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3332 = igen_1_io_fire ? _GEN_2308 : _GEN_1284; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3333 = igen_1_io_fire ? _GEN_2309 : _GEN_1285; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3334 = igen_1_io_fire ? _GEN_2310 : _GEN_1286; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3335 = igen_1_io_fire ? _GEN_2311 : _GEN_1287; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3336 = igen_1_io_fire ? _GEN_2312 : _GEN_1288; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3337 = igen_1_io_fire ? _GEN_2313 : _GEN_1289; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3338 = igen_1_io_fire ? _GEN_2314 : _GEN_1290; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3339 = igen_1_io_fire ? _GEN_2315 : _GEN_1291; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3340 = igen_1_io_fire ? _GEN_2316 : _GEN_1292; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3341 = igen_1_io_fire ? _GEN_2317 : _GEN_1293; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3342 = igen_1_io_fire ? _GEN_2318 : _GEN_1294; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3343 = igen_1_io_fire ? _GEN_2319 : _GEN_1295; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3344 = igen_1_io_fire ? _GEN_2320 : _GEN_1296; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3345 = igen_1_io_fire ? _GEN_2321 : _GEN_1297; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3346 = igen_1_io_fire ? _GEN_2322 : _GEN_1298; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3347 = igen_1_io_fire ? _GEN_2323 : _GEN_1299; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3348 = igen_1_io_fire ? _GEN_2324 : _GEN_1300; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3349 = igen_1_io_fire ? _GEN_2325 : _GEN_1301; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3350 = igen_1_io_fire ? _GEN_2326 : _GEN_1302; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3351 = igen_1_io_fire ? _GEN_2327 : _GEN_1303; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3352 = igen_1_io_fire ? _GEN_2328 : _GEN_1304; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3353 = igen_1_io_fire ? _GEN_2329 : _GEN_1305; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3354 = igen_1_io_fire ? _GEN_2330 : _GEN_1306; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3355 = igen_1_io_fire ? _GEN_2331 : _GEN_1307; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3356 = igen_1_io_fire ? _GEN_2332 : _GEN_1308; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3357 = igen_1_io_fire ? _GEN_2333 : _GEN_1309; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3358 = igen_1_io_fire ? _GEN_2334 : _GEN_1310; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3359 = igen_1_io_fire ? _GEN_2335 : _GEN_1311; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3360 = igen_1_io_fire ? _GEN_2336 : _GEN_1312; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3361 = igen_1_io_fire ? _GEN_2337 : _GEN_1313; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3362 = igen_1_io_fire ? _GEN_2338 : _GEN_1314; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3363 = igen_1_io_fire ? _GEN_2339 : _GEN_1315; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3364 = igen_1_io_fire ? _GEN_2340 : _GEN_1316; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3365 = igen_1_io_fire ? _GEN_2341 : _GEN_1317; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3366 = igen_1_io_fire ? _GEN_2342 : _GEN_1318; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3367 = igen_1_io_fire ? _GEN_2343 : _GEN_1319; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3368 = igen_1_io_fire ? _GEN_2344 : _GEN_1320; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3369 = igen_1_io_fire ? _GEN_2345 : _GEN_1321; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3370 = igen_1_io_fire ? _GEN_2346 : _GEN_1322; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3371 = igen_1_io_fire ? _GEN_2347 : _GEN_1323; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3372 = igen_1_io_fire ? _GEN_2348 : _GEN_1324; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3373 = igen_1_io_fire ? _GEN_2349 : _GEN_1325; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3374 = igen_1_io_fire ? _GEN_2350 : _GEN_1326; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3375 = igen_1_io_fire ? _GEN_2351 : _GEN_1327; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3376 = igen_1_io_fire ? _GEN_2352 : _GEN_1328; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3377 = igen_1_io_fire ? _GEN_2353 : _GEN_1329; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3378 = igen_1_io_fire ? _GEN_2354 : _GEN_1330; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3379 = igen_1_io_fire ? _GEN_2355 : _GEN_1331; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3380 = igen_1_io_fire ? _GEN_2356 : _GEN_1332; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3381 = igen_1_io_fire ? _GEN_2357 : _GEN_1333; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3382 = igen_1_io_fire ? _GEN_2358 : _GEN_1334; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3383 = igen_1_io_fire ? _GEN_2359 : _GEN_1335; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3384 = igen_1_io_fire ? _GEN_2360 : _GEN_1336; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3385 = igen_1_io_fire ? _GEN_2361 : _GEN_1337; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3386 = igen_1_io_fire ? _GEN_2362 : _GEN_1338; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3387 = igen_1_io_fire ? _GEN_2363 : _GEN_1339; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3388 = igen_1_io_fire ? _GEN_2364 : _GEN_1340; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3389 = igen_1_io_fire ? _GEN_2365 : _GEN_1341; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3390 = igen_1_io_fire ? _GEN_2366 : _GEN_1342; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3391 = igen_1_io_fire ? _GEN_2367 : _GEN_1343; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3392 = igen_1_io_fire ? _GEN_2368 : _GEN_1344; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3393 = igen_1_io_fire ? _GEN_2369 : _GEN_1345; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3394 = igen_1_io_fire ? _GEN_2370 : _GEN_1346; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3395 = igen_1_io_fire ? _GEN_2371 : _GEN_1347; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3396 = igen_1_io_fire ? _GEN_2372 : _GEN_1348; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3397 = igen_1_io_fire ? _GEN_2373 : _GEN_1349; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3398 = igen_1_io_fire ? _GEN_2374 : _GEN_1350; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3399 = igen_1_io_fire ? _GEN_2375 : _GEN_1351; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3400 = igen_1_io_fire ? _GEN_2376 : _GEN_1352; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3401 = igen_1_io_fire ? _GEN_2377 : _GEN_1353; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3402 = igen_1_io_fire ? _GEN_2378 : _GEN_1354; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3403 = igen_1_io_fire ? _GEN_2379 : _GEN_1355; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3404 = igen_1_io_fire ? _GEN_2380 : _GEN_1356; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3405 = igen_1_io_fire ? _GEN_2381 : _GEN_1357; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3406 = igen_1_io_fire ? _GEN_2382 : _GEN_1358; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3407 = igen_1_io_fire ? _GEN_2383 : _GEN_1359; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3408 = igen_1_io_fire ? _GEN_2384 : _GEN_1360; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3409 = igen_1_io_fire ? _GEN_2385 : _GEN_1361; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3410 = igen_1_io_fire ? _GEN_2386 : _GEN_1362; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3411 = igen_1_io_fire ? _GEN_2387 : _GEN_1363; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3412 = igen_1_io_fire ? _GEN_2388 : _GEN_1364; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3413 = igen_1_io_fire ? _GEN_2389 : _GEN_1365; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3414 = igen_1_io_fire ? _GEN_2390 : _GEN_1366; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3415 = igen_1_io_fire ? _GEN_2391 : _GEN_1367; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3416 = igen_1_io_fire ? _GEN_2392 : _GEN_1368; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3417 = igen_1_io_fire ? _GEN_2393 : _GEN_1369; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3418 = igen_1_io_fire ? _GEN_2394 : _GEN_1370; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3419 = igen_1_io_fire ? _GEN_2395 : _GEN_1371; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3420 = igen_1_io_fire ? _GEN_2396 : _GEN_1372; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3421 = igen_1_io_fire ? _GEN_2397 : _GEN_1373; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3422 = igen_1_io_fire ? _GEN_2398 : _GEN_1374; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3423 = igen_1_io_fire ? _GEN_2399 : _GEN_1375; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3424 = igen_1_io_fire ? _GEN_2400 : _GEN_1376; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3425 = igen_1_io_fire ? _GEN_2401 : _GEN_1377; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3426 = igen_1_io_fire ? _GEN_2402 : _GEN_1378; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3427 = igen_1_io_fire ? _GEN_2403 : _GEN_1379; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3428 = igen_1_io_fire ? _GEN_2404 : _GEN_1380; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3429 = igen_1_io_fire ? _GEN_2405 : _GEN_1381; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3430 = igen_1_io_fire ? _GEN_2406 : _GEN_1382; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3431 = igen_1_io_fire ? _GEN_2407 : _GEN_1383; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3432 = igen_1_io_fire ? _GEN_2408 : _GEN_1384; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3433 = igen_1_io_fire ? _GEN_2409 : _GEN_1385; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3434 = igen_1_io_fire ? _GEN_2410 : _GEN_1386; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3435 = igen_1_io_fire ? _GEN_2411 : _GEN_1387; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3436 = igen_1_io_fire ? _GEN_2412 : _GEN_1388; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3437 = igen_1_io_fire ? _GEN_2413 : _GEN_1389; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3438 = igen_1_io_fire ? _GEN_2414 : _GEN_1390; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3439 = igen_1_io_fire ? _GEN_2415 : _GEN_1391; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3440 = igen_1_io_fire ? _GEN_2416 : _GEN_1392; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3441 = igen_1_io_fire ? _GEN_2417 : _GEN_1393; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3442 = igen_1_io_fire ? _GEN_2418 : _GEN_1394; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3443 = igen_1_io_fire ? _GEN_2419 : _GEN_1395; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3444 = igen_1_io_fire ? _GEN_2420 : _GEN_1396; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3445 = igen_1_io_fire ? _GEN_2421 : _GEN_1397; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3446 = igen_1_io_fire ? _GEN_2422 : _GEN_1398; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3447 = igen_1_io_fire ? _GEN_2423 : _GEN_1399; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3448 = igen_1_io_fire ? _GEN_2424 : _GEN_1400; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3449 = igen_1_io_fire ? _GEN_2425 : _GEN_1401; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3450 = igen_1_io_fire ? _GEN_2426 : _GEN_1402; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3451 = igen_1_io_fire ? _GEN_2427 : _GEN_1403; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3452 = igen_1_io_fire ? _GEN_2428 : _GEN_1404; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3453 = igen_1_io_fire ? _GEN_2429 : _GEN_1405; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3454 = igen_1_io_fire ? _GEN_2430 : _GEN_1406; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3455 = igen_1_io_fire ? _GEN_2431 : _GEN_1407; // @[TestHarness.scala 178:25]
  wire [15:0] _GEN_3456 = igen_1_io_fire ? _GEN_2432 : _GEN_1408; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3841 = igen_1_io_fire ? _GEN_2817 : _GEN_1793; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3842 = igen_1_io_fire ? _GEN_2818 : _GEN_1794; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3843 = igen_1_io_fire ? _GEN_2819 : _GEN_1795; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3844 = igen_1_io_fire ? _GEN_2820 : _GEN_1796; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3845 = igen_1_io_fire ? _GEN_2821 : _GEN_1797; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3846 = igen_1_io_fire ? _GEN_2822 : _GEN_1798; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3847 = igen_1_io_fire ? _GEN_2823 : _GEN_1799; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3848 = igen_1_io_fire ? _GEN_2824 : _GEN_1800; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3849 = igen_1_io_fire ? _GEN_2825 : _GEN_1801; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3850 = igen_1_io_fire ? _GEN_2826 : _GEN_1802; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3851 = igen_1_io_fire ? _GEN_2827 : _GEN_1803; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3852 = igen_1_io_fire ? _GEN_2828 : _GEN_1804; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3853 = igen_1_io_fire ? _GEN_2829 : _GEN_1805; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3854 = igen_1_io_fire ? _GEN_2830 : _GEN_1806; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3855 = igen_1_io_fire ? _GEN_2831 : _GEN_1807; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3856 = igen_1_io_fire ? _GEN_2832 : _GEN_1808; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3857 = igen_1_io_fire ? _GEN_2833 : _GEN_1809; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3858 = igen_1_io_fire ? _GEN_2834 : _GEN_1810; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3859 = igen_1_io_fire ? _GEN_2835 : _GEN_1811; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3860 = igen_1_io_fire ? _GEN_2836 : _GEN_1812; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3861 = igen_1_io_fire ? _GEN_2837 : _GEN_1813; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3862 = igen_1_io_fire ? _GEN_2838 : _GEN_1814; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3863 = igen_1_io_fire ? _GEN_2839 : _GEN_1815; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3864 = igen_1_io_fire ? _GEN_2840 : _GEN_1816; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3865 = igen_1_io_fire ? _GEN_2841 : _GEN_1817; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3866 = igen_1_io_fire ? _GEN_2842 : _GEN_1818; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3867 = igen_1_io_fire ? _GEN_2843 : _GEN_1819; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3868 = igen_1_io_fire ? _GEN_2844 : _GEN_1820; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3869 = igen_1_io_fire ? _GEN_2845 : _GEN_1821; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3870 = igen_1_io_fire ? _GEN_2846 : _GEN_1822; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3871 = igen_1_io_fire ? _GEN_2847 : _GEN_1823; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3872 = igen_1_io_fire ? _GEN_2848 : _GEN_1824; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3873 = igen_1_io_fire ? _GEN_2849 : _GEN_1825; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3874 = igen_1_io_fire ? _GEN_2850 : _GEN_1826; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3875 = igen_1_io_fire ? _GEN_2851 : _GEN_1827; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3876 = igen_1_io_fire ? _GEN_2852 : _GEN_1828; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3877 = igen_1_io_fire ? _GEN_2853 : _GEN_1829; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3878 = igen_1_io_fire ? _GEN_2854 : _GEN_1830; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3879 = igen_1_io_fire ? _GEN_2855 : _GEN_1831; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3880 = igen_1_io_fire ? _GEN_2856 : _GEN_1832; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3881 = igen_1_io_fire ? _GEN_2857 : _GEN_1833; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3882 = igen_1_io_fire ? _GEN_2858 : _GEN_1834; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3883 = igen_1_io_fire ? _GEN_2859 : _GEN_1835; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3884 = igen_1_io_fire ? _GEN_2860 : _GEN_1836; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3885 = igen_1_io_fire ? _GEN_2861 : _GEN_1837; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3886 = igen_1_io_fire ? _GEN_2862 : _GEN_1838; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3887 = igen_1_io_fire ? _GEN_2863 : _GEN_1839; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3888 = igen_1_io_fire ? _GEN_2864 : _GEN_1840; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3889 = igen_1_io_fire ? _GEN_2865 : _GEN_1841; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3890 = igen_1_io_fire ? _GEN_2866 : _GEN_1842; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3891 = igen_1_io_fire ? _GEN_2867 : _GEN_1843; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3892 = igen_1_io_fire ? _GEN_2868 : _GEN_1844; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3893 = igen_1_io_fire ? _GEN_2869 : _GEN_1845; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3894 = igen_1_io_fire ? _GEN_2870 : _GEN_1846; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3895 = igen_1_io_fire ? _GEN_2871 : _GEN_1847; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3896 = igen_1_io_fire ? _GEN_2872 : _GEN_1848; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3897 = igen_1_io_fire ? _GEN_2873 : _GEN_1849; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3898 = igen_1_io_fire ? _GEN_2874 : _GEN_1850; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3899 = igen_1_io_fire ? _GEN_2875 : _GEN_1851; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3900 = igen_1_io_fire ? _GEN_2876 : _GEN_1852; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3901 = igen_1_io_fire ? _GEN_2877 : _GEN_1853; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3902 = igen_1_io_fire ? _GEN_2878 : _GEN_1854; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3903 = igen_1_io_fire ? _GEN_2879 : _GEN_1855; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3904 = igen_1_io_fire ? _GEN_2880 : _GEN_1856; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3905 = igen_1_io_fire ? _GEN_2881 : _GEN_1857; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3906 = igen_1_io_fire ? _GEN_2882 : _GEN_1858; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3907 = igen_1_io_fire ? _GEN_2883 : _GEN_1859; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3908 = igen_1_io_fire ? _GEN_2884 : _GEN_1860; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3909 = igen_1_io_fire ? _GEN_2885 : _GEN_1861; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3910 = igen_1_io_fire ? _GEN_2886 : _GEN_1862; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3911 = igen_1_io_fire ? _GEN_2887 : _GEN_1863; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3912 = igen_1_io_fire ? _GEN_2888 : _GEN_1864; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3913 = igen_1_io_fire ? _GEN_2889 : _GEN_1865; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3914 = igen_1_io_fire ? _GEN_2890 : _GEN_1866; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3915 = igen_1_io_fire ? _GEN_2891 : _GEN_1867; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3916 = igen_1_io_fire ? _GEN_2892 : _GEN_1868; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3917 = igen_1_io_fire ? _GEN_2893 : _GEN_1869; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3918 = igen_1_io_fire ? _GEN_2894 : _GEN_1870; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3919 = igen_1_io_fire ? _GEN_2895 : _GEN_1871; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3920 = igen_1_io_fire ? _GEN_2896 : _GEN_1872; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3921 = igen_1_io_fire ? _GEN_2897 : _GEN_1873; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3922 = igen_1_io_fire ? _GEN_2898 : _GEN_1874; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3923 = igen_1_io_fire ? _GEN_2899 : _GEN_1875; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3924 = igen_1_io_fire ? _GEN_2900 : _GEN_1876; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3925 = igen_1_io_fire ? _GEN_2901 : _GEN_1877; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3926 = igen_1_io_fire ? _GEN_2902 : _GEN_1878; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3927 = igen_1_io_fire ? _GEN_2903 : _GEN_1879; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3928 = igen_1_io_fire ? _GEN_2904 : _GEN_1880; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3929 = igen_1_io_fire ? _GEN_2905 : _GEN_1881; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3930 = igen_1_io_fire ? _GEN_2906 : _GEN_1882; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3931 = igen_1_io_fire ? _GEN_2907 : _GEN_1883; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3932 = igen_1_io_fire ? _GEN_2908 : _GEN_1884; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3933 = igen_1_io_fire ? _GEN_2909 : _GEN_1885; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3934 = igen_1_io_fire ? _GEN_2910 : _GEN_1886; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3935 = igen_1_io_fire ? _GEN_2911 : _GEN_1887; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3936 = igen_1_io_fire ? _GEN_2912 : _GEN_1888; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3937 = igen_1_io_fire ? _GEN_2913 : _GEN_1889; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3938 = igen_1_io_fire ? _GEN_2914 : _GEN_1890; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3939 = igen_1_io_fire ? _GEN_2915 : _GEN_1891; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3940 = igen_1_io_fire ? _GEN_2916 : _GEN_1892; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3941 = igen_1_io_fire ? _GEN_2917 : _GEN_1893; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3942 = igen_1_io_fire ? _GEN_2918 : _GEN_1894; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3943 = igen_1_io_fire ? _GEN_2919 : _GEN_1895; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3944 = igen_1_io_fire ? _GEN_2920 : _GEN_1896; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3945 = igen_1_io_fire ? _GEN_2921 : _GEN_1897; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3946 = igen_1_io_fire ? _GEN_2922 : _GEN_1898; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3947 = igen_1_io_fire ? _GEN_2923 : _GEN_1899; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3948 = igen_1_io_fire ? _GEN_2924 : _GEN_1900; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3949 = igen_1_io_fire ? _GEN_2925 : _GEN_1901; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3950 = igen_1_io_fire ? _GEN_2926 : _GEN_1902; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3951 = igen_1_io_fire ? _GEN_2927 : _GEN_1903; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3952 = igen_1_io_fire ? _GEN_2928 : _GEN_1904; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3953 = igen_1_io_fire ? _GEN_2929 : _GEN_1905; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3954 = igen_1_io_fire ? _GEN_2930 : _GEN_1906; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3955 = igen_1_io_fire ? _GEN_2931 : _GEN_1907; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3956 = igen_1_io_fire ? _GEN_2932 : _GEN_1908; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3957 = igen_1_io_fire ? _GEN_2933 : _GEN_1909; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3958 = igen_1_io_fire ? _GEN_2934 : _GEN_1910; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3959 = igen_1_io_fire ? _GEN_2935 : _GEN_1911; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3960 = igen_1_io_fire ? _GEN_2936 : _GEN_1912; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3961 = igen_1_io_fire ? _GEN_2937 : _GEN_1913; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3962 = igen_1_io_fire ? _GEN_2938 : _GEN_1914; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3963 = igen_1_io_fire ? _GEN_2939 : _GEN_1915; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3964 = igen_1_io_fire ? _GEN_2940 : _GEN_1916; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3965 = igen_1_io_fire ? _GEN_2941 : _GEN_1917; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3966 = igen_1_io_fire ? _GEN_2942 : _GEN_1918; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3967 = igen_1_io_fire ? _GEN_2943 : _GEN_1919; // @[TestHarness.scala 178:25]
  wire [3:0] _GEN_3968 = igen_1_io_fire ? _GEN_2944 : _GEN_1920; // @[TestHarness.scala 178:25]
  wire  enable_print_latency = plusarg_reader_out; // @[TestHarness.scala 190:81]
  wire [31:0] out_payload_tsc = io_from_noc_0_flit_bits_payload[63:32]; // @[TestHarness.scala 194:51]
  reg  packet_valid; // @[TestHarness.scala 196:31]
  reg [6:0] packet_rob_idx; // @[TestHarness.scala 197:29]
  wire [127:0] _T_42 = rob_valids >> out_payload_rob_idx; // @[TestHarness.scala 201:24]
  wire [31:0] _GEN_4098 = 7'h1 == out_payload_rob_idx[6:0] ? rob_payload_1_tsc : rob_payload_0_tsc; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4099 = 7'h2 == out_payload_rob_idx[6:0] ? rob_payload_2_tsc : _GEN_4098; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4100 = 7'h3 == out_payload_rob_idx[6:0] ? rob_payload_3_tsc : _GEN_4099; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4101 = 7'h4 == out_payload_rob_idx[6:0] ? rob_payload_4_tsc : _GEN_4100; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4102 = 7'h5 == out_payload_rob_idx[6:0] ? rob_payload_5_tsc : _GEN_4101; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4103 = 7'h6 == out_payload_rob_idx[6:0] ? rob_payload_6_tsc : _GEN_4102; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4104 = 7'h7 == out_payload_rob_idx[6:0] ? rob_payload_7_tsc : _GEN_4103; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4105 = 7'h8 == out_payload_rob_idx[6:0] ? rob_payload_8_tsc : _GEN_4104; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4106 = 7'h9 == out_payload_rob_idx[6:0] ? rob_payload_9_tsc : _GEN_4105; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4107 = 7'ha == out_payload_rob_idx[6:0] ? rob_payload_10_tsc : _GEN_4106; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4108 = 7'hb == out_payload_rob_idx[6:0] ? rob_payload_11_tsc : _GEN_4107; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4109 = 7'hc == out_payload_rob_idx[6:0] ? rob_payload_12_tsc : _GEN_4108; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4110 = 7'hd == out_payload_rob_idx[6:0] ? rob_payload_13_tsc : _GEN_4109; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4111 = 7'he == out_payload_rob_idx[6:0] ? rob_payload_14_tsc : _GEN_4110; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4112 = 7'hf == out_payload_rob_idx[6:0] ? rob_payload_15_tsc : _GEN_4111; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4113 = 7'h10 == out_payload_rob_idx[6:0] ? rob_payload_16_tsc : _GEN_4112; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4114 = 7'h11 == out_payload_rob_idx[6:0] ? rob_payload_17_tsc : _GEN_4113; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4115 = 7'h12 == out_payload_rob_idx[6:0] ? rob_payload_18_tsc : _GEN_4114; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4116 = 7'h13 == out_payload_rob_idx[6:0] ? rob_payload_19_tsc : _GEN_4115; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4117 = 7'h14 == out_payload_rob_idx[6:0] ? rob_payload_20_tsc : _GEN_4116; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4118 = 7'h15 == out_payload_rob_idx[6:0] ? rob_payload_21_tsc : _GEN_4117; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4119 = 7'h16 == out_payload_rob_idx[6:0] ? rob_payload_22_tsc : _GEN_4118; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4120 = 7'h17 == out_payload_rob_idx[6:0] ? rob_payload_23_tsc : _GEN_4119; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4121 = 7'h18 == out_payload_rob_idx[6:0] ? rob_payload_24_tsc : _GEN_4120; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4122 = 7'h19 == out_payload_rob_idx[6:0] ? rob_payload_25_tsc : _GEN_4121; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4123 = 7'h1a == out_payload_rob_idx[6:0] ? rob_payload_26_tsc : _GEN_4122; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4124 = 7'h1b == out_payload_rob_idx[6:0] ? rob_payload_27_tsc : _GEN_4123; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4125 = 7'h1c == out_payload_rob_idx[6:0] ? rob_payload_28_tsc : _GEN_4124; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4126 = 7'h1d == out_payload_rob_idx[6:0] ? rob_payload_29_tsc : _GEN_4125; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4127 = 7'h1e == out_payload_rob_idx[6:0] ? rob_payload_30_tsc : _GEN_4126; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4128 = 7'h1f == out_payload_rob_idx[6:0] ? rob_payload_31_tsc : _GEN_4127; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4129 = 7'h20 == out_payload_rob_idx[6:0] ? rob_payload_32_tsc : _GEN_4128; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4130 = 7'h21 == out_payload_rob_idx[6:0] ? rob_payload_33_tsc : _GEN_4129; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4131 = 7'h22 == out_payload_rob_idx[6:0] ? rob_payload_34_tsc : _GEN_4130; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4132 = 7'h23 == out_payload_rob_idx[6:0] ? rob_payload_35_tsc : _GEN_4131; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4133 = 7'h24 == out_payload_rob_idx[6:0] ? rob_payload_36_tsc : _GEN_4132; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4134 = 7'h25 == out_payload_rob_idx[6:0] ? rob_payload_37_tsc : _GEN_4133; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4135 = 7'h26 == out_payload_rob_idx[6:0] ? rob_payload_38_tsc : _GEN_4134; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4136 = 7'h27 == out_payload_rob_idx[6:0] ? rob_payload_39_tsc : _GEN_4135; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4137 = 7'h28 == out_payload_rob_idx[6:0] ? rob_payload_40_tsc : _GEN_4136; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4138 = 7'h29 == out_payload_rob_idx[6:0] ? rob_payload_41_tsc : _GEN_4137; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4139 = 7'h2a == out_payload_rob_idx[6:0] ? rob_payload_42_tsc : _GEN_4138; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4140 = 7'h2b == out_payload_rob_idx[6:0] ? rob_payload_43_tsc : _GEN_4139; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4141 = 7'h2c == out_payload_rob_idx[6:0] ? rob_payload_44_tsc : _GEN_4140; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4142 = 7'h2d == out_payload_rob_idx[6:0] ? rob_payload_45_tsc : _GEN_4141; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4143 = 7'h2e == out_payload_rob_idx[6:0] ? rob_payload_46_tsc : _GEN_4142; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4144 = 7'h2f == out_payload_rob_idx[6:0] ? rob_payload_47_tsc : _GEN_4143; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4145 = 7'h30 == out_payload_rob_idx[6:0] ? rob_payload_48_tsc : _GEN_4144; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4146 = 7'h31 == out_payload_rob_idx[6:0] ? rob_payload_49_tsc : _GEN_4145; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4147 = 7'h32 == out_payload_rob_idx[6:0] ? rob_payload_50_tsc : _GEN_4146; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4148 = 7'h33 == out_payload_rob_idx[6:0] ? rob_payload_51_tsc : _GEN_4147; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4149 = 7'h34 == out_payload_rob_idx[6:0] ? rob_payload_52_tsc : _GEN_4148; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4150 = 7'h35 == out_payload_rob_idx[6:0] ? rob_payload_53_tsc : _GEN_4149; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4151 = 7'h36 == out_payload_rob_idx[6:0] ? rob_payload_54_tsc : _GEN_4150; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4152 = 7'h37 == out_payload_rob_idx[6:0] ? rob_payload_55_tsc : _GEN_4151; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4153 = 7'h38 == out_payload_rob_idx[6:0] ? rob_payload_56_tsc : _GEN_4152; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4154 = 7'h39 == out_payload_rob_idx[6:0] ? rob_payload_57_tsc : _GEN_4153; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4155 = 7'h3a == out_payload_rob_idx[6:0] ? rob_payload_58_tsc : _GEN_4154; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4156 = 7'h3b == out_payload_rob_idx[6:0] ? rob_payload_59_tsc : _GEN_4155; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4157 = 7'h3c == out_payload_rob_idx[6:0] ? rob_payload_60_tsc : _GEN_4156; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4158 = 7'h3d == out_payload_rob_idx[6:0] ? rob_payload_61_tsc : _GEN_4157; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4159 = 7'h3e == out_payload_rob_idx[6:0] ? rob_payload_62_tsc : _GEN_4158; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4160 = 7'h3f == out_payload_rob_idx[6:0] ? rob_payload_63_tsc : _GEN_4159; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4161 = 7'h40 == out_payload_rob_idx[6:0] ? rob_payload_64_tsc : _GEN_4160; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4162 = 7'h41 == out_payload_rob_idx[6:0] ? rob_payload_65_tsc : _GEN_4161; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4163 = 7'h42 == out_payload_rob_idx[6:0] ? rob_payload_66_tsc : _GEN_4162; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4164 = 7'h43 == out_payload_rob_idx[6:0] ? rob_payload_67_tsc : _GEN_4163; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4165 = 7'h44 == out_payload_rob_idx[6:0] ? rob_payload_68_tsc : _GEN_4164; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4166 = 7'h45 == out_payload_rob_idx[6:0] ? rob_payload_69_tsc : _GEN_4165; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4167 = 7'h46 == out_payload_rob_idx[6:0] ? rob_payload_70_tsc : _GEN_4166; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4168 = 7'h47 == out_payload_rob_idx[6:0] ? rob_payload_71_tsc : _GEN_4167; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4169 = 7'h48 == out_payload_rob_idx[6:0] ? rob_payload_72_tsc : _GEN_4168; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4170 = 7'h49 == out_payload_rob_idx[6:0] ? rob_payload_73_tsc : _GEN_4169; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4171 = 7'h4a == out_payload_rob_idx[6:0] ? rob_payload_74_tsc : _GEN_4170; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4172 = 7'h4b == out_payload_rob_idx[6:0] ? rob_payload_75_tsc : _GEN_4171; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4173 = 7'h4c == out_payload_rob_idx[6:0] ? rob_payload_76_tsc : _GEN_4172; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4174 = 7'h4d == out_payload_rob_idx[6:0] ? rob_payload_77_tsc : _GEN_4173; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4175 = 7'h4e == out_payload_rob_idx[6:0] ? rob_payload_78_tsc : _GEN_4174; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4176 = 7'h4f == out_payload_rob_idx[6:0] ? rob_payload_79_tsc : _GEN_4175; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4177 = 7'h50 == out_payload_rob_idx[6:0] ? rob_payload_80_tsc : _GEN_4176; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4178 = 7'h51 == out_payload_rob_idx[6:0] ? rob_payload_81_tsc : _GEN_4177; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4179 = 7'h52 == out_payload_rob_idx[6:0] ? rob_payload_82_tsc : _GEN_4178; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4180 = 7'h53 == out_payload_rob_idx[6:0] ? rob_payload_83_tsc : _GEN_4179; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4181 = 7'h54 == out_payload_rob_idx[6:0] ? rob_payload_84_tsc : _GEN_4180; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4182 = 7'h55 == out_payload_rob_idx[6:0] ? rob_payload_85_tsc : _GEN_4181; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4183 = 7'h56 == out_payload_rob_idx[6:0] ? rob_payload_86_tsc : _GEN_4182; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4184 = 7'h57 == out_payload_rob_idx[6:0] ? rob_payload_87_tsc : _GEN_4183; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4185 = 7'h58 == out_payload_rob_idx[6:0] ? rob_payload_88_tsc : _GEN_4184; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4186 = 7'h59 == out_payload_rob_idx[6:0] ? rob_payload_89_tsc : _GEN_4185; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4187 = 7'h5a == out_payload_rob_idx[6:0] ? rob_payload_90_tsc : _GEN_4186; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4188 = 7'h5b == out_payload_rob_idx[6:0] ? rob_payload_91_tsc : _GEN_4187; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4189 = 7'h5c == out_payload_rob_idx[6:0] ? rob_payload_92_tsc : _GEN_4188; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4190 = 7'h5d == out_payload_rob_idx[6:0] ? rob_payload_93_tsc : _GEN_4189; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4191 = 7'h5e == out_payload_rob_idx[6:0] ? rob_payload_94_tsc : _GEN_4190; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4192 = 7'h5f == out_payload_rob_idx[6:0] ? rob_payload_95_tsc : _GEN_4191; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4193 = 7'h60 == out_payload_rob_idx[6:0] ? rob_payload_96_tsc : _GEN_4192; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4194 = 7'h61 == out_payload_rob_idx[6:0] ? rob_payload_97_tsc : _GEN_4193; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4195 = 7'h62 == out_payload_rob_idx[6:0] ? rob_payload_98_tsc : _GEN_4194; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4196 = 7'h63 == out_payload_rob_idx[6:0] ? rob_payload_99_tsc : _GEN_4195; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4197 = 7'h64 == out_payload_rob_idx[6:0] ? rob_payload_100_tsc : _GEN_4196; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4198 = 7'h65 == out_payload_rob_idx[6:0] ? rob_payload_101_tsc : _GEN_4197; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4199 = 7'h66 == out_payload_rob_idx[6:0] ? rob_payload_102_tsc : _GEN_4198; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4200 = 7'h67 == out_payload_rob_idx[6:0] ? rob_payload_103_tsc : _GEN_4199; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4201 = 7'h68 == out_payload_rob_idx[6:0] ? rob_payload_104_tsc : _GEN_4200; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4202 = 7'h69 == out_payload_rob_idx[6:0] ? rob_payload_105_tsc : _GEN_4201; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4203 = 7'h6a == out_payload_rob_idx[6:0] ? rob_payload_106_tsc : _GEN_4202; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4204 = 7'h6b == out_payload_rob_idx[6:0] ? rob_payload_107_tsc : _GEN_4203; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4205 = 7'h6c == out_payload_rob_idx[6:0] ? rob_payload_108_tsc : _GEN_4204; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4206 = 7'h6d == out_payload_rob_idx[6:0] ? rob_payload_109_tsc : _GEN_4205; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4207 = 7'h6e == out_payload_rob_idx[6:0] ? rob_payload_110_tsc : _GEN_4206; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4208 = 7'h6f == out_payload_rob_idx[6:0] ? rob_payload_111_tsc : _GEN_4207; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4209 = 7'h70 == out_payload_rob_idx[6:0] ? rob_payload_112_tsc : _GEN_4208; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4210 = 7'h71 == out_payload_rob_idx[6:0] ? rob_payload_113_tsc : _GEN_4209; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4211 = 7'h72 == out_payload_rob_idx[6:0] ? rob_payload_114_tsc : _GEN_4210; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4212 = 7'h73 == out_payload_rob_idx[6:0] ? rob_payload_115_tsc : _GEN_4211; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4213 = 7'h74 == out_payload_rob_idx[6:0] ? rob_payload_116_tsc : _GEN_4212; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4214 = 7'h75 == out_payload_rob_idx[6:0] ? rob_payload_117_tsc : _GEN_4213; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4215 = 7'h76 == out_payload_rob_idx[6:0] ? rob_payload_118_tsc : _GEN_4214; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4216 = 7'h77 == out_payload_rob_idx[6:0] ? rob_payload_119_tsc : _GEN_4215; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4217 = 7'h78 == out_payload_rob_idx[6:0] ? rob_payload_120_tsc : _GEN_4216; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4218 = 7'h79 == out_payload_rob_idx[6:0] ? rob_payload_121_tsc : _GEN_4217; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4219 = 7'h7a == out_payload_rob_idx[6:0] ? rob_payload_122_tsc : _GEN_4218; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4220 = 7'h7b == out_payload_rob_idx[6:0] ? rob_payload_123_tsc : _GEN_4219; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4221 = 7'h7c == out_payload_rob_idx[6:0] ? rob_payload_124_tsc : _GEN_4220; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4222 = 7'h7d == out_payload_rob_idx[6:0] ? rob_payload_125_tsc : _GEN_4221; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4223 = 7'h7e == out_payload_rob_idx[6:0] ? rob_payload_126_tsc : _GEN_4222; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_4224 = 7'h7f == out_payload_rob_idx[6:0] ? rob_payload_127_tsc : _GEN_4223; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4226 = 7'h1 == out_payload_rob_idx[6:0] ? rob_payload_1_rob_idx : rob_payload_0_rob_idx; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4227 = 7'h2 == out_payload_rob_idx[6:0] ? rob_payload_2_rob_idx : _GEN_4226; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4228 = 7'h3 == out_payload_rob_idx[6:0] ? rob_payload_3_rob_idx : _GEN_4227; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4229 = 7'h4 == out_payload_rob_idx[6:0] ? rob_payload_4_rob_idx : _GEN_4228; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4230 = 7'h5 == out_payload_rob_idx[6:0] ? rob_payload_5_rob_idx : _GEN_4229; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4231 = 7'h6 == out_payload_rob_idx[6:0] ? rob_payload_6_rob_idx : _GEN_4230; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4232 = 7'h7 == out_payload_rob_idx[6:0] ? rob_payload_7_rob_idx : _GEN_4231; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4233 = 7'h8 == out_payload_rob_idx[6:0] ? rob_payload_8_rob_idx : _GEN_4232; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4234 = 7'h9 == out_payload_rob_idx[6:0] ? rob_payload_9_rob_idx : _GEN_4233; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4235 = 7'ha == out_payload_rob_idx[6:0] ? rob_payload_10_rob_idx : _GEN_4234; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4236 = 7'hb == out_payload_rob_idx[6:0] ? rob_payload_11_rob_idx : _GEN_4235; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4237 = 7'hc == out_payload_rob_idx[6:0] ? rob_payload_12_rob_idx : _GEN_4236; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4238 = 7'hd == out_payload_rob_idx[6:0] ? rob_payload_13_rob_idx : _GEN_4237; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4239 = 7'he == out_payload_rob_idx[6:0] ? rob_payload_14_rob_idx : _GEN_4238; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4240 = 7'hf == out_payload_rob_idx[6:0] ? rob_payload_15_rob_idx : _GEN_4239; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4241 = 7'h10 == out_payload_rob_idx[6:0] ? rob_payload_16_rob_idx : _GEN_4240; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4242 = 7'h11 == out_payload_rob_idx[6:0] ? rob_payload_17_rob_idx : _GEN_4241; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4243 = 7'h12 == out_payload_rob_idx[6:0] ? rob_payload_18_rob_idx : _GEN_4242; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4244 = 7'h13 == out_payload_rob_idx[6:0] ? rob_payload_19_rob_idx : _GEN_4243; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4245 = 7'h14 == out_payload_rob_idx[6:0] ? rob_payload_20_rob_idx : _GEN_4244; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4246 = 7'h15 == out_payload_rob_idx[6:0] ? rob_payload_21_rob_idx : _GEN_4245; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4247 = 7'h16 == out_payload_rob_idx[6:0] ? rob_payload_22_rob_idx : _GEN_4246; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4248 = 7'h17 == out_payload_rob_idx[6:0] ? rob_payload_23_rob_idx : _GEN_4247; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4249 = 7'h18 == out_payload_rob_idx[6:0] ? rob_payload_24_rob_idx : _GEN_4248; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4250 = 7'h19 == out_payload_rob_idx[6:0] ? rob_payload_25_rob_idx : _GEN_4249; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4251 = 7'h1a == out_payload_rob_idx[6:0] ? rob_payload_26_rob_idx : _GEN_4250; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4252 = 7'h1b == out_payload_rob_idx[6:0] ? rob_payload_27_rob_idx : _GEN_4251; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4253 = 7'h1c == out_payload_rob_idx[6:0] ? rob_payload_28_rob_idx : _GEN_4252; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4254 = 7'h1d == out_payload_rob_idx[6:0] ? rob_payload_29_rob_idx : _GEN_4253; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4255 = 7'h1e == out_payload_rob_idx[6:0] ? rob_payload_30_rob_idx : _GEN_4254; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4256 = 7'h1f == out_payload_rob_idx[6:0] ? rob_payload_31_rob_idx : _GEN_4255; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4257 = 7'h20 == out_payload_rob_idx[6:0] ? rob_payload_32_rob_idx : _GEN_4256; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4258 = 7'h21 == out_payload_rob_idx[6:0] ? rob_payload_33_rob_idx : _GEN_4257; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4259 = 7'h22 == out_payload_rob_idx[6:0] ? rob_payload_34_rob_idx : _GEN_4258; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4260 = 7'h23 == out_payload_rob_idx[6:0] ? rob_payload_35_rob_idx : _GEN_4259; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4261 = 7'h24 == out_payload_rob_idx[6:0] ? rob_payload_36_rob_idx : _GEN_4260; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4262 = 7'h25 == out_payload_rob_idx[6:0] ? rob_payload_37_rob_idx : _GEN_4261; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4263 = 7'h26 == out_payload_rob_idx[6:0] ? rob_payload_38_rob_idx : _GEN_4262; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4264 = 7'h27 == out_payload_rob_idx[6:0] ? rob_payload_39_rob_idx : _GEN_4263; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4265 = 7'h28 == out_payload_rob_idx[6:0] ? rob_payload_40_rob_idx : _GEN_4264; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4266 = 7'h29 == out_payload_rob_idx[6:0] ? rob_payload_41_rob_idx : _GEN_4265; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4267 = 7'h2a == out_payload_rob_idx[6:0] ? rob_payload_42_rob_idx : _GEN_4266; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4268 = 7'h2b == out_payload_rob_idx[6:0] ? rob_payload_43_rob_idx : _GEN_4267; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4269 = 7'h2c == out_payload_rob_idx[6:0] ? rob_payload_44_rob_idx : _GEN_4268; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4270 = 7'h2d == out_payload_rob_idx[6:0] ? rob_payload_45_rob_idx : _GEN_4269; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4271 = 7'h2e == out_payload_rob_idx[6:0] ? rob_payload_46_rob_idx : _GEN_4270; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4272 = 7'h2f == out_payload_rob_idx[6:0] ? rob_payload_47_rob_idx : _GEN_4271; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4273 = 7'h30 == out_payload_rob_idx[6:0] ? rob_payload_48_rob_idx : _GEN_4272; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4274 = 7'h31 == out_payload_rob_idx[6:0] ? rob_payload_49_rob_idx : _GEN_4273; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4275 = 7'h32 == out_payload_rob_idx[6:0] ? rob_payload_50_rob_idx : _GEN_4274; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4276 = 7'h33 == out_payload_rob_idx[6:0] ? rob_payload_51_rob_idx : _GEN_4275; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4277 = 7'h34 == out_payload_rob_idx[6:0] ? rob_payload_52_rob_idx : _GEN_4276; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4278 = 7'h35 == out_payload_rob_idx[6:0] ? rob_payload_53_rob_idx : _GEN_4277; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4279 = 7'h36 == out_payload_rob_idx[6:0] ? rob_payload_54_rob_idx : _GEN_4278; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4280 = 7'h37 == out_payload_rob_idx[6:0] ? rob_payload_55_rob_idx : _GEN_4279; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4281 = 7'h38 == out_payload_rob_idx[6:0] ? rob_payload_56_rob_idx : _GEN_4280; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4282 = 7'h39 == out_payload_rob_idx[6:0] ? rob_payload_57_rob_idx : _GEN_4281; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4283 = 7'h3a == out_payload_rob_idx[6:0] ? rob_payload_58_rob_idx : _GEN_4282; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4284 = 7'h3b == out_payload_rob_idx[6:0] ? rob_payload_59_rob_idx : _GEN_4283; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4285 = 7'h3c == out_payload_rob_idx[6:0] ? rob_payload_60_rob_idx : _GEN_4284; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4286 = 7'h3d == out_payload_rob_idx[6:0] ? rob_payload_61_rob_idx : _GEN_4285; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4287 = 7'h3e == out_payload_rob_idx[6:0] ? rob_payload_62_rob_idx : _GEN_4286; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4288 = 7'h3f == out_payload_rob_idx[6:0] ? rob_payload_63_rob_idx : _GEN_4287; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4289 = 7'h40 == out_payload_rob_idx[6:0] ? rob_payload_64_rob_idx : _GEN_4288; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4290 = 7'h41 == out_payload_rob_idx[6:0] ? rob_payload_65_rob_idx : _GEN_4289; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4291 = 7'h42 == out_payload_rob_idx[6:0] ? rob_payload_66_rob_idx : _GEN_4290; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4292 = 7'h43 == out_payload_rob_idx[6:0] ? rob_payload_67_rob_idx : _GEN_4291; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4293 = 7'h44 == out_payload_rob_idx[6:0] ? rob_payload_68_rob_idx : _GEN_4292; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4294 = 7'h45 == out_payload_rob_idx[6:0] ? rob_payload_69_rob_idx : _GEN_4293; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4295 = 7'h46 == out_payload_rob_idx[6:0] ? rob_payload_70_rob_idx : _GEN_4294; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4296 = 7'h47 == out_payload_rob_idx[6:0] ? rob_payload_71_rob_idx : _GEN_4295; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4297 = 7'h48 == out_payload_rob_idx[6:0] ? rob_payload_72_rob_idx : _GEN_4296; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4298 = 7'h49 == out_payload_rob_idx[6:0] ? rob_payload_73_rob_idx : _GEN_4297; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4299 = 7'h4a == out_payload_rob_idx[6:0] ? rob_payload_74_rob_idx : _GEN_4298; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4300 = 7'h4b == out_payload_rob_idx[6:0] ? rob_payload_75_rob_idx : _GEN_4299; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4301 = 7'h4c == out_payload_rob_idx[6:0] ? rob_payload_76_rob_idx : _GEN_4300; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4302 = 7'h4d == out_payload_rob_idx[6:0] ? rob_payload_77_rob_idx : _GEN_4301; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4303 = 7'h4e == out_payload_rob_idx[6:0] ? rob_payload_78_rob_idx : _GEN_4302; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4304 = 7'h4f == out_payload_rob_idx[6:0] ? rob_payload_79_rob_idx : _GEN_4303; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4305 = 7'h50 == out_payload_rob_idx[6:0] ? rob_payload_80_rob_idx : _GEN_4304; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4306 = 7'h51 == out_payload_rob_idx[6:0] ? rob_payload_81_rob_idx : _GEN_4305; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4307 = 7'h52 == out_payload_rob_idx[6:0] ? rob_payload_82_rob_idx : _GEN_4306; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4308 = 7'h53 == out_payload_rob_idx[6:0] ? rob_payload_83_rob_idx : _GEN_4307; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4309 = 7'h54 == out_payload_rob_idx[6:0] ? rob_payload_84_rob_idx : _GEN_4308; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4310 = 7'h55 == out_payload_rob_idx[6:0] ? rob_payload_85_rob_idx : _GEN_4309; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4311 = 7'h56 == out_payload_rob_idx[6:0] ? rob_payload_86_rob_idx : _GEN_4310; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4312 = 7'h57 == out_payload_rob_idx[6:0] ? rob_payload_87_rob_idx : _GEN_4311; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4313 = 7'h58 == out_payload_rob_idx[6:0] ? rob_payload_88_rob_idx : _GEN_4312; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4314 = 7'h59 == out_payload_rob_idx[6:0] ? rob_payload_89_rob_idx : _GEN_4313; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4315 = 7'h5a == out_payload_rob_idx[6:0] ? rob_payload_90_rob_idx : _GEN_4314; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4316 = 7'h5b == out_payload_rob_idx[6:0] ? rob_payload_91_rob_idx : _GEN_4315; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4317 = 7'h5c == out_payload_rob_idx[6:0] ? rob_payload_92_rob_idx : _GEN_4316; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4318 = 7'h5d == out_payload_rob_idx[6:0] ? rob_payload_93_rob_idx : _GEN_4317; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4319 = 7'h5e == out_payload_rob_idx[6:0] ? rob_payload_94_rob_idx : _GEN_4318; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4320 = 7'h5f == out_payload_rob_idx[6:0] ? rob_payload_95_rob_idx : _GEN_4319; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4321 = 7'h60 == out_payload_rob_idx[6:0] ? rob_payload_96_rob_idx : _GEN_4320; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4322 = 7'h61 == out_payload_rob_idx[6:0] ? rob_payload_97_rob_idx : _GEN_4321; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4323 = 7'h62 == out_payload_rob_idx[6:0] ? rob_payload_98_rob_idx : _GEN_4322; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4324 = 7'h63 == out_payload_rob_idx[6:0] ? rob_payload_99_rob_idx : _GEN_4323; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4325 = 7'h64 == out_payload_rob_idx[6:0] ? rob_payload_100_rob_idx : _GEN_4324; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4326 = 7'h65 == out_payload_rob_idx[6:0] ? rob_payload_101_rob_idx : _GEN_4325; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4327 = 7'h66 == out_payload_rob_idx[6:0] ? rob_payload_102_rob_idx : _GEN_4326; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4328 = 7'h67 == out_payload_rob_idx[6:0] ? rob_payload_103_rob_idx : _GEN_4327; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4329 = 7'h68 == out_payload_rob_idx[6:0] ? rob_payload_104_rob_idx : _GEN_4328; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4330 = 7'h69 == out_payload_rob_idx[6:0] ? rob_payload_105_rob_idx : _GEN_4329; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4331 = 7'h6a == out_payload_rob_idx[6:0] ? rob_payload_106_rob_idx : _GEN_4330; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4332 = 7'h6b == out_payload_rob_idx[6:0] ? rob_payload_107_rob_idx : _GEN_4331; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4333 = 7'h6c == out_payload_rob_idx[6:0] ? rob_payload_108_rob_idx : _GEN_4332; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4334 = 7'h6d == out_payload_rob_idx[6:0] ? rob_payload_109_rob_idx : _GEN_4333; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4335 = 7'h6e == out_payload_rob_idx[6:0] ? rob_payload_110_rob_idx : _GEN_4334; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4336 = 7'h6f == out_payload_rob_idx[6:0] ? rob_payload_111_rob_idx : _GEN_4335; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4337 = 7'h70 == out_payload_rob_idx[6:0] ? rob_payload_112_rob_idx : _GEN_4336; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4338 = 7'h71 == out_payload_rob_idx[6:0] ? rob_payload_113_rob_idx : _GEN_4337; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4339 = 7'h72 == out_payload_rob_idx[6:0] ? rob_payload_114_rob_idx : _GEN_4338; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4340 = 7'h73 == out_payload_rob_idx[6:0] ? rob_payload_115_rob_idx : _GEN_4339; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4341 = 7'h74 == out_payload_rob_idx[6:0] ? rob_payload_116_rob_idx : _GEN_4340; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4342 = 7'h75 == out_payload_rob_idx[6:0] ? rob_payload_117_rob_idx : _GEN_4341; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4343 = 7'h76 == out_payload_rob_idx[6:0] ? rob_payload_118_rob_idx : _GEN_4342; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4344 = 7'h77 == out_payload_rob_idx[6:0] ? rob_payload_119_rob_idx : _GEN_4343; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4345 = 7'h78 == out_payload_rob_idx[6:0] ? rob_payload_120_rob_idx : _GEN_4344; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4346 = 7'h79 == out_payload_rob_idx[6:0] ? rob_payload_121_rob_idx : _GEN_4345; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4347 = 7'h7a == out_payload_rob_idx[6:0] ? rob_payload_122_rob_idx : _GEN_4346; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4348 = 7'h7b == out_payload_rob_idx[6:0] ? rob_payload_123_rob_idx : _GEN_4347; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4349 = 7'h7c == out_payload_rob_idx[6:0] ? rob_payload_124_rob_idx : _GEN_4348; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4350 = 7'h7d == out_payload_rob_idx[6:0] ? rob_payload_125_rob_idx : _GEN_4349; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4351 = 7'h7e == out_payload_rob_idx[6:0] ? rob_payload_126_rob_idx : _GEN_4350; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4352 = 7'h7f == out_payload_rob_idx[6:0] ? rob_payload_127_rob_idx : _GEN_4351; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4354 = 7'h1 == out_payload_rob_idx[6:0] ? rob_payload_1_flits_fired : rob_payload_0_flits_fired; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4355 = 7'h2 == out_payload_rob_idx[6:0] ? rob_payload_2_flits_fired : _GEN_4354; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4356 = 7'h3 == out_payload_rob_idx[6:0] ? rob_payload_3_flits_fired : _GEN_4355; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4357 = 7'h4 == out_payload_rob_idx[6:0] ? rob_payload_4_flits_fired : _GEN_4356; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4358 = 7'h5 == out_payload_rob_idx[6:0] ? rob_payload_5_flits_fired : _GEN_4357; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4359 = 7'h6 == out_payload_rob_idx[6:0] ? rob_payload_6_flits_fired : _GEN_4358; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4360 = 7'h7 == out_payload_rob_idx[6:0] ? rob_payload_7_flits_fired : _GEN_4359; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4361 = 7'h8 == out_payload_rob_idx[6:0] ? rob_payload_8_flits_fired : _GEN_4360; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4362 = 7'h9 == out_payload_rob_idx[6:0] ? rob_payload_9_flits_fired : _GEN_4361; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4363 = 7'ha == out_payload_rob_idx[6:0] ? rob_payload_10_flits_fired : _GEN_4362; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4364 = 7'hb == out_payload_rob_idx[6:0] ? rob_payload_11_flits_fired : _GEN_4363; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4365 = 7'hc == out_payload_rob_idx[6:0] ? rob_payload_12_flits_fired : _GEN_4364; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4366 = 7'hd == out_payload_rob_idx[6:0] ? rob_payload_13_flits_fired : _GEN_4365; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4367 = 7'he == out_payload_rob_idx[6:0] ? rob_payload_14_flits_fired : _GEN_4366; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4368 = 7'hf == out_payload_rob_idx[6:0] ? rob_payload_15_flits_fired : _GEN_4367; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4369 = 7'h10 == out_payload_rob_idx[6:0] ? rob_payload_16_flits_fired : _GEN_4368; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4370 = 7'h11 == out_payload_rob_idx[6:0] ? rob_payload_17_flits_fired : _GEN_4369; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4371 = 7'h12 == out_payload_rob_idx[6:0] ? rob_payload_18_flits_fired : _GEN_4370; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4372 = 7'h13 == out_payload_rob_idx[6:0] ? rob_payload_19_flits_fired : _GEN_4371; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4373 = 7'h14 == out_payload_rob_idx[6:0] ? rob_payload_20_flits_fired : _GEN_4372; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4374 = 7'h15 == out_payload_rob_idx[6:0] ? rob_payload_21_flits_fired : _GEN_4373; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4375 = 7'h16 == out_payload_rob_idx[6:0] ? rob_payload_22_flits_fired : _GEN_4374; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4376 = 7'h17 == out_payload_rob_idx[6:0] ? rob_payload_23_flits_fired : _GEN_4375; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4377 = 7'h18 == out_payload_rob_idx[6:0] ? rob_payload_24_flits_fired : _GEN_4376; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4378 = 7'h19 == out_payload_rob_idx[6:0] ? rob_payload_25_flits_fired : _GEN_4377; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4379 = 7'h1a == out_payload_rob_idx[6:0] ? rob_payload_26_flits_fired : _GEN_4378; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4380 = 7'h1b == out_payload_rob_idx[6:0] ? rob_payload_27_flits_fired : _GEN_4379; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4381 = 7'h1c == out_payload_rob_idx[6:0] ? rob_payload_28_flits_fired : _GEN_4380; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4382 = 7'h1d == out_payload_rob_idx[6:0] ? rob_payload_29_flits_fired : _GEN_4381; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4383 = 7'h1e == out_payload_rob_idx[6:0] ? rob_payload_30_flits_fired : _GEN_4382; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4384 = 7'h1f == out_payload_rob_idx[6:0] ? rob_payload_31_flits_fired : _GEN_4383; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4385 = 7'h20 == out_payload_rob_idx[6:0] ? rob_payload_32_flits_fired : _GEN_4384; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4386 = 7'h21 == out_payload_rob_idx[6:0] ? rob_payload_33_flits_fired : _GEN_4385; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4387 = 7'h22 == out_payload_rob_idx[6:0] ? rob_payload_34_flits_fired : _GEN_4386; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4388 = 7'h23 == out_payload_rob_idx[6:0] ? rob_payload_35_flits_fired : _GEN_4387; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4389 = 7'h24 == out_payload_rob_idx[6:0] ? rob_payload_36_flits_fired : _GEN_4388; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4390 = 7'h25 == out_payload_rob_idx[6:0] ? rob_payload_37_flits_fired : _GEN_4389; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4391 = 7'h26 == out_payload_rob_idx[6:0] ? rob_payload_38_flits_fired : _GEN_4390; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4392 = 7'h27 == out_payload_rob_idx[6:0] ? rob_payload_39_flits_fired : _GEN_4391; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4393 = 7'h28 == out_payload_rob_idx[6:0] ? rob_payload_40_flits_fired : _GEN_4392; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4394 = 7'h29 == out_payload_rob_idx[6:0] ? rob_payload_41_flits_fired : _GEN_4393; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4395 = 7'h2a == out_payload_rob_idx[6:0] ? rob_payload_42_flits_fired : _GEN_4394; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4396 = 7'h2b == out_payload_rob_idx[6:0] ? rob_payload_43_flits_fired : _GEN_4395; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4397 = 7'h2c == out_payload_rob_idx[6:0] ? rob_payload_44_flits_fired : _GEN_4396; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4398 = 7'h2d == out_payload_rob_idx[6:0] ? rob_payload_45_flits_fired : _GEN_4397; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4399 = 7'h2e == out_payload_rob_idx[6:0] ? rob_payload_46_flits_fired : _GEN_4398; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4400 = 7'h2f == out_payload_rob_idx[6:0] ? rob_payload_47_flits_fired : _GEN_4399; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4401 = 7'h30 == out_payload_rob_idx[6:0] ? rob_payload_48_flits_fired : _GEN_4400; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4402 = 7'h31 == out_payload_rob_idx[6:0] ? rob_payload_49_flits_fired : _GEN_4401; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4403 = 7'h32 == out_payload_rob_idx[6:0] ? rob_payload_50_flits_fired : _GEN_4402; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4404 = 7'h33 == out_payload_rob_idx[6:0] ? rob_payload_51_flits_fired : _GEN_4403; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4405 = 7'h34 == out_payload_rob_idx[6:0] ? rob_payload_52_flits_fired : _GEN_4404; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4406 = 7'h35 == out_payload_rob_idx[6:0] ? rob_payload_53_flits_fired : _GEN_4405; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4407 = 7'h36 == out_payload_rob_idx[6:0] ? rob_payload_54_flits_fired : _GEN_4406; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4408 = 7'h37 == out_payload_rob_idx[6:0] ? rob_payload_55_flits_fired : _GEN_4407; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4409 = 7'h38 == out_payload_rob_idx[6:0] ? rob_payload_56_flits_fired : _GEN_4408; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4410 = 7'h39 == out_payload_rob_idx[6:0] ? rob_payload_57_flits_fired : _GEN_4409; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4411 = 7'h3a == out_payload_rob_idx[6:0] ? rob_payload_58_flits_fired : _GEN_4410; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4412 = 7'h3b == out_payload_rob_idx[6:0] ? rob_payload_59_flits_fired : _GEN_4411; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4413 = 7'h3c == out_payload_rob_idx[6:0] ? rob_payload_60_flits_fired : _GEN_4412; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4414 = 7'h3d == out_payload_rob_idx[6:0] ? rob_payload_61_flits_fired : _GEN_4413; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4415 = 7'h3e == out_payload_rob_idx[6:0] ? rob_payload_62_flits_fired : _GEN_4414; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4416 = 7'h3f == out_payload_rob_idx[6:0] ? rob_payload_63_flits_fired : _GEN_4415; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4417 = 7'h40 == out_payload_rob_idx[6:0] ? rob_payload_64_flits_fired : _GEN_4416; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4418 = 7'h41 == out_payload_rob_idx[6:0] ? rob_payload_65_flits_fired : _GEN_4417; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4419 = 7'h42 == out_payload_rob_idx[6:0] ? rob_payload_66_flits_fired : _GEN_4418; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4420 = 7'h43 == out_payload_rob_idx[6:0] ? rob_payload_67_flits_fired : _GEN_4419; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4421 = 7'h44 == out_payload_rob_idx[6:0] ? rob_payload_68_flits_fired : _GEN_4420; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4422 = 7'h45 == out_payload_rob_idx[6:0] ? rob_payload_69_flits_fired : _GEN_4421; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4423 = 7'h46 == out_payload_rob_idx[6:0] ? rob_payload_70_flits_fired : _GEN_4422; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4424 = 7'h47 == out_payload_rob_idx[6:0] ? rob_payload_71_flits_fired : _GEN_4423; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4425 = 7'h48 == out_payload_rob_idx[6:0] ? rob_payload_72_flits_fired : _GEN_4424; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4426 = 7'h49 == out_payload_rob_idx[6:0] ? rob_payload_73_flits_fired : _GEN_4425; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4427 = 7'h4a == out_payload_rob_idx[6:0] ? rob_payload_74_flits_fired : _GEN_4426; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4428 = 7'h4b == out_payload_rob_idx[6:0] ? rob_payload_75_flits_fired : _GEN_4427; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4429 = 7'h4c == out_payload_rob_idx[6:0] ? rob_payload_76_flits_fired : _GEN_4428; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4430 = 7'h4d == out_payload_rob_idx[6:0] ? rob_payload_77_flits_fired : _GEN_4429; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4431 = 7'h4e == out_payload_rob_idx[6:0] ? rob_payload_78_flits_fired : _GEN_4430; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4432 = 7'h4f == out_payload_rob_idx[6:0] ? rob_payload_79_flits_fired : _GEN_4431; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4433 = 7'h50 == out_payload_rob_idx[6:0] ? rob_payload_80_flits_fired : _GEN_4432; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4434 = 7'h51 == out_payload_rob_idx[6:0] ? rob_payload_81_flits_fired : _GEN_4433; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4435 = 7'h52 == out_payload_rob_idx[6:0] ? rob_payload_82_flits_fired : _GEN_4434; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4436 = 7'h53 == out_payload_rob_idx[6:0] ? rob_payload_83_flits_fired : _GEN_4435; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4437 = 7'h54 == out_payload_rob_idx[6:0] ? rob_payload_84_flits_fired : _GEN_4436; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4438 = 7'h55 == out_payload_rob_idx[6:0] ? rob_payload_85_flits_fired : _GEN_4437; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4439 = 7'h56 == out_payload_rob_idx[6:0] ? rob_payload_86_flits_fired : _GEN_4438; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4440 = 7'h57 == out_payload_rob_idx[6:0] ? rob_payload_87_flits_fired : _GEN_4439; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4441 = 7'h58 == out_payload_rob_idx[6:0] ? rob_payload_88_flits_fired : _GEN_4440; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4442 = 7'h59 == out_payload_rob_idx[6:0] ? rob_payload_89_flits_fired : _GEN_4441; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4443 = 7'h5a == out_payload_rob_idx[6:0] ? rob_payload_90_flits_fired : _GEN_4442; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4444 = 7'h5b == out_payload_rob_idx[6:0] ? rob_payload_91_flits_fired : _GEN_4443; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4445 = 7'h5c == out_payload_rob_idx[6:0] ? rob_payload_92_flits_fired : _GEN_4444; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4446 = 7'h5d == out_payload_rob_idx[6:0] ? rob_payload_93_flits_fired : _GEN_4445; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4447 = 7'h5e == out_payload_rob_idx[6:0] ? rob_payload_94_flits_fired : _GEN_4446; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4448 = 7'h5f == out_payload_rob_idx[6:0] ? rob_payload_95_flits_fired : _GEN_4447; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4449 = 7'h60 == out_payload_rob_idx[6:0] ? rob_payload_96_flits_fired : _GEN_4448; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4450 = 7'h61 == out_payload_rob_idx[6:0] ? rob_payload_97_flits_fired : _GEN_4449; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4451 = 7'h62 == out_payload_rob_idx[6:0] ? rob_payload_98_flits_fired : _GEN_4450; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4452 = 7'h63 == out_payload_rob_idx[6:0] ? rob_payload_99_flits_fired : _GEN_4451; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4453 = 7'h64 == out_payload_rob_idx[6:0] ? rob_payload_100_flits_fired : _GEN_4452; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4454 = 7'h65 == out_payload_rob_idx[6:0] ? rob_payload_101_flits_fired : _GEN_4453; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4455 = 7'h66 == out_payload_rob_idx[6:0] ? rob_payload_102_flits_fired : _GEN_4454; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4456 = 7'h67 == out_payload_rob_idx[6:0] ? rob_payload_103_flits_fired : _GEN_4455; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4457 = 7'h68 == out_payload_rob_idx[6:0] ? rob_payload_104_flits_fired : _GEN_4456; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4458 = 7'h69 == out_payload_rob_idx[6:0] ? rob_payload_105_flits_fired : _GEN_4457; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4459 = 7'h6a == out_payload_rob_idx[6:0] ? rob_payload_106_flits_fired : _GEN_4458; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4460 = 7'h6b == out_payload_rob_idx[6:0] ? rob_payload_107_flits_fired : _GEN_4459; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4461 = 7'h6c == out_payload_rob_idx[6:0] ? rob_payload_108_flits_fired : _GEN_4460; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4462 = 7'h6d == out_payload_rob_idx[6:0] ? rob_payload_109_flits_fired : _GEN_4461; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4463 = 7'h6e == out_payload_rob_idx[6:0] ? rob_payload_110_flits_fired : _GEN_4462; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4464 = 7'h6f == out_payload_rob_idx[6:0] ? rob_payload_111_flits_fired : _GEN_4463; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4465 = 7'h70 == out_payload_rob_idx[6:0] ? rob_payload_112_flits_fired : _GEN_4464; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4466 = 7'h71 == out_payload_rob_idx[6:0] ? rob_payload_113_flits_fired : _GEN_4465; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4467 = 7'h72 == out_payload_rob_idx[6:0] ? rob_payload_114_flits_fired : _GEN_4466; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4468 = 7'h73 == out_payload_rob_idx[6:0] ? rob_payload_115_flits_fired : _GEN_4467; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4469 = 7'h74 == out_payload_rob_idx[6:0] ? rob_payload_116_flits_fired : _GEN_4468; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4470 = 7'h75 == out_payload_rob_idx[6:0] ? rob_payload_117_flits_fired : _GEN_4469; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4471 = 7'h76 == out_payload_rob_idx[6:0] ? rob_payload_118_flits_fired : _GEN_4470; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4472 = 7'h77 == out_payload_rob_idx[6:0] ? rob_payload_119_flits_fired : _GEN_4471; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4473 = 7'h78 == out_payload_rob_idx[6:0] ? rob_payload_120_flits_fired : _GEN_4472; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4474 = 7'h79 == out_payload_rob_idx[6:0] ? rob_payload_121_flits_fired : _GEN_4473; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4475 = 7'h7a == out_payload_rob_idx[6:0] ? rob_payload_122_flits_fired : _GEN_4474; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4476 = 7'h7b == out_payload_rob_idx[6:0] ? rob_payload_123_flits_fired : _GEN_4475; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4477 = 7'h7c == out_payload_rob_idx[6:0] ? rob_payload_124_flits_fired : _GEN_4476; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4478 = 7'h7d == out_payload_rob_idx[6:0] ? rob_payload_125_flits_fired : _GEN_4477; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4479 = 7'h7e == out_payload_rob_idx[6:0] ? rob_payload_126_flits_fired : _GEN_4478; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_4480 = 7'h7f == out_payload_rob_idx[6:0] ? rob_payload_127_flits_fired : _GEN_4479; // @[TestHarness.scala 202:{35,35}]
  wire [63:0] _T_48 = {_GEN_4224,_GEN_4352,_GEN_4480}; // @[TestHarness.scala 202:35]
  wire  _GEN_4482 = 7'h1 == out_payload_rob_idx[6:0] ? rob_ingress_id_1 : rob_ingress_id_0; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4483 = 7'h2 == out_payload_rob_idx[6:0] ? rob_ingress_id_2 : _GEN_4482; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4484 = 7'h3 == out_payload_rob_idx[6:0] ? rob_ingress_id_3 : _GEN_4483; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4485 = 7'h4 == out_payload_rob_idx[6:0] ? rob_ingress_id_4 : _GEN_4484; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4486 = 7'h5 == out_payload_rob_idx[6:0] ? rob_ingress_id_5 : _GEN_4485; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4487 = 7'h6 == out_payload_rob_idx[6:0] ? rob_ingress_id_6 : _GEN_4486; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4488 = 7'h7 == out_payload_rob_idx[6:0] ? rob_ingress_id_7 : _GEN_4487; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4489 = 7'h8 == out_payload_rob_idx[6:0] ? rob_ingress_id_8 : _GEN_4488; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4490 = 7'h9 == out_payload_rob_idx[6:0] ? rob_ingress_id_9 : _GEN_4489; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4491 = 7'ha == out_payload_rob_idx[6:0] ? rob_ingress_id_10 : _GEN_4490; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4492 = 7'hb == out_payload_rob_idx[6:0] ? rob_ingress_id_11 : _GEN_4491; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4493 = 7'hc == out_payload_rob_idx[6:0] ? rob_ingress_id_12 : _GEN_4492; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4494 = 7'hd == out_payload_rob_idx[6:0] ? rob_ingress_id_13 : _GEN_4493; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4495 = 7'he == out_payload_rob_idx[6:0] ? rob_ingress_id_14 : _GEN_4494; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4496 = 7'hf == out_payload_rob_idx[6:0] ? rob_ingress_id_15 : _GEN_4495; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4497 = 7'h10 == out_payload_rob_idx[6:0] ? rob_ingress_id_16 : _GEN_4496; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4498 = 7'h11 == out_payload_rob_idx[6:0] ? rob_ingress_id_17 : _GEN_4497; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4499 = 7'h12 == out_payload_rob_idx[6:0] ? rob_ingress_id_18 : _GEN_4498; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4500 = 7'h13 == out_payload_rob_idx[6:0] ? rob_ingress_id_19 : _GEN_4499; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4501 = 7'h14 == out_payload_rob_idx[6:0] ? rob_ingress_id_20 : _GEN_4500; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4502 = 7'h15 == out_payload_rob_idx[6:0] ? rob_ingress_id_21 : _GEN_4501; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4503 = 7'h16 == out_payload_rob_idx[6:0] ? rob_ingress_id_22 : _GEN_4502; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4504 = 7'h17 == out_payload_rob_idx[6:0] ? rob_ingress_id_23 : _GEN_4503; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4505 = 7'h18 == out_payload_rob_idx[6:0] ? rob_ingress_id_24 : _GEN_4504; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4506 = 7'h19 == out_payload_rob_idx[6:0] ? rob_ingress_id_25 : _GEN_4505; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4507 = 7'h1a == out_payload_rob_idx[6:0] ? rob_ingress_id_26 : _GEN_4506; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4508 = 7'h1b == out_payload_rob_idx[6:0] ? rob_ingress_id_27 : _GEN_4507; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4509 = 7'h1c == out_payload_rob_idx[6:0] ? rob_ingress_id_28 : _GEN_4508; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4510 = 7'h1d == out_payload_rob_idx[6:0] ? rob_ingress_id_29 : _GEN_4509; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4511 = 7'h1e == out_payload_rob_idx[6:0] ? rob_ingress_id_30 : _GEN_4510; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4512 = 7'h1f == out_payload_rob_idx[6:0] ? rob_ingress_id_31 : _GEN_4511; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4513 = 7'h20 == out_payload_rob_idx[6:0] ? rob_ingress_id_32 : _GEN_4512; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4514 = 7'h21 == out_payload_rob_idx[6:0] ? rob_ingress_id_33 : _GEN_4513; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4515 = 7'h22 == out_payload_rob_idx[6:0] ? rob_ingress_id_34 : _GEN_4514; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4516 = 7'h23 == out_payload_rob_idx[6:0] ? rob_ingress_id_35 : _GEN_4515; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4517 = 7'h24 == out_payload_rob_idx[6:0] ? rob_ingress_id_36 : _GEN_4516; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4518 = 7'h25 == out_payload_rob_idx[6:0] ? rob_ingress_id_37 : _GEN_4517; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4519 = 7'h26 == out_payload_rob_idx[6:0] ? rob_ingress_id_38 : _GEN_4518; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4520 = 7'h27 == out_payload_rob_idx[6:0] ? rob_ingress_id_39 : _GEN_4519; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4521 = 7'h28 == out_payload_rob_idx[6:0] ? rob_ingress_id_40 : _GEN_4520; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4522 = 7'h29 == out_payload_rob_idx[6:0] ? rob_ingress_id_41 : _GEN_4521; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4523 = 7'h2a == out_payload_rob_idx[6:0] ? rob_ingress_id_42 : _GEN_4522; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4524 = 7'h2b == out_payload_rob_idx[6:0] ? rob_ingress_id_43 : _GEN_4523; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4525 = 7'h2c == out_payload_rob_idx[6:0] ? rob_ingress_id_44 : _GEN_4524; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4526 = 7'h2d == out_payload_rob_idx[6:0] ? rob_ingress_id_45 : _GEN_4525; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4527 = 7'h2e == out_payload_rob_idx[6:0] ? rob_ingress_id_46 : _GEN_4526; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4528 = 7'h2f == out_payload_rob_idx[6:0] ? rob_ingress_id_47 : _GEN_4527; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4529 = 7'h30 == out_payload_rob_idx[6:0] ? rob_ingress_id_48 : _GEN_4528; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4530 = 7'h31 == out_payload_rob_idx[6:0] ? rob_ingress_id_49 : _GEN_4529; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4531 = 7'h32 == out_payload_rob_idx[6:0] ? rob_ingress_id_50 : _GEN_4530; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4532 = 7'h33 == out_payload_rob_idx[6:0] ? rob_ingress_id_51 : _GEN_4531; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4533 = 7'h34 == out_payload_rob_idx[6:0] ? rob_ingress_id_52 : _GEN_4532; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4534 = 7'h35 == out_payload_rob_idx[6:0] ? rob_ingress_id_53 : _GEN_4533; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4535 = 7'h36 == out_payload_rob_idx[6:0] ? rob_ingress_id_54 : _GEN_4534; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4536 = 7'h37 == out_payload_rob_idx[6:0] ? rob_ingress_id_55 : _GEN_4535; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4537 = 7'h38 == out_payload_rob_idx[6:0] ? rob_ingress_id_56 : _GEN_4536; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4538 = 7'h39 == out_payload_rob_idx[6:0] ? rob_ingress_id_57 : _GEN_4537; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4539 = 7'h3a == out_payload_rob_idx[6:0] ? rob_ingress_id_58 : _GEN_4538; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4540 = 7'h3b == out_payload_rob_idx[6:0] ? rob_ingress_id_59 : _GEN_4539; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4541 = 7'h3c == out_payload_rob_idx[6:0] ? rob_ingress_id_60 : _GEN_4540; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4542 = 7'h3d == out_payload_rob_idx[6:0] ? rob_ingress_id_61 : _GEN_4541; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4543 = 7'h3e == out_payload_rob_idx[6:0] ? rob_ingress_id_62 : _GEN_4542; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4544 = 7'h3f == out_payload_rob_idx[6:0] ? rob_ingress_id_63 : _GEN_4543; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4545 = 7'h40 == out_payload_rob_idx[6:0] ? rob_ingress_id_64 : _GEN_4544; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4546 = 7'h41 == out_payload_rob_idx[6:0] ? rob_ingress_id_65 : _GEN_4545; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4547 = 7'h42 == out_payload_rob_idx[6:0] ? rob_ingress_id_66 : _GEN_4546; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4548 = 7'h43 == out_payload_rob_idx[6:0] ? rob_ingress_id_67 : _GEN_4547; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4549 = 7'h44 == out_payload_rob_idx[6:0] ? rob_ingress_id_68 : _GEN_4548; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4550 = 7'h45 == out_payload_rob_idx[6:0] ? rob_ingress_id_69 : _GEN_4549; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4551 = 7'h46 == out_payload_rob_idx[6:0] ? rob_ingress_id_70 : _GEN_4550; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4552 = 7'h47 == out_payload_rob_idx[6:0] ? rob_ingress_id_71 : _GEN_4551; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4553 = 7'h48 == out_payload_rob_idx[6:0] ? rob_ingress_id_72 : _GEN_4552; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4554 = 7'h49 == out_payload_rob_idx[6:0] ? rob_ingress_id_73 : _GEN_4553; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4555 = 7'h4a == out_payload_rob_idx[6:0] ? rob_ingress_id_74 : _GEN_4554; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4556 = 7'h4b == out_payload_rob_idx[6:0] ? rob_ingress_id_75 : _GEN_4555; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4557 = 7'h4c == out_payload_rob_idx[6:0] ? rob_ingress_id_76 : _GEN_4556; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4558 = 7'h4d == out_payload_rob_idx[6:0] ? rob_ingress_id_77 : _GEN_4557; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4559 = 7'h4e == out_payload_rob_idx[6:0] ? rob_ingress_id_78 : _GEN_4558; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4560 = 7'h4f == out_payload_rob_idx[6:0] ? rob_ingress_id_79 : _GEN_4559; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4561 = 7'h50 == out_payload_rob_idx[6:0] ? rob_ingress_id_80 : _GEN_4560; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4562 = 7'h51 == out_payload_rob_idx[6:0] ? rob_ingress_id_81 : _GEN_4561; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4563 = 7'h52 == out_payload_rob_idx[6:0] ? rob_ingress_id_82 : _GEN_4562; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4564 = 7'h53 == out_payload_rob_idx[6:0] ? rob_ingress_id_83 : _GEN_4563; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4565 = 7'h54 == out_payload_rob_idx[6:0] ? rob_ingress_id_84 : _GEN_4564; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4566 = 7'h55 == out_payload_rob_idx[6:0] ? rob_ingress_id_85 : _GEN_4565; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4567 = 7'h56 == out_payload_rob_idx[6:0] ? rob_ingress_id_86 : _GEN_4566; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4568 = 7'h57 == out_payload_rob_idx[6:0] ? rob_ingress_id_87 : _GEN_4567; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4569 = 7'h58 == out_payload_rob_idx[6:0] ? rob_ingress_id_88 : _GEN_4568; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4570 = 7'h59 == out_payload_rob_idx[6:0] ? rob_ingress_id_89 : _GEN_4569; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4571 = 7'h5a == out_payload_rob_idx[6:0] ? rob_ingress_id_90 : _GEN_4570; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4572 = 7'h5b == out_payload_rob_idx[6:0] ? rob_ingress_id_91 : _GEN_4571; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4573 = 7'h5c == out_payload_rob_idx[6:0] ? rob_ingress_id_92 : _GEN_4572; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4574 = 7'h5d == out_payload_rob_idx[6:0] ? rob_ingress_id_93 : _GEN_4573; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4575 = 7'h5e == out_payload_rob_idx[6:0] ? rob_ingress_id_94 : _GEN_4574; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4576 = 7'h5f == out_payload_rob_idx[6:0] ? rob_ingress_id_95 : _GEN_4575; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4577 = 7'h60 == out_payload_rob_idx[6:0] ? rob_ingress_id_96 : _GEN_4576; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4578 = 7'h61 == out_payload_rob_idx[6:0] ? rob_ingress_id_97 : _GEN_4577; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4579 = 7'h62 == out_payload_rob_idx[6:0] ? rob_ingress_id_98 : _GEN_4578; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4580 = 7'h63 == out_payload_rob_idx[6:0] ? rob_ingress_id_99 : _GEN_4579; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4581 = 7'h64 == out_payload_rob_idx[6:0] ? rob_ingress_id_100 : _GEN_4580; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4582 = 7'h65 == out_payload_rob_idx[6:0] ? rob_ingress_id_101 : _GEN_4581; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4583 = 7'h66 == out_payload_rob_idx[6:0] ? rob_ingress_id_102 : _GEN_4582; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4584 = 7'h67 == out_payload_rob_idx[6:0] ? rob_ingress_id_103 : _GEN_4583; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4585 = 7'h68 == out_payload_rob_idx[6:0] ? rob_ingress_id_104 : _GEN_4584; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4586 = 7'h69 == out_payload_rob_idx[6:0] ? rob_ingress_id_105 : _GEN_4585; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4587 = 7'h6a == out_payload_rob_idx[6:0] ? rob_ingress_id_106 : _GEN_4586; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4588 = 7'h6b == out_payload_rob_idx[6:0] ? rob_ingress_id_107 : _GEN_4587; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4589 = 7'h6c == out_payload_rob_idx[6:0] ? rob_ingress_id_108 : _GEN_4588; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4590 = 7'h6d == out_payload_rob_idx[6:0] ? rob_ingress_id_109 : _GEN_4589; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4591 = 7'h6e == out_payload_rob_idx[6:0] ? rob_ingress_id_110 : _GEN_4590; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4592 = 7'h6f == out_payload_rob_idx[6:0] ? rob_ingress_id_111 : _GEN_4591; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4593 = 7'h70 == out_payload_rob_idx[6:0] ? rob_ingress_id_112 : _GEN_4592; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4594 = 7'h71 == out_payload_rob_idx[6:0] ? rob_ingress_id_113 : _GEN_4593; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4595 = 7'h72 == out_payload_rob_idx[6:0] ? rob_ingress_id_114 : _GEN_4594; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4596 = 7'h73 == out_payload_rob_idx[6:0] ? rob_ingress_id_115 : _GEN_4595; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4597 = 7'h74 == out_payload_rob_idx[6:0] ? rob_ingress_id_116 : _GEN_4596; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4598 = 7'h75 == out_payload_rob_idx[6:0] ? rob_ingress_id_117 : _GEN_4597; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4599 = 7'h76 == out_payload_rob_idx[6:0] ? rob_ingress_id_118 : _GEN_4598; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4600 = 7'h77 == out_payload_rob_idx[6:0] ? rob_ingress_id_119 : _GEN_4599; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4601 = 7'h78 == out_payload_rob_idx[6:0] ? rob_ingress_id_120 : _GEN_4600; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4602 = 7'h79 == out_payload_rob_idx[6:0] ? rob_ingress_id_121 : _GEN_4601; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4603 = 7'h7a == out_payload_rob_idx[6:0] ? rob_ingress_id_122 : _GEN_4602; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4604 = 7'h7b == out_payload_rob_idx[6:0] ? rob_ingress_id_123 : _GEN_4603; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4605 = 7'h7c == out_payload_rob_idx[6:0] ? rob_ingress_id_124 : _GEN_4604; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4606 = 7'h7d == out_payload_rob_idx[6:0] ? rob_ingress_id_125 : _GEN_4605; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4607 = 7'h7e == out_payload_rob_idx[6:0] ? rob_ingress_id_126 : _GEN_4606; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4608 = 7'h7f == out_payload_rob_idx[6:0] ? rob_ingress_id_127 : _GEN_4607; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_4610 = 7'h1 == out_payload_rob_idx[6:0] ? rob_egress_id_1 : rob_egress_id_0; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4611 = 7'h2 == out_payload_rob_idx[6:0] ? rob_egress_id_2 : _GEN_4610; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4612 = 7'h3 == out_payload_rob_idx[6:0] ? rob_egress_id_3 : _GEN_4611; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4613 = 7'h4 == out_payload_rob_idx[6:0] ? rob_egress_id_4 : _GEN_4612; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4614 = 7'h5 == out_payload_rob_idx[6:0] ? rob_egress_id_5 : _GEN_4613; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4615 = 7'h6 == out_payload_rob_idx[6:0] ? rob_egress_id_6 : _GEN_4614; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4616 = 7'h7 == out_payload_rob_idx[6:0] ? rob_egress_id_7 : _GEN_4615; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4617 = 7'h8 == out_payload_rob_idx[6:0] ? rob_egress_id_8 : _GEN_4616; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4618 = 7'h9 == out_payload_rob_idx[6:0] ? rob_egress_id_9 : _GEN_4617; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4619 = 7'ha == out_payload_rob_idx[6:0] ? rob_egress_id_10 : _GEN_4618; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4620 = 7'hb == out_payload_rob_idx[6:0] ? rob_egress_id_11 : _GEN_4619; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4621 = 7'hc == out_payload_rob_idx[6:0] ? rob_egress_id_12 : _GEN_4620; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4622 = 7'hd == out_payload_rob_idx[6:0] ? rob_egress_id_13 : _GEN_4621; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4623 = 7'he == out_payload_rob_idx[6:0] ? rob_egress_id_14 : _GEN_4622; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4624 = 7'hf == out_payload_rob_idx[6:0] ? rob_egress_id_15 : _GEN_4623; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4625 = 7'h10 == out_payload_rob_idx[6:0] ? rob_egress_id_16 : _GEN_4624; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4626 = 7'h11 == out_payload_rob_idx[6:0] ? rob_egress_id_17 : _GEN_4625; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4627 = 7'h12 == out_payload_rob_idx[6:0] ? rob_egress_id_18 : _GEN_4626; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4628 = 7'h13 == out_payload_rob_idx[6:0] ? rob_egress_id_19 : _GEN_4627; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4629 = 7'h14 == out_payload_rob_idx[6:0] ? rob_egress_id_20 : _GEN_4628; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4630 = 7'h15 == out_payload_rob_idx[6:0] ? rob_egress_id_21 : _GEN_4629; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4631 = 7'h16 == out_payload_rob_idx[6:0] ? rob_egress_id_22 : _GEN_4630; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4632 = 7'h17 == out_payload_rob_idx[6:0] ? rob_egress_id_23 : _GEN_4631; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4633 = 7'h18 == out_payload_rob_idx[6:0] ? rob_egress_id_24 : _GEN_4632; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4634 = 7'h19 == out_payload_rob_idx[6:0] ? rob_egress_id_25 : _GEN_4633; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4635 = 7'h1a == out_payload_rob_idx[6:0] ? rob_egress_id_26 : _GEN_4634; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4636 = 7'h1b == out_payload_rob_idx[6:0] ? rob_egress_id_27 : _GEN_4635; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4637 = 7'h1c == out_payload_rob_idx[6:0] ? rob_egress_id_28 : _GEN_4636; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4638 = 7'h1d == out_payload_rob_idx[6:0] ? rob_egress_id_29 : _GEN_4637; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4639 = 7'h1e == out_payload_rob_idx[6:0] ? rob_egress_id_30 : _GEN_4638; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4640 = 7'h1f == out_payload_rob_idx[6:0] ? rob_egress_id_31 : _GEN_4639; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4641 = 7'h20 == out_payload_rob_idx[6:0] ? rob_egress_id_32 : _GEN_4640; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4642 = 7'h21 == out_payload_rob_idx[6:0] ? rob_egress_id_33 : _GEN_4641; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4643 = 7'h22 == out_payload_rob_idx[6:0] ? rob_egress_id_34 : _GEN_4642; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4644 = 7'h23 == out_payload_rob_idx[6:0] ? rob_egress_id_35 : _GEN_4643; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4645 = 7'h24 == out_payload_rob_idx[6:0] ? rob_egress_id_36 : _GEN_4644; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4646 = 7'h25 == out_payload_rob_idx[6:0] ? rob_egress_id_37 : _GEN_4645; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4647 = 7'h26 == out_payload_rob_idx[6:0] ? rob_egress_id_38 : _GEN_4646; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4648 = 7'h27 == out_payload_rob_idx[6:0] ? rob_egress_id_39 : _GEN_4647; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4649 = 7'h28 == out_payload_rob_idx[6:0] ? rob_egress_id_40 : _GEN_4648; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4650 = 7'h29 == out_payload_rob_idx[6:0] ? rob_egress_id_41 : _GEN_4649; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4651 = 7'h2a == out_payload_rob_idx[6:0] ? rob_egress_id_42 : _GEN_4650; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4652 = 7'h2b == out_payload_rob_idx[6:0] ? rob_egress_id_43 : _GEN_4651; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4653 = 7'h2c == out_payload_rob_idx[6:0] ? rob_egress_id_44 : _GEN_4652; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4654 = 7'h2d == out_payload_rob_idx[6:0] ? rob_egress_id_45 : _GEN_4653; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4655 = 7'h2e == out_payload_rob_idx[6:0] ? rob_egress_id_46 : _GEN_4654; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4656 = 7'h2f == out_payload_rob_idx[6:0] ? rob_egress_id_47 : _GEN_4655; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4657 = 7'h30 == out_payload_rob_idx[6:0] ? rob_egress_id_48 : _GEN_4656; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4658 = 7'h31 == out_payload_rob_idx[6:0] ? rob_egress_id_49 : _GEN_4657; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4659 = 7'h32 == out_payload_rob_idx[6:0] ? rob_egress_id_50 : _GEN_4658; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4660 = 7'h33 == out_payload_rob_idx[6:0] ? rob_egress_id_51 : _GEN_4659; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4661 = 7'h34 == out_payload_rob_idx[6:0] ? rob_egress_id_52 : _GEN_4660; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4662 = 7'h35 == out_payload_rob_idx[6:0] ? rob_egress_id_53 : _GEN_4661; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4663 = 7'h36 == out_payload_rob_idx[6:0] ? rob_egress_id_54 : _GEN_4662; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4664 = 7'h37 == out_payload_rob_idx[6:0] ? rob_egress_id_55 : _GEN_4663; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4665 = 7'h38 == out_payload_rob_idx[6:0] ? rob_egress_id_56 : _GEN_4664; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4666 = 7'h39 == out_payload_rob_idx[6:0] ? rob_egress_id_57 : _GEN_4665; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4667 = 7'h3a == out_payload_rob_idx[6:0] ? rob_egress_id_58 : _GEN_4666; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4668 = 7'h3b == out_payload_rob_idx[6:0] ? rob_egress_id_59 : _GEN_4667; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4669 = 7'h3c == out_payload_rob_idx[6:0] ? rob_egress_id_60 : _GEN_4668; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4670 = 7'h3d == out_payload_rob_idx[6:0] ? rob_egress_id_61 : _GEN_4669; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4671 = 7'h3e == out_payload_rob_idx[6:0] ? rob_egress_id_62 : _GEN_4670; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4672 = 7'h3f == out_payload_rob_idx[6:0] ? rob_egress_id_63 : _GEN_4671; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4673 = 7'h40 == out_payload_rob_idx[6:0] ? rob_egress_id_64 : _GEN_4672; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4674 = 7'h41 == out_payload_rob_idx[6:0] ? rob_egress_id_65 : _GEN_4673; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4675 = 7'h42 == out_payload_rob_idx[6:0] ? rob_egress_id_66 : _GEN_4674; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4676 = 7'h43 == out_payload_rob_idx[6:0] ? rob_egress_id_67 : _GEN_4675; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4677 = 7'h44 == out_payload_rob_idx[6:0] ? rob_egress_id_68 : _GEN_4676; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4678 = 7'h45 == out_payload_rob_idx[6:0] ? rob_egress_id_69 : _GEN_4677; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4679 = 7'h46 == out_payload_rob_idx[6:0] ? rob_egress_id_70 : _GEN_4678; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4680 = 7'h47 == out_payload_rob_idx[6:0] ? rob_egress_id_71 : _GEN_4679; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4681 = 7'h48 == out_payload_rob_idx[6:0] ? rob_egress_id_72 : _GEN_4680; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4682 = 7'h49 == out_payload_rob_idx[6:0] ? rob_egress_id_73 : _GEN_4681; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4683 = 7'h4a == out_payload_rob_idx[6:0] ? rob_egress_id_74 : _GEN_4682; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4684 = 7'h4b == out_payload_rob_idx[6:0] ? rob_egress_id_75 : _GEN_4683; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4685 = 7'h4c == out_payload_rob_idx[6:0] ? rob_egress_id_76 : _GEN_4684; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4686 = 7'h4d == out_payload_rob_idx[6:0] ? rob_egress_id_77 : _GEN_4685; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4687 = 7'h4e == out_payload_rob_idx[6:0] ? rob_egress_id_78 : _GEN_4686; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4688 = 7'h4f == out_payload_rob_idx[6:0] ? rob_egress_id_79 : _GEN_4687; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4689 = 7'h50 == out_payload_rob_idx[6:0] ? rob_egress_id_80 : _GEN_4688; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4690 = 7'h51 == out_payload_rob_idx[6:0] ? rob_egress_id_81 : _GEN_4689; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4691 = 7'h52 == out_payload_rob_idx[6:0] ? rob_egress_id_82 : _GEN_4690; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4692 = 7'h53 == out_payload_rob_idx[6:0] ? rob_egress_id_83 : _GEN_4691; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4693 = 7'h54 == out_payload_rob_idx[6:0] ? rob_egress_id_84 : _GEN_4692; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4694 = 7'h55 == out_payload_rob_idx[6:0] ? rob_egress_id_85 : _GEN_4693; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4695 = 7'h56 == out_payload_rob_idx[6:0] ? rob_egress_id_86 : _GEN_4694; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4696 = 7'h57 == out_payload_rob_idx[6:0] ? rob_egress_id_87 : _GEN_4695; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4697 = 7'h58 == out_payload_rob_idx[6:0] ? rob_egress_id_88 : _GEN_4696; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4698 = 7'h59 == out_payload_rob_idx[6:0] ? rob_egress_id_89 : _GEN_4697; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4699 = 7'h5a == out_payload_rob_idx[6:0] ? rob_egress_id_90 : _GEN_4698; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4700 = 7'h5b == out_payload_rob_idx[6:0] ? rob_egress_id_91 : _GEN_4699; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4701 = 7'h5c == out_payload_rob_idx[6:0] ? rob_egress_id_92 : _GEN_4700; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4702 = 7'h5d == out_payload_rob_idx[6:0] ? rob_egress_id_93 : _GEN_4701; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4703 = 7'h5e == out_payload_rob_idx[6:0] ? rob_egress_id_94 : _GEN_4702; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4704 = 7'h5f == out_payload_rob_idx[6:0] ? rob_egress_id_95 : _GEN_4703; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4705 = 7'h60 == out_payload_rob_idx[6:0] ? rob_egress_id_96 : _GEN_4704; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4706 = 7'h61 == out_payload_rob_idx[6:0] ? rob_egress_id_97 : _GEN_4705; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4707 = 7'h62 == out_payload_rob_idx[6:0] ? rob_egress_id_98 : _GEN_4706; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4708 = 7'h63 == out_payload_rob_idx[6:0] ? rob_egress_id_99 : _GEN_4707; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4709 = 7'h64 == out_payload_rob_idx[6:0] ? rob_egress_id_100 : _GEN_4708; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4710 = 7'h65 == out_payload_rob_idx[6:0] ? rob_egress_id_101 : _GEN_4709; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4711 = 7'h66 == out_payload_rob_idx[6:0] ? rob_egress_id_102 : _GEN_4710; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4712 = 7'h67 == out_payload_rob_idx[6:0] ? rob_egress_id_103 : _GEN_4711; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4713 = 7'h68 == out_payload_rob_idx[6:0] ? rob_egress_id_104 : _GEN_4712; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4714 = 7'h69 == out_payload_rob_idx[6:0] ? rob_egress_id_105 : _GEN_4713; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4715 = 7'h6a == out_payload_rob_idx[6:0] ? rob_egress_id_106 : _GEN_4714; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4716 = 7'h6b == out_payload_rob_idx[6:0] ? rob_egress_id_107 : _GEN_4715; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4717 = 7'h6c == out_payload_rob_idx[6:0] ? rob_egress_id_108 : _GEN_4716; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4718 = 7'h6d == out_payload_rob_idx[6:0] ? rob_egress_id_109 : _GEN_4717; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4719 = 7'h6e == out_payload_rob_idx[6:0] ? rob_egress_id_110 : _GEN_4718; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4720 = 7'h6f == out_payload_rob_idx[6:0] ? rob_egress_id_111 : _GEN_4719; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4721 = 7'h70 == out_payload_rob_idx[6:0] ? rob_egress_id_112 : _GEN_4720; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4722 = 7'h71 == out_payload_rob_idx[6:0] ? rob_egress_id_113 : _GEN_4721; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4723 = 7'h72 == out_payload_rob_idx[6:0] ? rob_egress_id_114 : _GEN_4722; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4724 = 7'h73 == out_payload_rob_idx[6:0] ? rob_egress_id_115 : _GEN_4723; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4725 = 7'h74 == out_payload_rob_idx[6:0] ? rob_egress_id_116 : _GEN_4724; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4726 = 7'h75 == out_payload_rob_idx[6:0] ? rob_egress_id_117 : _GEN_4725; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4727 = 7'h76 == out_payload_rob_idx[6:0] ? rob_egress_id_118 : _GEN_4726; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4728 = 7'h77 == out_payload_rob_idx[6:0] ? rob_egress_id_119 : _GEN_4727; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4729 = 7'h78 == out_payload_rob_idx[6:0] ? rob_egress_id_120 : _GEN_4728; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4730 = 7'h79 == out_payload_rob_idx[6:0] ? rob_egress_id_121 : _GEN_4729; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4731 = 7'h7a == out_payload_rob_idx[6:0] ? rob_egress_id_122 : _GEN_4730; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4732 = 7'h7b == out_payload_rob_idx[6:0] ? rob_egress_id_123 : _GEN_4731; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4733 = 7'h7c == out_payload_rob_idx[6:0] ? rob_egress_id_124 : _GEN_4732; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4734 = 7'h7d == out_payload_rob_idx[6:0] ? rob_egress_id_125 : _GEN_4733; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4735 = 7'h7e == out_payload_rob_idx[6:0] ? rob_egress_id_126 : _GEN_4734; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_4736 = 7'h7f == out_payload_rob_idx[6:0] ? rob_egress_id_127 : _GEN_4735; // @[TestHarness.scala 204:{18,18}]
  wire [3:0] _GEN_4738 = 7'h1 == out_payload_rob_idx[6:0] ? rob_flits_returned_1 : rob_flits_returned_0; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4739 = 7'h2 == out_payload_rob_idx[6:0] ? rob_flits_returned_2 : _GEN_4738; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4740 = 7'h3 == out_payload_rob_idx[6:0] ? rob_flits_returned_3 : _GEN_4739; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4741 = 7'h4 == out_payload_rob_idx[6:0] ? rob_flits_returned_4 : _GEN_4740; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4742 = 7'h5 == out_payload_rob_idx[6:0] ? rob_flits_returned_5 : _GEN_4741; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4743 = 7'h6 == out_payload_rob_idx[6:0] ? rob_flits_returned_6 : _GEN_4742; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4744 = 7'h7 == out_payload_rob_idx[6:0] ? rob_flits_returned_7 : _GEN_4743; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4745 = 7'h8 == out_payload_rob_idx[6:0] ? rob_flits_returned_8 : _GEN_4744; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4746 = 7'h9 == out_payload_rob_idx[6:0] ? rob_flits_returned_9 : _GEN_4745; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4747 = 7'ha == out_payload_rob_idx[6:0] ? rob_flits_returned_10 : _GEN_4746; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4748 = 7'hb == out_payload_rob_idx[6:0] ? rob_flits_returned_11 : _GEN_4747; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4749 = 7'hc == out_payload_rob_idx[6:0] ? rob_flits_returned_12 : _GEN_4748; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4750 = 7'hd == out_payload_rob_idx[6:0] ? rob_flits_returned_13 : _GEN_4749; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4751 = 7'he == out_payload_rob_idx[6:0] ? rob_flits_returned_14 : _GEN_4750; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4752 = 7'hf == out_payload_rob_idx[6:0] ? rob_flits_returned_15 : _GEN_4751; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4753 = 7'h10 == out_payload_rob_idx[6:0] ? rob_flits_returned_16 : _GEN_4752; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4754 = 7'h11 == out_payload_rob_idx[6:0] ? rob_flits_returned_17 : _GEN_4753; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4755 = 7'h12 == out_payload_rob_idx[6:0] ? rob_flits_returned_18 : _GEN_4754; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4756 = 7'h13 == out_payload_rob_idx[6:0] ? rob_flits_returned_19 : _GEN_4755; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4757 = 7'h14 == out_payload_rob_idx[6:0] ? rob_flits_returned_20 : _GEN_4756; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4758 = 7'h15 == out_payload_rob_idx[6:0] ? rob_flits_returned_21 : _GEN_4757; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4759 = 7'h16 == out_payload_rob_idx[6:0] ? rob_flits_returned_22 : _GEN_4758; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4760 = 7'h17 == out_payload_rob_idx[6:0] ? rob_flits_returned_23 : _GEN_4759; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4761 = 7'h18 == out_payload_rob_idx[6:0] ? rob_flits_returned_24 : _GEN_4760; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4762 = 7'h19 == out_payload_rob_idx[6:0] ? rob_flits_returned_25 : _GEN_4761; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4763 = 7'h1a == out_payload_rob_idx[6:0] ? rob_flits_returned_26 : _GEN_4762; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4764 = 7'h1b == out_payload_rob_idx[6:0] ? rob_flits_returned_27 : _GEN_4763; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4765 = 7'h1c == out_payload_rob_idx[6:0] ? rob_flits_returned_28 : _GEN_4764; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4766 = 7'h1d == out_payload_rob_idx[6:0] ? rob_flits_returned_29 : _GEN_4765; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4767 = 7'h1e == out_payload_rob_idx[6:0] ? rob_flits_returned_30 : _GEN_4766; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4768 = 7'h1f == out_payload_rob_idx[6:0] ? rob_flits_returned_31 : _GEN_4767; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4769 = 7'h20 == out_payload_rob_idx[6:0] ? rob_flits_returned_32 : _GEN_4768; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4770 = 7'h21 == out_payload_rob_idx[6:0] ? rob_flits_returned_33 : _GEN_4769; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4771 = 7'h22 == out_payload_rob_idx[6:0] ? rob_flits_returned_34 : _GEN_4770; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4772 = 7'h23 == out_payload_rob_idx[6:0] ? rob_flits_returned_35 : _GEN_4771; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4773 = 7'h24 == out_payload_rob_idx[6:0] ? rob_flits_returned_36 : _GEN_4772; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4774 = 7'h25 == out_payload_rob_idx[6:0] ? rob_flits_returned_37 : _GEN_4773; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4775 = 7'h26 == out_payload_rob_idx[6:0] ? rob_flits_returned_38 : _GEN_4774; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4776 = 7'h27 == out_payload_rob_idx[6:0] ? rob_flits_returned_39 : _GEN_4775; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4777 = 7'h28 == out_payload_rob_idx[6:0] ? rob_flits_returned_40 : _GEN_4776; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4778 = 7'h29 == out_payload_rob_idx[6:0] ? rob_flits_returned_41 : _GEN_4777; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4779 = 7'h2a == out_payload_rob_idx[6:0] ? rob_flits_returned_42 : _GEN_4778; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4780 = 7'h2b == out_payload_rob_idx[6:0] ? rob_flits_returned_43 : _GEN_4779; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4781 = 7'h2c == out_payload_rob_idx[6:0] ? rob_flits_returned_44 : _GEN_4780; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4782 = 7'h2d == out_payload_rob_idx[6:0] ? rob_flits_returned_45 : _GEN_4781; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4783 = 7'h2e == out_payload_rob_idx[6:0] ? rob_flits_returned_46 : _GEN_4782; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4784 = 7'h2f == out_payload_rob_idx[6:0] ? rob_flits_returned_47 : _GEN_4783; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4785 = 7'h30 == out_payload_rob_idx[6:0] ? rob_flits_returned_48 : _GEN_4784; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4786 = 7'h31 == out_payload_rob_idx[6:0] ? rob_flits_returned_49 : _GEN_4785; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4787 = 7'h32 == out_payload_rob_idx[6:0] ? rob_flits_returned_50 : _GEN_4786; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4788 = 7'h33 == out_payload_rob_idx[6:0] ? rob_flits_returned_51 : _GEN_4787; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4789 = 7'h34 == out_payload_rob_idx[6:0] ? rob_flits_returned_52 : _GEN_4788; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4790 = 7'h35 == out_payload_rob_idx[6:0] ? rob_flits_returned_53 : _GEN_4789; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4791 = 7'h36 == out_payload_rob_idx[6:0] ? rob_flits_returned_54 : _GEN_4790; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4792 = 7'h37 == out_payload_rob_idx[6:0] ? rob_flits_returned_55 : _GEN_4791; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4793 = 7'h38 == out_payload_rob_idx[6:0] ? rob_flits_returned_56 : _GEN_4792; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4794 = 7'h39 == out_payload_rob_idx[6:0] ? rob_flits_returned_57 : _GEN_4793; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4795 = 7'h3a == out_payload_rob_idx[6:0] ? rob_flits_returned_58 : _GEN_4794; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4796 = 7'h3b == out_payload_rob_idx[6:0] ? rob_flits_returned_59 : _GEN_4795; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4797 = 7'h3c == out_payload_rob_idx[6:0] ? rob_flits_returned_60 : _GEN_4796; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4798 = 7'h3d == out_payload_rob_idx[6:0] ? rob_flits_returned_61 : _GEN_4797; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4799 = 7'h3e == out_payload_rob_idx[6:0] ? rob_flits_returned_62 : _GEN_4798; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4800 = 7'h3f == out_payload_rob_idx[6:0] ? rob_flits_returned_63 : _GEN_4799; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4801 = 7'h40 == out_payload_rob_idx[6:0] ? rob_flits_returned_64 : _GEN_4800; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4802 = 7'h41 == out_payload_rob_idx[6:0] ? rob_flits_returned_65 : _GEN_4801; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4803 = 7'h42 == out_payload_rob_idx[6:0] ? rob_flits_returned_66 : _GEN_4802; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4804 = 7'h43 == out_payload_rob_idx[6:0] ? rob_flits_returned_67 : _GEN_4803; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4805 = 7'h44 == out_payload_rob_idx[6:0] ? rob_flits_returned_68 : _GEN_4804; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4806 = 7'h45 == out_payload_rob_idx[6:0] ? rob_flits_returned_69 : _GEN_4805; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4807 = 7'h46 == out_payload_rob_idx[6:0] ? rob_flits_returned_70 : _GEN_4806; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4808 = 7'h47 == out_payload_rob_idx[6:0] ? rob_flits_returned_71 : _GEN_4807; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4809 = 7'h48 == out_payload_rob_idx[6:0] ? rob_flits_returned_72 : _GEN_4808; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4810 = 7'h49 == out_payload_rob_idx[6:0] ? rob_flits_returned_73 : _GEN_4809; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4811 = 7'h4a == out_payload_rob_idx[6:0] ? rob_flits_returned_74 : _GEN_4810; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4812 = 7'h4b == out_payload_rob_idx[6:0] ? rob_flits_returned_75 : _GEN_4811; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4813 = 7'h4c == out_payload_rob_idx[6:0] ? rob_flits_returned_76 : _GEN_4812; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4814 = 7'h4d == out_payload_rob_idx[6:0] ? rob_flits_returned_77 : _GEN_4813; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4815 = 7'h4e == out_payload_rob_idx[6:0] ? rob_flits_returned_78 : _GEN_4814; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4816 = 7'h4f == out_payload_rob_idx[6:0] ? rob_flits_returned_79 : _GEN_4815; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4817 = 7'h50 == out_payload_rob_idx[6:0] ? rob_flits_returned_80 : _GEN_4816; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4818 = 7'h51 == out_payload_rob_idx[6:0] ? rob_flits_returned_81 : _GEN_4817; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4819 = 7'h52 == out_payload_rob_idx[6:0] ? rob_flits_returned_82 : _GEN_4818; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4820 = 7'h53 == out_payload_rob_idx[6:0] ? rob_flits_returned_83 : _GEN_4819; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4821 = 7'h54 == out_payload_rob_idx[6:0] ? rob_flits_returned_84 : _GEN_4820; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4822 = 7'h55 == out_payload_rob_idx[6:0] ? rob_flits_returned_85 : _GEN_4821; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4823 = 7'h56 == out_payload_rob_idx[6:0] ? rob_flits_returned_86 : _GEN_4822; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4824 = 7'h57 == out_payload_rob_idx[6:0] ? rob_flits_returned_87 : _GEN_4823; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4825 = 7'h58 == out_payload_rob_idx[6:0] ? rob_flits_returned_88 : _GEN_4824; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4826 = 7'h59 == out_payload_rob_idx[6:0] ? rob_flits_returned_89 : _GEN_4825; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4827 = 7'h5a == out_payload_rob_idx[6:0] ? rob_flits_returned_90 : _GEN_4826; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4828 = 7'h5b == out_payload_rob_idx[6:0] ? rob_flits_returned_91 : _GEN_4827; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4829 = 7'h5c == out_payload_rob_idx[6:0] ? rob_flits_returned_92 : _GEN_4828; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4830 = 7'h5d == out_payload_rob_idx[6:0] ? rob_flits_returned_93 : _GEN_4829; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4831 = 7'h5e == out_payload_rob_idx[6:0] ? rob_flits_returned_94 : _GEN_4830; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4832 = 7'h5f == out_payload_rob_idx[6:0] ? rob_flits_returned_95 : _GEN_4831; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4833 = 7'h60 == out_payload_rob_idx[6:0] ? rob_flits_returned_96 : _GEN_4832; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4834 = 7'h61 == out_payload_rob_idx[6:0] ? rob_flits_returned_97 : _GEN_4833; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4835 = 7'h62 == out_payload_rob_idx[6:0] ? rob_flits_returned_98 : _GEN_4834; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4836 = 7'h63 == out_payload_rob_idx[6:0] ? rob_flits_returned_99 : _GEN_4835; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4837 = 7'h64 == out_payload_rob_idx[6:0] ? rob_flits_returned_100 : _GEN_4836; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4838 = 7'h65 == out_payload_rob_idx[6:0] ? rob_flits_returned_101 : _GEN_4837; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4839 = 7'h66 == out_payload_rob_idx[6:0] ? rob_flits_returned_102 : _GEN_4838; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4840 = 7'h67 == out_payload_rob_idx[6:0] ? rob_flits_returned_103 : _GEN_4839; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4841 = 7'h68 == out_payload_rob_idx[6:0] ? rob_flits_returned_104 : _GEN_4840; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4842 = 7'h69 == out_payload_rob_idx[6:0] ? rob_flits_returned_105 : _GEN_4841; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4843 = 7'h6a == out_payload_rob_idx[6:0] ? rob_flits_returned_106 : _GEN_4842; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4844 = 7'h6b == out_payload_rob_idx[6:0] ? rob_flits_returned_107 : _GEN_4843; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4845 = 7'h6c == out_payload_rob_idx[6:0] ? rob_flits_returned_108 : _GEN_4844; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4846 = 7'h6d == out_payload_rob_idx[6:0] ? rob_flits_returned_109 : _GEN_4845; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4847 = 7'h6e == out_payload_rob_idx[6:0] ? rob_flits_returned_110 : _GEN_4846; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4848 = 7'h6f == out_payload_rob_idx[6:0] ? rob_flits_returned_111 : _GEN_4847; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4849 = 7'h70 == out_payload_rob_idx[6:0] ? rob_flits_returned_112 : _GEN_4848; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4850 = 7'h71 == out_payload_rob_idx[6:0] ? rob_flits_returned_113 : _GEN_4849; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4851 = 7'h72 == out_payload_rob_idx[6:0] ? rob_flits_returned_114 : _GEN_4850; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4852 = 7'h73 == out_payload_rob_idx[6:0] ? rob_flits_returned_115 : _GEN_4851; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4853 = 7'h74 == out_payload_rob_idx[6:0] ? rob_flits_returned_116 : _GEN_4852; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4854 = 7'h75 == out_payload_rob_idx[6:0] ? rob_flits_returned_117 : _GEN_4853; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4855 = 7'h76 == out_payload_rob_idx[6:0] ? rob_flits_returned_118 : _GEN_4854; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4856 = 7'h77 == out_payload_rob_idx[6:0] ? rob_flits_returned_119 : _GEN_4855; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4857 = 7'h78 == out_payload_rob_idx[6:0] ? rob_flits_returned_120 : _GEN_4856; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4858 = 7'h79 == out_payload_rob_idx[6:0] ? rob_flits_returned_121 : _GEN_4857; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4859 = 7'h7a == out_payload_rob_idx[6:0] ? rob_flits_returned_122 : _GEN_4858; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4860 = 7'h7b == out_payload_rob_idx[6:0] ? rob_flits_returned_123 : _GEN_4859; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4861 = 7'h7c == out_payload_rob_idx[6:0] ? rob_flits_returned_124 : _GEN_4860; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4862 = 7'h7d == out_payload_rob_idx[6:0] ? rob_flits_returned_125 : _GEN_4861; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4863 = 7'h7e == out_payload_rob_idx[6:0] ? rob_flits_returned_126 : _GEN_4862; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4864 = 7'h7f == out_payload_rob_idx[6:0] ? rob_flits_returned_127 : _GEN_4863; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4866 = 7'h1 == out_payload_rob_idx[6:0] ? rob_n_flits_1 : rob_n_flits_0; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4867 = 7'h2 == out_payload_rob_idx[6:0] ? rob_n_flits_2 : _GEN_4866; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4868 = 7'h3 == out_payload_rob_idx[6:0] ? rob_n_flits_3 : _GEN_4867; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4869 = 7'h4 == out_payload_rob_idx[6:0] ? rob_n_flits_4 : _GEN_4868; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4870 = 7'h5 == out_payload_rob_idx[6:0] ? rob_n_flits_5 : _GEN_4869; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4871 = 7'h6 == out_payload_rob_idx[6:0] ? rob_n_flits_6 : _GEN_4870; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4872 = 7'h7 == out_payload_rob_idx[6:0] ? rob_n_flits_7 : _GEN_4871; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4873 = 7'h8 == out_payload_rob_idx[6:0] ? rob_n_flits_8 : _GEN_4872; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4874 = 7'h9 == out_payload_rob_idx[6:0] ? rob_n_flits_9 : _GEN_4873; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4875 = 7'ha == out_payload_rob_idx[6:0] ? rob_n_flits_10 : _GEN_4874; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4876 = 7'hb == out_payload_rob_idx[6:0] ? rob_n_flits_11 : _GEN_4875; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4877 = 7'hc == out_payload_rob_idx[6:0] ? rob_n_flits_12 : _GEN_4876; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4878 = 7'hd == out_payload_rob_idx[6:0] ? rob_n_flits_13 : _GEN_4877; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4879 = 7'he == out_payload_rob_idx[6:0] ? rob_n_flits_14 : _GEN_4878; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4880 = 7'hf == out_payload_rob_idx[6:0] ? rob_n_flits_15 : _GEN_4879; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4881 = 7'h10 == out_payload_rob_idx[6:0] ? rob_n_flits_16 : _GEN_4880; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4882 = 7'h11 == out_payload_rob_idx[6:0] ? rob_n_flits_17 : _GEN_4881; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4883 = 7'h12 == out_payload_rob_idx[6:0] ? rob_n_flits_18 : _GEN_4882; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4884 = 7'h13 == out_payload_rob_idx[6:0] ? rob_n_flits_19 : _GEN_4883; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4885 = 7'h14 == out_payload_rob_idx[6:0] ? rob_n_flits_20 : _GEN_4884; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4886 = 7'h15 == out_payload_rob_idx[6:0] ? rob_n_flits_21 : _GEN_4885; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4887 = 7'h16 == out_payload_rob_idx[6:0] ? rob_n_flits_22 : _GEN_4886; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4888 = 7'h17 == out_payload_rob_idx[6:0] ? rob_n_flits_23 : _GEN_4887; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4889 = 7'h18 == out_payload_rob_idx[6:0] ? rob_n_flits_24 : _GEN_4888; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4890 = 7'h19 == out_payload_rob_idx[6:0] ? rob_n_flits_25 : _GEN_4889; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4891 = 7'h1a == out_payload_rob_idx[6:0] ? rob_n_flits_26 : _GEN_4890; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4892 = 7'h1b == out_payload_rob_idx[6:0] ? rob_n_flits_27 : _GEN_4891; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4893 = 7'h1c == out_payload_rob_idx[6:0] ? rob_n_flits_28 : _GEN_4892; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4894 = 7'h1d == out_payload_rob_idx[6:0] ? rob_n_flits_29 : _GEN_4893; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4895 = 7'h1e == out_payload_rob_idx[6:0] ? rob_n_flits_30 : _GEN_4894; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4896 = 7'h1f == out_payload_rob_idx[6:0] ? rob_n_flits_31 : _GEN_4895; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4897 = 7'h20 == out_payload_rob_idx[6:0] ? rob_n_flits_32 : _GEN_4896; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4898 = 7'h21 == out_payload_rob_idx[6:0] ? rob_n_flits_33 : _GEN_4897; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4899 = 7'h22 == out_payload_rob_idx[6:0] ? rob_n_flits_34 : _GEN_4898; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4900 = 7'h23 == out_payload_rob_idx[6:0] ? rob_n_flits_35 : _GEN_4899; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4901 = 7'h24 == out_payload_rob_idx[6:0] ? rob_n_flits_36 : _GEN_4900; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4902 = 7'h25 == out_payload_rob_idx[6:0] ? rob_n_flits_37 : _GEN_4901; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4903 = 7'h26 == out_payload_rob_idx[6:0] ? rob_n_flits_38 : _GEN_4902; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4904 = 7'h27 == out_payload_rob_idx[6:0] ? rob_n_flits_39 : _GEN_4903; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4905 = 7'h28 == out_payload_rob_idx[6:0] ? rob_n_flits_40 : _GEN_4904; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4906 = 7'h29 == out_payload_rob_idx[6:0] ? rob_n_flits_41 : _GEN_4905; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4907 = 7'h2a == out_payload_rob_idx[6:0] ? rob_n_flits_42 : _GEN_4906; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4908 = 7'h2b == out_payload_rob_idx[6:0] ? rob_n_flits_43 : _GEN_4907; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4909 = 7'h2c == out_payload_rob_idx[6:0] ? rob_n_flits_44 : _GEN_4908; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4910 = 7'h2d == out_payload_rob_idx[6:0] ? rob_n_flits_45 : _GEN_4909; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4911 = 7'h2e == out_payload_rob_idx[6:0] ? rob_n_flits_46 : _GEN_4910; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4912 = 7'h2f == out_payload_rob_idx[6:0] ? rob_n_flits_47 : _GEN_4911; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4913 = 7'h30 == out_payload_rob_idx[6:0] ? rob_n_flits_48 : _GEN_4912; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4914 = 7'h31 == out_payload_rob_idx[6:0] ? rob_n_flits_49 : _GEN_4913; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4915 = 7'h32 == out_payload_rob_idx[6:0] ? rob_n_flits_50 : _GEN_4914; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4916 = 7'h33 == out_payload_rob_idx[6:0] ? rob_n_flits_51 : _GEN_4915; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4917 = 7'h34 == out_payload_rob_idx[6:0] ? rob_n_flits_52 : _GEN_4916; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4918 = 7'h35 == out_payload_rob_idx[6:0] ? rob_n_flits_53 : _GEN_4917; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4919 = 7'h36 == out_payload_rob_idx[6:0] ? rob_n_flits_54 : _GEN_4918; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4920 = 7'h37 == out_payload_rob_idx[6:0] ? rob_n_flits_55 : _GEN_4919; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4921 = 7'h38 == out_payload_rob_idx[6:0] ? rob_n_flits_56 : _GEN_4920; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4922 = 7'h39 == out_payload_rob_idx[6:0] ? rob_n_flits_57 : _GEN_4921; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4923 = 7'h3a == out_payload_rob_idx[6:0] ? rob_n_flits_58 : _GEN_4922; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4924 = 7'h3b == out_payload_rob_idx[6:0] ? rob_n_flits_59 : _GEN_4923; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4925 = 7'h3c == out_payload_rob_idx[6:0] ? rob_n_flits_60 : _GEN_4924; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4926 = 7'h3d == out_payload_rob_idx[6:0] ? rob_n_flits_61 : _GEN_4925; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4927 = 7'h3e == out_payload_rob_idx[6:0] ? rob_n_flits_62 : _GEN_4926; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4928 = 7'h3f == out_payload_rob_idx[6:0] ? rob_n_flits_63 : _GEN_4927; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4929 = 7'h40 == out_payload_rob_idx[6:0] ? rob_n_flits_64 : _GEN_4928; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4930 = 7'h41 == out_payload_rob_idx[6:0] ? rob_n_flits_65 : _GEN_4929; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4931 = 7'h42 == out_payload_rob_idx[6:0] ? rob_n_flits_66 : _GEN_4930; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4932 = 7'h43 == out_payload_rob_idx[6:0] ? rob_n_flits_67 : _GEN_4931; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4933 = 7'h44 == out_payload_rob_idx[6:0] ? rob_n_flits_68 : _GEN_4932; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4934 = 7'h45 == out_payload_rob_idx[6:0] ? rob_n_flits_69 : _GEN_4933; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4935 = 7'h46 == out_payload_rob_idx[6:0] ? rob_n_flits_70 : _GEN_4934; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4936 = 7'h47 == out_payload_rob_idx[6:0] ? rob_n_flits_71 : _GEN_4935; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4937 = 7'h48 == out_payload_rob_idx[6:0] ? rob_n_flits_72 : _GEN_4936; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4938 = 7'h49 == out_payload_rob_idx[6:0] ? rob_n_flits_73 : _GEN_4937; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4939 = 7'h4a == out_payload_rob_idx[6:0] ? rob_n_flits_74 : _GEN_4938; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4940 = 7'h4b == out_payload_rob_idx[6:0] ? rob_n_flits_75 : _GEN_4939; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4941 = 7'h4c == out_payload_rob_idx[6:0] ? rob_n_flits_76 : _GEN_4940; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4942 = 7'h4d == out_payload_rob_idx[6:0] ? rob_n_flits_77 : _GEN_4941; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4943 = 7'h4e == out_payload_rob_idx[6:0] ? rob_n_flits_78 : _GEN_4942; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4944 = 7'h4f == out_payload_rob_idx[6:0] ? rob_n_flits_79 : _GEN_4943; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4945 = 7'h50 == out_payload_rob_idx[6:0] ? rob_n_flits_80 : _GEN_4944; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4946 = 7'h51 == out_payload_rob_idx[6:0] ? rob_n_flits_81 : _GEN_4945; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4947 = 7'h52 == out_payload_rob_idx[6:0] ? rob_n_flits_82 : _GEN_4946; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4948 = 7'h53 == out_payload_rob_idx[6:0] ? rob_n_flits_83 : _GEN_4947; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4949 = 7'h54 == out_payload_rob_idx[6:0] ? rob_n_flits_84 : _GEN_4948; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4950 = 7'h55 == out_payload_rob_idx[6:0] ? rob_n_flits_85 : _GEN_4949; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4951 = 7'h56 == out_payload_rob_idx[6:0] ? rob_n_flits_86 : _GEN_4950; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4952 = 7'h57 == out_payload_rob_idx[6:0] ? rob_n_flits_87 : _GEN_4951; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4953 = 7'h58 == out_payload_rob_idx[6:0] ? rob_n_flits_88 : _GEN_4952; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4954 = 7'h59 == out_payload_rob_idx[6:0] ? rob_n_flits_89 : _GEN_4953; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4955 = 7'h5a == out_payload_rob_idx[6:0] ? rob_n_flits_90 : _GEN_4954; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4956 = 7'h5b == out_payload_rob_idx[6:0] ? rob_n_flits_91 : _GEN_4955; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4957 = 7'h5c == out_payload_rob_idx[6:0] ? rob_n_flits_92 : _GEN_4956; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4958 = 7'h5d == out_payload_rob_idx[6:0] ? rob_n_flits_93 : _GEN_4957; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4959 = 7'h5e == out_payload_rob_idx[6:0] ? rob_n_flits_94 : _GEN_4958; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4960 = 7'h5f == out_payload_rob_idx[6:0] ? rob_n_flits_95 : _GEN_4959; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4961 = 7'h60 == out_payload_rob_idx[6:0] ? rob_n_flits_96 : _GEN_4960; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4962 = 7'h61 == out_payload_rob_idx[6:0] ? rob_n_flits_97 : _GEN_4961; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4963 = 7'h62 == out_payload_rob_idx[6:0] ? rob_n_flits_98 : _GEN_4962; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4964 = 7'h63 == out_payload_rob_idx[6:0] ? rob_n_flits_99 : _GEN_4963; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4965 = 7'h64 == out_payload_rob_idx[6:0] ? rob_n_flits_100 : _GEN_4964; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4966 = 7'h65 == out_payload_rob_idx[6:0] ? rob_n_flits_101 : _GEN_4965; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4967 = 7'h66 == out_payload_rob_idx[6:0] ? rob_n_flits_102 : _GEN_4966; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4968 = 7'h67 == out_payload_rob_idx[6:0] ? rob_n_flits_103 : _GEN_4967; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4969 = 7'h68 == out_payload_rob_idx[6:0] ? rob_n_flits_104 : _GEN_4968; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4970 = 7'h69 == out_payload_rob_idx[6:0] ? rob_n_flits_105 : _GEN_4969; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4971 = 7'h6a == out_payload_rob_idx[6:0] ? rob_n_flits_106 : _GEN_4970; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4972 = 7'h6b == out_payload_rob_idx[6:0] ? rob_n_flits_107 : _GEN_4971; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4973 = 7'h6c == out_payload_rob_idx[6:0] ? rob_n_flits_108 : _GEN_4972; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4974 = 7'h6d == out_payload_rob_idx[6:0] ? rob_n_flits_109 : _GEN_4973; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4975 = 7'h6e == out_payload_rob_idx[6:0] ? rob_n_flits_110 : _GEN_4974; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4976 = 7'h6f == out_payload_rob_idx[6:0] ? rob_n_flits_111 : _GEN_4975; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4977 = 7'h70 == out_payload_rob_idx[6:0] ? rob_n_flits_112 : _GEN_4976; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4978 = 7'h71 == out_payload_rob_idx[6:0] ? rob_n_flits_113 : _GEN_4977; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4979 = 7'h72 == out_payload_rob_idx[6:0] ? rob_n_flits_114 : _GEN_4978; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4980 = 7'h73 == out_payload_rob_idx[6:0] ? rob_n_flits_115 : _GEN_4979; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4981 = 7'h74 == out_payload_rob_idx[6:0] ? rob_n_flits_116 : _GEN_4980; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4982 = 7'h75 == out_payload_rob_idx[6:0] ? rob_n_flits_117 : _GEN_4981; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4983 = 7'h76 == out_payload_rob_idx[6:0] ? rob_n_flits_118 : _GEN_4982; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4984 = 7'h77 == out_payload_rob_idx[6:0] ? rob_n_flits_119 : _GEN_4983; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4985 = 7'h78 == out_payload_rob_idx[6:0] ? rob_n_flits_120 : _GEN_4984; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4986 = 7'h79 == out_payload_rob_idx[6:0] ? rob_n_flits_121 : _GEN_4985; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4987 = 7'h7a == out_payload_rob_idx[6:0] ? rob_n_flits_122 : _GEN_4986; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4988 = 7'h7b == out_payload_rob_idx[6:0] ? rob_n_flits_123 : _GEN_4987; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4989 = 7'h7c == out_payload_rob_idx[6:0] ? rob_n_flits_124 : _GEN_4988; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4990 = 7'h7d == out_payload_rob_idx[6:0] ? rob_n_flits_125 : _GEN_4989; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4991 = 7'h7e == out_payload_rob_idx[6:0] ? rob_n_flits_126 : _GEN_4990; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_4992 = 7'h7f == out_payload_rob_idx[6:0] ? rob_n_flits_127 : _GEN_4991; // @[TestHarness.scala 205:{42,42}]
  wire [15:0] _GEN_7819 = {{9'd0}, packet_rob_idx}; // @[TestHarness.scala 206:61]
  wire  _T_76 = io_from_noc_0_flit_bits_head & enable_print_latency; // @[TestHarness.scala 208:30]
  wire [3:0] _rob_flits_returned_T_2 = _GEN_4864 + 4'h1; // @[TestHarness.scala 213:66]
  wire [3:0] _GEN_5249 = 7'h0 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3841; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5250 = 7'h1 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3842; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5251 = 7'h2 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3843; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5252 = 7'h3 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3844; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5253 = 7'h4 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3845; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5254 = 7'h5 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3846; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5255 = 7'h6 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3847; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5256 = 7'h7 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3848; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5257 = 7'h8 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3849; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5258 = 7'h9 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3850; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5259 = 7'ha == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3851; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5260 = 7'hb == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3852; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5261 = 7'hc == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3853; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5262 = 7'hd == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3854; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5263 = 7'he == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3855; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5264 = 7'hf == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3856; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5265 = 7'h10 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3857; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5266 = 7'h11 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3858; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5267 = 7'h12 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3859; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5268 = 7'h13 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3860; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5269 = 7'h14 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3861; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5270 = 7'h15 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3862; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5271 = 7'h16 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3863; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5272 = 7'h17 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3864; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5273 = 7'h18 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3865; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5274 = 7'h19 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3866; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5275 = 7'h1a == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3867; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5276 = 7'h1b == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3868; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5277 = 7'h1c == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3869; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5278 = 7'h1d == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3870; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5279 = 7'h1e == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3871; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5280 = 7'h1f == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3872; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5281 = 7'h20 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3873; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5282 = 7'h21 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3874; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5283 = 7'h22 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3875; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5284 = 7'h23 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3876; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5285 = 7'h24 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3877; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5286 = 7'h25 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3878; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5287 = 7'h26 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3879; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5288 = 7'h27 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3880; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5289 = 7'h28 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3881; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5290 = 7'h29 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3882; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5291 = 7'h2a == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3883; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5292 = 7'h2b == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3884; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5293 = 7'h2c == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3885; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5294 = 7'h2d == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3886; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5295 = 7'h2e == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3887; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5296 = 7'h2f == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3888; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5297 = 7'h30 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3889; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5298 = 7'h31 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3890; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5299 = 7'h32 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3891; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5300 = 7'h33 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3892; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5301 = 7'h34 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3893; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5302 = 7'h35 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3894; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5303 = 7'h36 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3895; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5304 = 7'h37 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3896; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5305 = 7'h38 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3897; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5306 = 7'h39 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3898; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5307 = 7'h3a == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3899; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5308 = 7'h3b == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3900; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5309 = 7'h3c == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3901; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5310 = 7'h3d == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3902; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5311 = 7'h3e == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3903; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5312 = 7'h3f == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3904; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5313 = 7'h40 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3905; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5314 = 7'h41 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3906; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5315 = 7'h42 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3907; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5316 = 7'h43 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3908; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5317 = 7'h44 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3909; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5318 = 7'h45 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3910; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5319 = 7'h46 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3911; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5320 = 7'h47 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3912; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5321 = 7'h48 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3913; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5322 = 7'h49 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3914; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5323 = 7'h4a == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3915; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5324 = 7'h4b == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3916; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5325 = 7'h4c == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3917; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5326 = 7'h4d == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3918; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5327 = 7'h4e == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3919; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5328 = 7'h4f == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3920; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5329 = 7'h50 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3921; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5330 = 7'h51 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3922; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5331 = 7'h52 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3923; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5332 = 7'h53 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3924; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5333 = 7'h54 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3925; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5334 = 7'h55 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3926; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5335 = 7'h56 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3927; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5336 = 7'h57 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3928; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5337 = 7'h58 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3929; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5338 = 7'h59 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3930; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5339 = 7'h5a == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3931; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5340 = 7'h5b == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3932; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5341 = 7'h5c == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3933; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5342 = 7'h5d == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3934; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5343 = 7'h5e == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3935; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5344 = 7'h5f == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3936; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5345 = 7'h60 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3937; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5346 = 7'h61 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3938; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5347 = 7'h62 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3939; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5348 = 7'h63 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3940; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5349 = 7'h64 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3941; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5350 = 7'h65 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3942; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5351 = 7'h66 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3943; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5352 = 7'h67 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3944; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5353 = 7'h68 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3945; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5354 = 7'h69 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3946; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5355 = 7'h6a == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3947; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5356 = 7'h6b == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3948; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5357 = 7'h6c == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3949; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5358 = 7'h6d == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3950; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5359 = 7'h6e == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3951; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5360 = 7'h6f == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3952; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5361 = 7'h70 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3953; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5362 = 7'h71 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3954; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5363 = 7'h72 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3955; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5364 = 7'h73 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3956; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5365 = 7'h74 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3957; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5366 = 7'h75 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3958; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5367 = 7'h76 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3959; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5368 = 7'h77 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3960; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5369 = 7'h78 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3961; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5370 = 7'h79 == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3962; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5371 = 7'h7a == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3963; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5372 = 7'h7b == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3964; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5373 = 7'h7c == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3965; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5374 = 7'h7d == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3966; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5375 = 7'h7e == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3967; // @[TestHarness.scala 213:{35,35}]
  wire [3:0] _GEN_5376 = 7'h7f == out_payload_rob_idx[6:0] ? _rob_flits_returned_T_2 : _GEN_3968; // @[TestHarness.scala 213:{35,35}]
  wire [15:0] _rob_payload_flits_fired_T_2 = _GEN_4480 + 16'h1; // @[TestHarness.scala 214:76]
  wire [15:0] _GEN_5505 = 7'h0 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3329; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5506 = 7'h1 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3330; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5507 = 7'h2 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3331; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5508 = 7'h3 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3332; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5509 = 7'h4 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3333; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5510 = 7'h5 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3334; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5511 = 7'h6 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3335; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5512 = 7'h7 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3336; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5513 = 7'h8 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3337; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5514 = 7'h9 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3338; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5515 = 7'ha == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3339; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5516 = 7'hb == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3340; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5517 = 7'hc == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3341; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5518 = 7'hd == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3342; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5519 = 7'he == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3343; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5520 = 7'hf == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3344; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5521 = 7'h10 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3345; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5522 = 7'h11 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3346; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5523 = 7'h12 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3347; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5524 = 7'h13 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3348; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5525 = 7'h14 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3349; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5526 = 7'h15 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3350; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5527 = 7'h16 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3351; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5528 = 7'h17 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3352; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5529 = 7'h18 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3353; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5530 = 7'h19 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3354; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5531 = 7'h1a == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3355; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5532 = 7'h1b == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3356; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5533 = 7'h1c == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3357; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5534 = 7'h1d == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3358; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5535 = 7'h1e == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3359; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5536 = 7'h1f == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3360; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5537 = 7'h20 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3361; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5538 = 7'h21 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3362; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5539 = 7'h22 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3363; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5540 = 7'h23 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3364; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5541 = 7'h24 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3365; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5542 = 7'h25 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3366; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5543 = 7'h26 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3367; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5544 = 7'h27 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3368; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5545 = 7'h28 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3369; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5546 = 7'h29 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3370; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5547 = 7'h2a == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3371; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5548 = 7'h2b == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3372; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5549 = 7'h2c == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3373; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5550 = 7'h2d == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3374; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5551 = 7'h2e == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3375; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5552 = 7'h2f == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3376; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5553 = 7'h30 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3377; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5554 = 7'h31 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3378; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5555 = 7'h32 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3379; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5556 = 7'h33 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3380; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5557 = 7'h34 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3381; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5558 = 7'h35 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3382; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5559 = 7'h36 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3383; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5560 = 7'h37 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3384; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5561 = 7'h38 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3385; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5562 = 7'h39 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3386; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5563 = 7'h3a == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3387; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5564 = 7'h3b == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3388; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5565 = 7'h3c == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3389; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5566 = 7'h3d == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3390; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5567 = 7'h3e == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3391; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5568 = 7'h3f == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3392; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5569 = 7'h40 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3393; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5570 = 7'h41 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3394; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5571 = 7'h42 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3395; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5572 = 7'h43 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3396; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5573 = 7'h44 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3397; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5574 = 7'h45 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3398; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5575 = 7'h46 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3399; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5576 = 7'h47 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3400; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5577 = 7'h48 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3401; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5578 = 7'h49 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3402; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5579 = 7'h4a == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3403; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5580 = 7'h4b == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3404; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5581 = 7'h4c == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3405; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5582 = 7'h4d == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3406; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5583 = 7'h4e == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3407; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5584 = 7'h4f == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3408; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5585 = 7'h50 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3409; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5586 = 7'h51 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3410; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5587 = 7'h52 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3411; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5588 = 7'h53 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3412; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5589 = 7'h54 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3413; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5590 = 7'h55 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3414; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5591 = 7'h56 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3415; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5592 = 7'h57 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3416; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5593 = 7'h58 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3417; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5594 = 7'h59 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3418; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5595 = 7'h5a == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3419; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5596 = 7'h5b == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3420; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5597 = 7'h5c == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3421; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5598 = 7'h5d == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3422; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5599 = 7'h5e == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3423; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5600 = 7'h5f == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3424; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5601 = 7'h60 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3425; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5602 = 7'h61 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3426; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5603 = 7'h62 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3427; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5604 = 7'h63 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3428; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5605 = 7'h64 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3429; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5606 = 7'h65 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3430; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5607 = 7'h66 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3431; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5608 = 7'h67 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3432; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5609 = 7'h68 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3433; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5610 = 7'h69 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3434; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5611 = 7'h6a == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3435; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5612 = 7'h6b == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3436; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5613 = 7'h6c == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3437; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5614 = 7'h6d == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3438; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5615 = 7'h6e == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3439; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5616 = 7'h6f == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3440; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5617 = 7'h70 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3441; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5618 = 7'h71 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3442; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5619 = 7'h72 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3443; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5620 = 7'h73 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3444; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5621 = 7'h74 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3445; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5622 = 7'h75 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3446; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5623 = 7'h76 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3447; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5624 = 7'h77 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3448; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5625 = 7'h78 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3449; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5626 = 7'h79 == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3450; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5627 = 7'h7a == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3451; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5628 = 7'h7b == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3452; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5629 = 7'h7c == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3453; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5630 = 7'h7d == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3454; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5631 = 7'h7e == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3455; // @[TestHarness.scala 214:{40,40}]
  wire [15:0] _GEN_5632 = 7'h7f == out_payload_rob_idx[6:0] ? _rob_payload_flits_fired_T_2 : _GEN_3456; // @[TestHarness.scala 214:{40,40}]
  wire  _GEN_5633 = io_from_noc_0_flit_bits_head | packet_valid; // @[TestHarness.scala 196:31 215:{31,46}]
  wire [15:0] _GEN_5634 = io_from_noc_0_flit_bits_head ? out_payload_rob_idx : {{9'd0}, packet_rob_idx}; // @[TestHarness.scala 197:29 215:{31,72}]
  wire [3:0] _GEN_5636 = _T_84 ? _GEN_5249 : _GEN_3841; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5637 = _T_84 ? _GEN_5250 : _GEN_3842; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5638 = _T_84 ? _GEN_5251 : _GEN_3843; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5639 = _T_84 ? _GEN_5252 : _GEN_3844; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5640 = _T_84 ? _GEN_5253 : _GEN_3845; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5641 = _T_84 ? _GEN_5254 : _GEN_3846; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5642 = _T_84 ? _GEN_5255 : _GEN_3847; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5643 = _T_84 ? _GEN_5256 : _GEN_3848; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5644 = _T_84 ? _GEN_5257 : _GEN_3849; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5645 = _T_84 ? _GEN_5258 : _GEN_3850; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5646 = _T_84 ? _GEN_5259 : _GEN_3851; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5647 = _T_84 ? _GEN_5260 : _GEN_3852; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5648 = _T_84 ? _GEN_5261 : _GEN_3853; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5649 = _T_84 ? _GEN_5262 : _GEN_3854; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5650 = _T_84 ? _GEN_5263 : _GEN_3855; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5651 = _T_84 ? _GEN_5264 : _GEN_3856; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5652 = _T_84 ? _GEN_5265 : _GEN_3857; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5653 = _T_84 ? _GEN_5266 : _GEN_3858; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5654 = _T_84 ? _GEN_5267 : _GEN_3859; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5655 = _T_84 ? _GEN_5268 : _GEN_3860; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5656 = _T_84 ? _GEN_5269 : _GEN_3861; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5657 = _T_84 ? _GEN_5270 : _GEN_3862; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5658 = _T_84 ? _GEN_5271 : _GEN_3863; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5659 = _T_84 ? _GEN_5272 : _GEN_3864; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5660 = _T_84 ? _GEN_5273 : _GEN_3865; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5661 = _T_84 ? _GEN_5274 : _GEN_3866; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5662 = _T_84 ? _GEN_5275 : _GEN_3867; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5663 = _T_84 ? _GEN_5276 : _GEN_3868; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5664 = _T_84 ? _GEN_5277 : _GEN_3869; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5665 = _T_84 ? _GEN_5278 : _GEN_3870; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5666 = _T_84 ? _GEN_5279 : _GEN_3871; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5667 = _T_84 ? _GEN_5280 : _GEN_3872; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5668 = _T_84 ? _GEN_5281 : _GEN_3873; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5669 = _T_84 ? _GEN_5282 : _GEN_3874; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5670 = _T_84 ? _GEN_5283 : _GEN_3875; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5671 = _T_84 ? _GEN_5284 : _GEN_3876; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5672 = _T_84 ? _GEN_5285 : _GEN_3877; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5673 = _T_84 ? _GEN_5286 : _GEN_3878; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5674 = _T_84 ? _GEN_5287 : _GEN_3879; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5675 = _T_84 ? _GEN_5288 : _GEN_3880; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5676 = _T_84 ? _GEN_5289 : _GEN_3881; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5677 = _T_84 ? _GEN_5290 : _GEN_3882; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5678 = _T_84 ? _GEN_5291 : _GEN_3883; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5679 = _T_84 ? _GEN_5292 : _GEN_3884; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5680 = _T_84 ? _GEN_5293 : _GEN_3885; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5681 = _T_84 ? _GEN_5294 : _GEN_3886; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5682 = _T_84 ? _GEN_5295 : _GEN_3887; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5683 = _T_84 ? _GEN_5296 : _GEN_3888; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5684 = _T_84 ? _GEN_5297 : _GEN_3889; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5685 = _T_84 ? _GEN_5298 : _GEN_3890; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5686 = _T_84 ? _GEN_5299 : _GEN_3891; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5687 = _T_84 ? _GEN_5300 : _GEN_3892; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5688 = _T_84 ? _GEN_5301 : _GEN_3893; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5689 = _T_84 ? _GEN_5302 : _GEN_3894; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5690 = _T_84 ? _GEN_5303 : _GEN_3895; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5691 = _T_84 ? _GEN_5304 : _GEN_3896; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5692 = _T_84 ? _GEN_5305 : _GEN_3897; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5693 = _T_84 ? _GEN_5306 : _GEN_3898; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5694 = _T_84 ? _GEN_5307 : _GEN_3899; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5695 = _T_84 ? _GEN_5308 : _GEN_3900; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5696 = _T_84 ? _GEN_5309 : _GEN_3901; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5697 = _T_84 ? _GEN_5310 : _GEN_3902; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5698 = _T_84 ? _GEN_5311 : _GEN_3903; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5699 = _T_84 ? _GEN_5312 : _GEN_3904; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5700 = _T_84 ? _GEN_5313 : _GEN_3905; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5701 = _T_84 ? _GEN_5314 : _GEN_3906; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5702 = _T_84 ? _GEN_5315 : _GEN_3907; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5703 = _T_84 ? _GEN_5316 : _GEN_3908; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5704 = _T_84 ? _GEN_5317 : _GEN_3909; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5705 = _T_84 ? _GEN_5318 : _GEN_3910; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5706 = _T_84 ? _GEN_5319 : _GEN_3911; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5707 = _T_84 ? _GEN_5320 : _GEN_3912; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5708 = _T_84 ? _GEN_5321 : _GEN_3913; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5709 = _T_84 ? _GEN_5322 : _GEN_3914; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5710 = _T_84 ? _GEN_5323 : _GEN_3915; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5711 = _T_84 ? _GEN_5324 : _GEN_3916; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5712 = _T_84 ? _GEN_5325 : _GEN_3917; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5713 = _T_84 ? _GEN_5326 : _GEN_3918; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5714 = _T_84 ? _GEN_5327 : _GEN_3919; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5715 = _T_84 ? _GEN_5328 : _GEN_3920; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5716 = _T_84 ? _GEN_5329 : _GEN_3921; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5717 = _T_84 ? _GEN_5330 : _GEN_3922; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5718 = _T_84 ? _GEN_5331 : _GEN_3923; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5719 = _T_84 ? _GEN_5332 : _GEN_3924; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5720 = _T_84 ? _GEN_5333 : _GEN_3925; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5721 = _T_84 ? _GEN_5334 : _GEN_3926; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5722 = _T_84 ? _GEN_5335 : _GEN_3927; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5723 = _T_84 ? _GEN_5336 : _GEN_3928; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5724 = _T_84 ? _GEN_5337 : _GEN_3929; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5725 = _T_84 ? _GEN_5338 : _GEN_3930; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5726 = _T_84 ? _GEN_5339 : _GEN_3931; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5727 = _T_84 ? _GEN_5340 : _GEN_3932; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5728 = _T_84 ? _GEN_5341 : _GEN_3933; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5729 = _T_84 ? _GEN_5342 : _GEN_3934; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5730 = _T_84 ? _GEN_5343 : _GEN_3935; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5731 = _T_84 ? _GEN_5344 : _GEN_3936; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5732 = _T_84 ? _GEN_5345 : _GEN_3937; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5733 = _T_84 ? _GEN_5346 : _GEN_3938; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5734 = _T_84 ? _GEN_5347 : _GEN_3939; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5735 = _T_84 ? _GEN_5348 : _GEN_3940; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5736 = _T_84 ? _GEN_5349 : _GEN_3941; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5737 = _T_84 ? _GEN_5350 : _GEN_3942; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5738 = _T_84 ? _GEN_5351 : _GEN_3943; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5739 = _T_84 ? _GEN_5352 : _GEN_3944; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5740 = _T_84 ? _GEN_5353 : _GEN_3945; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5741 = _T_84 ? _GEN_5354 : _GEN_3946; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5742 = _T_84 ? _GEN_5355 : _GEN_3947; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5743 = _T_84 ? _GEN_5356 : _GEN_3948; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5744 = _T_84 ? _GEN_5357 : _GEN_3949; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5745 = _T_84 ? _GEN_5358 : _GEN_3950; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5746 = _T_84 ? _GEN_5359 : _GEN_3951; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5747 = _T_84 ? _GEN_5360 : _GEN_3952; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5748 = _T_84 ? _GEN_5361 : _GEN_3953; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5749 = _T_84 ? _GEN_5362 : _GEN_3954; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5750 = _T_84 ? _GEN_5363 : _GEN_3955; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5751 = _T_84 ? _GEN_5364 : _GEN_3956; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5752 = _T_84 ? _GEN_5365 : _GEN_3957; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5753 = _T_84 ? _GEN_5366 : _GEN_3958; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5754 = _T_84 ? _GEN_5367 : _GEN_3959; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5755 = _T_84 ? _GEN_5368 : _GEN_3960; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5756 = _T_84 ? _GEN_5369 : _GEN_3961; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5757 = _T_84 ? _GEN_5370 : _GEN_3962; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5758 = _T_84 ? _GEN_5371 : _GEN_3963; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5759 = _T_84 ? _GEN_5372 : _GEN_3964; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5760 = _T_84 ? _GEN_5373 : _GEN_3965; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5761 = _T_84 ? _GEN_5374 : _GEN_3966; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5762 = _T_84 ? _GEN_5375 : _GEN_3967; // @[TestHarness.scala 199:26]
  wire [3:0] _GEN_5763 = _T_84 ? _GEN_5376 : _GEN_3968; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5764 = _T_84 ? _GEN_5505 : _GEN_3329; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5765 = _T_84 ? _GEN_5506 : _GEN_3330; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5766 = _T_84 ? _GEN_5507 : _GEN_3331; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5767 = _T_84 ? _GEN_5508 : _GEN_3332; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5768 = _T_84 ? _GEN_5509 : _GEN_3333; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5769 = _T_84 ? _GEN_5510 : _GEN_3334; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5770 = _T_84 ? _GEN_5511 : _GEN_3335; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5771 = _T_84 ? _GEN_5512 : _GEN_3336; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5772 = _T_84 ? _GEN_5513 : _GEN_3337; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5773 = _T_84 ? _GEN_5514 : _GEN_3338; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5774 = _T_84 ? _GEN_5515 : _GEN_3339; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5775 = _T_84 ? _GEN_5516 : _GEN_3340; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5776 = _T_84 ? _GEN_5517 : _GEN_3341; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5777 = _T_84 ? _GEN_5518 : _GEN_3342; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5778 = _T_84 ? _GEN_5519 : _GEN_3343; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5779 = _T_84 ? _GEN_5520 : _GEN_3344; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5780 = _T_84 ? _GEN_5521 : _GEN_3345; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5781 = _T_84 ? _GEN_5522 : _GEN_3346; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5782 = _T_84 ? _GEN_5523 : _GEN_3347; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5783 = _T_84 ? _GEN_5524 : _GEN_3348; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5784 = _T_84 ? _GEN_5525 : _GEN_3349; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5785 = _T_84 ? _GEN_5526 : _GEN_3350; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5786 = _T_84 ? _GEN_5527 : _GEN_3351; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5787 = _T_84 ? _GEN_5528 : _GEN_3352; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5788 = _T_84 ? _GEN_5529 : _GEN_3353; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5789 = _T_84 ? _GEN_5530 : _GEN_3354; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5790 = _T_84 ? _GEN_5531 : _GEN_3355; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5791 = _T_84 ? _GEN_5532 : _GEN_3356; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5792 = _T_84 ? _GEN_5533 : _GEN_3357; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5793 = _T_84 ? _GEN_5534 : _GEN_3358; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5794 = _T_84 ? _GEN_5535 : _GEN_3359; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5795 = _T_84 ? _GEN_5536 : _GEN_3360; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5796 = _T_84 ? _GEN_5537 : _GEN_3361; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5797 = _T_84 ? _GEN_5538 : _GEN_3362; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5798 = _T_84 ? _GEN_5539 : _GEN_3363; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5799 = _T_84 ? _GEN_5540 : _GEN_3364; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5800 = _T_84 ? _GEN_5541 : _GEN_3365; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5801 = _T_84 ? _GEN_5542 : _GEN_3366; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5802 = _T_84 ? _GEN_5543 : _GEN_3367; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5803 = _T_84 ? _GEN_5544 : _GEN_3368; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5804 = _T_84 ? _GEN_5545 : _GEN_3369; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5805 = _T_84 ? _GEN_5546 : _GEN_3370; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5806 = _T_84 ? _GEN_5547 : _GEN_3371; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5807 = _T_84 ? _GEN_5548 : _GEN_3372; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5808 = _T_84 ? _GEN_5549 : _GEN_3373; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5809 = _T_84 ? _GEN_5550 : _GEN_3374; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5810 = _T_84 ? _GEN_5551 : _GEN_3375; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5811 = _T_84 ? _GEN_5552 : _GEN_3376; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5812 = _T_84 ? _GEN_5553 : _GEN_3377; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5813 = _T_84 ? _GEN_5554 : _GEN_3378; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5814 = _T_84 ? _GEN_5555 : _GEN_3379; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5815 = _T_84 ? _GEN_5556 : _GEN_3380; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5816 = _T_84 ? _GEN_5557 : _GEN_3381; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5817 = _T_84 ? _GEN_5558 : _GEN_3382; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5818 = _T_84 ? _GEN_5559 : _GEN_3383; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5819 = _T_84 ? _GEN_5560 : _GEN_3384; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5820 = _T_84 ? _GEN_5561 : _GEN_3385; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5821 = _T_84 ? _GEN_5562 : _GEN_3386; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5822 = _T_84 ? _GEN_5563 : _GEN_3387; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5823 = _T_84 ? _GEN_5564 : _GEN_3388; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5824 = _T_84 ? _GEN_5565 : _GEN_3389; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5825 = _T_84 ? _GEN_5566 : _GEN_3390; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5826 = _T_84 ? _GEN_5567 : _GEN_3391; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5827 = _T_84 ? _GEN_5568 : _GEN_3392; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5828 = _T_84 ? _GEN_5569 : _GEN_3393; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5829 = _T_84 ? _GEN_5570 : _GEN_3394; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5830 = _T_84 ? _GEN_5571 : _GEN_3395; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5831 = _T_84 ? _GEN_5572 : _GEN_3396; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5832 = _T_84 ? _GEN_5573 : _GEN_3397; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5833 = _T_84 ? _GEN_5574 : _GEN_3398; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5834 = _T_84 ? _GEN_5575 : _GEN_3399; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5835 = _T_84 ? _GEN_5576 : _GEN_3400; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5836 = _T_84 ? _GEN_5577 : _GEN_3401; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5837 = _T_84 ? _GEN_5578 : _GEN_3402; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5838 = _T_84 ? _GEN_5579 : _GEN_3403; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5839 = _T_84 ? _GEN_5580 : _GEN_3404; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5840 = _T_84 ? _GEN_5581 : _GEN_3405; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5841 = _T_84 ? _GEN_5582 : _GEN_3406; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5842 = _T_84 ? _GEN_5583 : _GEN_3407; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5843 = _T_84 ? _GEN_5584 : _GEN_3408; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5844 = _T_84 ? _GEN_5585 : _GEN_3409; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5845 = _T_84 ? _GEN_5586 : _GEN_3410; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5846 = _T_84 ? _GEN_5587 : _GEN_3411; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5847 = _T_84 ? _GEN_5588 : _GEN_3412; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5848 = _T_84 ? _GEN_5589 : _GEN_3413; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5849 = _T_84 ? _GEN_5590 : _GEN_3414; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5850 = _T_84 ? _GEN_5591 : _GEN_3415; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5851 = _T_84 ? _GEN_5592 : _GEN_3416; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5852 = _T_84 ? _GEN_5593 : _GEN_3417; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5853 = _T_84 ? _GEN_5594 : _GEN_3418; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5854 = _T_84 ? _GEN_5595 : _GEN_3419; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5855 = _T_84 ? _GEN_5596 : _GEN_3420; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5856 = _T_84 ? _GEN_5597 : _GEN_3421; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5857 = _T_84 ? _GEN_5598 : _GEN_3422; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5858 = _T_84 ? _GEN_5599 : _GEN_3423; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5859 = _T_84 ? _GEN_5600 : _GEN_3424; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5860 = _T_84 ? _GEN_5601 : _GEN_3425; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5861 = _T_84 ? _GEN_5602 : _GEN_3426; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5862 = _T_84 ? _GEN_5603 : _GEN_3427; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5863 = _T_84 ? _GEN_5604 : _GEN_3428; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5864 = _T_84 ? _GEN_5605 : _GEN_3429; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5865 = _T_84 ? _GEN_5606 : _GEN_3430; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5866 = _T_84 ? _GEN_5607 : _GEN_3431; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5867 = _T_84 ? _GEN_5608 : _GEN_3432; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5868 = _T_84 ? _GEN_5609 : _GEN_3433; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5869 = _T_84 ? _GEN_5610 : _GEN_3434; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5870 = _T_84 ? _GEN_5611 : _GEN_3435; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5871 = _T_84 ? _GEN_5612 : _GEN_3436; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5872 = _T_84 ? _GEN_5613 : _GEN_3437; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5873 = _T_84 ? _GEN_5614 : _GEN_3438; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5874 = _T_84 ? _GEN_5615 : _GEN_3439; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5875 = _T_84 ? _GEN_5616 : _GEN_3440; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5876 = _T_84 ? _GEN_5617 : _GEN_3441; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5877 = _T_84 ? _GEN_5618 : _GEN_3442; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5878 = _T_84 ? _GEN_5619 : _GEN_3443; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5879 = _T_84 ? _GEN_5620 : _GEN_3444; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5880 = _T_84 ? _GEN_5621 : _GEN_3445; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5881 = _T_84 ? _GEN_5622 : _GEN_3446; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5882 = _T_84 ? _GEN_5623 : _GEN_3447; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5883 = _T_84 ? _GEN_5624 : _GEN_3448; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5884 = _T_84 ? _GEN_5625 : _GEN_3449; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5885 = _T_84 ? _GEN_5626 : _GEN_3450; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5886 = _T_84 ? _GEN_5627 : _GEN_3451; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5887 = _T_84 ? _GEN_5628 : _GEN_3452; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5888 = _T_84 ? _GEN_5629 : _GEN_3453; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5889 = _T_84 ? _GEN_5630 : _GEN_3454; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5890 = _T_84 ? _GEN_5631 : _GEN_3455; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5891 = _T_84 ? _GEN_5632 : _GEN_3456; // @[TestHarness.scala 199:26]
  wire [15:0] _GEN_5893 = _T_84 ? _GEN_5634 : {{9'd0}, packet_rob_idx}; // @[TestHarness.scala 199:26 197:29]
  wire [31:0] out_payload_1_tsc = io_from_noc_1_flit_bits_payload[63:32]; // @[TestHarness.scala 194:51]
  reg  packet_valid_1; // @[TestHarness.scala 196:31]
  reg [6:0] packet_rob_idx_1; // @[TestHarness.scala 197:29]
  wire [127:0] _T_89 = rob_valids >> out_payload_1_rob_idx; // @[TestHarness.scala 201:24]
  wire [31:0] _GEN_5895 = 7'h1 == out_payload_1_rob_idx[6:0] ? rob_payload_1_tsc : rob_payload_0_tsc; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5896 = 7'h2 == out_payload_1_rob_idx[6:0] ? rob_payload_2_tsc : _GEN_5895; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5897 = 7'h3 == out_payload_1_rob_idx[6:0] ? rob_payload_3_tsc : _GEN_5896; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5898 = 7'h4 == out_payload_1_rob_idx[6:0] ? rob_payload_4_tsc : _GEN_5897; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5899 = 7'h5 == out_payload_1_rob_idx[6:0] ? rob_payload_5_tsc : _GEN_5898; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5900 = 7'h6 == out_payload_1_rob_idx[6:0] ? rob_payload_6_tsc : _GEN_5899; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5901 = 7'h7 == out_payload_1_rob_idx[6:0] ? rob_payload_7_tsc : _GEN_5900; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5902 = 7'h8 == out_payload_1_rob_idx[6:0] ? rob_payload_8_tsc : _GEN_5901; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5903 = 7'h9 == out_payload_1_rob_idx[6:0] ? rob_payload_9_tsc : _GEN_5902; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5904 = 7'ha == out_payload_1_rob_idx[6:0] ? rob_payload_10_tsc : _GEN_5903; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5905 = 7'hb == out_payload_1_rob_idx[6:0] ? rob_payload_11_tsc : _GEN_5904; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5906 = 7'hc == out_payload_1_rob_idx[6:0] ? rob_payload_12_tsc : _GEN_5905; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5907 = 7'hd == out_payload_1_rob_idx[6:0] ? rob_payload_13_tsc : _GEN_5906; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5908 = 7'he == out_payload_1_rob_idx[6:0] ? rob_payload_14_tsc : _GEN_5907; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5909 = 7'hf == out_payload_1_rob_idx[6:0] ? rob_payload_15_tsc : _GEN_5908; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5910 = 7'h10 == out_payload_1_rob_idx[6:0] ? rob_payload_16_tsc : _GEN_5909; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5911 = 7'h11 == out_payload_1_rob_idx[6:0] ? rob_payload_17_tsc : _GEN_5910; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5912 = 7'h12 == out_payload_1_rob_idx[6:0] ? rob_payload_18_tsc : _GEN_5911; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5913 = 7'h13 == out_payload_1_rob_idx[6:0] ? rob_payload_19_tsc : _GEN_5912; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5914 = 7'h14 == out_payload_1_rob_idx[6:0] ? rob_payload_20_tsc : _GEN_5913; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5915 = 7'h15 == out_payload_1_rob_idx[6:0] ? rob_payload_21_tsc : _GEN_5914; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5916 = 7'h16 == out_payload_1_rob_idx[6:0] ? rob_payload_22_tsc : _GEN_5915; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5917 = 7'h17 == out_payload_1_rob_idx[6:0] ? rob_payload_23_tsc : _GEN_5916; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5918 = 7'h18 == out_payload_1_rob_idx[6:0] ? rob_payload_24_tsc : _GEN_5917; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5919 = 7'h19 == out_payload_1_rob_idx[6:0] ? rob_payload_25_tsc : _GEN_5918; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5920 = 7'h1a == out_payload_1_rob_idx[6:0] ? rob_payload_26_tsc : _GEN_5919; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5921 = 7'h1b == out_payload_1_rob_idx[6:0] ? rob_payload_27_tsc : _GEN_5920; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5922 = 7'h1c == out_payload_1_rob_idx[6:0] ? rob_payload_28_tsc : _GEN_5921; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5923 = 7'h1d == out_payload_1_rob_idx[6:0] ? rob_payload_29_tsc : _GEN_5922; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5924 = 7'h1e == out_payload_1_rob_idx[6:0] ? rob_payload_30_tsc : _GEN_5923; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5925 = 7'h1f == out_payload_1_rob_idx[6:0] ? rob_payload_31_tsc : _GEN_5924; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5926 = 7'h20 == out_payload_1_rob_idx[6:0] ? rob_payload_32_tsc : _GEN_5925; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5927 = 7'h21 == out_payload_1_rob_idx[6:0] ? rob_payload_33_tsc : _GEN_5926; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5928 = 7'h22 == out_payload_1_rob_idx[6:0] ? rob_payload_34_tsc : _GEN_5927; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5929 = 7'h23 == out_payload_1_rob_idx[6:0] ? rob_payload_35_tsc : _GEN_5928; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5930 = 7'h24 == out_payload_1_rob_idx[6:0] ? rob_payload_36_tsc : _GEN_5929; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5931 = 7'h25 == out_payload_1_rob_idx[6:0] ? rob_payload_37_tsc : _GEN_5930; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5932 = 7'h26 == out_payload_1_rob_idx[6:0] ? rob_payload_38_tsc : _GEN_5931; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5933 = 7'h27 == out_payload_1_rob_idx[6:0] ? rob_payload_39_tsc : _GEN_5932; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5934 = 7'h28 == out_payload_1_rob_idx[6:0] ? rob_payload_40_tsc : _GEN_5933; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5935 = 7'h29 == out_payload_1_rob_idx[6:0] ? rob_payload_41_tsc : _GEN_5934; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5936 = 7'h2a == out_payload_1_rob_idx[6:0] ? rob_payload_42_tsc : _GEN_5935; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5937 = 7'h2b == out_payload_1_rob_idx[6:0] ? rob_payload_43_tsc : _GEN_5936; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5938 = 7'h2c == out_payload_1_rob_idx[6:0] ? rob_payload_44_tsc : _GEN_5937; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5939 = 7'h2d == out_payload_1_rob_idx[6:0] ? rob_payload_45_tsc : _GEN_5938; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5940 = 7'h2e == out_payload_1_rob_idx[6:0] ? rob_payload_46_tsc : _GEN_5939; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5941 = 7'h2f == out_payload_1_rob_idx[6:0] ? rob_payload_47_tsc : _GEN_5940; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5942 = 7'h30 == out_payload_1_rob_idx[6:0] ? rob_payload_48_tsc : _GEN_5941; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5943 = 7'h31 == out_payload_1_rob_idx[6:0] ? rob_payload_49_tsc : _GEN_5942; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5944 = 7'h32 == out_payload_1_rob_idx[6:0] ? rob_payload_50_tsc : _GEN_5943; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5945 = 7'h33 == out_payload_1_rob_idx[6:0] ? rob_payload_51_tsc : _GEN_5944; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5946 = 7'h34 == out_payload_1_rob_idx[6:0] ? rob_payload_52_tsc : _GEN_5945; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5947 = 7'h35 == out_payload_1_rob_idx[6:0] ? rob_payload_53_tsc : _GEN_5946; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5948 = 7'h36 == out_payload_1_rob_idx[6:0] ? rob_payload_54_tsc : _GEN_5947; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5949 = 7'h37 == out_payload_1_rob_idx[6:0] ? rob_payload_55_tsc : _GEN_5948; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5950 = 7'h38 == out_payload_1_rob_idx[6:0] ? rob_payload_56_tsc : _GEN_5949; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5951 = 7'h39 == out_payload_1_rob_idx[6:0] ? rob_payload_57_tsc : _GEN_5950; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5952 = 7'h3a == out_payload_1_rob_idx[6:0] ? rob_payload_58_tsc : _GEN_5951; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5953 = 7'h3b == out_payload_1_rob_idx[6:0] ? rob_payload_59_tsc : _GEN_5952; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5954 = 7'h3c == out_payload_1_rob_idx[6:0] ? rob_payload_60_tsc : _GEN_5953; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5955 = 7'h3d == out_payload_1_rob_idx[6:0] ? rob_payload_61_tsc : _GEN_5954; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5956 = 7'h3e == out_payload_1_rob_idx[6:0] ? rob_payload_62_tsc : _GEN_5955; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5957 = 7'h3f == out_payload_1_rob_idx[6:0] ? rob_payload_63_tsc : _GEN_5956; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5958 = 7'h40 == out_payload_1_rob_idx[6:0] ? rob_payload_64_tsc : _GEN_5957; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5959 = 7'h41 == out_payload_1_rob_idx[6:0] ? rob_payload_65_tsc : _GEN_5958; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5960 = 7'h42 == out_payload_1_rob_idx[6:0] ? rob_payload_66_tsc : _GEN_5959; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5961 = 7'h43 == out_payload_1_rob_idx[6:0] ? rob_payload_67_tsc : _GEN_5960; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5962 = 7'h44 == out_payload_1_rob_idx[6:0] ? rob_payload_68_tsc : _GEN_5961; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5963 = 7'h45 == out_payload_1_rob_idx[6:0] ? rob_payload_69_tsc : _GEN_5962; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5964 = 7'h46 == out_payload_1_rob_idx[6:0] ? rob_payload_70_tsc : _GEN_5963; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5965 = 7'h47 == out_payload_1_rob_idx[6:0] ? rob_payload_71_tsc : _GEN_5964; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5966 = 7'h48 == out_payload_1_rob_idx[6:0] ? rob_payload_72_tsc : _GEN_5965; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5967 = 7'h49 == out_payload_1_rob_idx[6:0] ? rob_payload_73_tsc : _GEN_5966; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5968 = 7'h4a == out_payload_1_rob_idx[6:0] ? rob_payload_74_tsc : _GEN_5967; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5969 = 7'h4b == out_payload_1_rob_idx[6:0] ? rob_payload_75_tsc : _GEN_5968; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5970 = 7'h4c == out_payload_1_rob_idx[6:0] ? rob_payload_76_tsc : _GEN_5969; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5971 = 7'h4d == out_payload_1_rob_idx[6:0] ? rob_payload_77_tsc : _GEN_5970; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5972 = 7'h4e == out_payload_1_rob_idx[6:0] ? rob_payload_78_tsc : _GEN_5971; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5973 = 7'h4f == out_payload_1_rob_idx[6:0] ? rob_payload_79_tsc : _GEN_5972; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5974 = 7'h50 == out_payload_1_rob_idx[6:0] ? rob_payload_80_tsc : _GEN_5973; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5975 = 7'h51 == out_payload_1_rob_idx[6:0] ? rob_payload_81_tsc : _GEN_5974; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5976 = 7'h52 == out_payload_1_rob_idx[6:0] ? rob_payload_82_tsc : _GEN_5975; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5977 = 7'h53 == out_payload_1_rob_idx[6:0] ? rob_payload_83_tsc : _GEN_5976; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5978 = 7'h54 == out_payload_1_rob_idx[6:0] ? rob_payload_84_tsc : _GEN_5977; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5979 = 7'h55 == out_payload_1_rob_idx[6:0] ? rob_payload_85_tsc : _GEN_5978; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5980 = 7'h56 == out_payload_1_rob_idx[6:0] ? rob_payload_86_tsc : _GEN_5979; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5981 = 7'h57 == out_payload_1_rob_idx[6:0] ? rob_payload_87_tsc : _GEN_5980; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5982 = 7'h58 == out_payload_1_rob_idx[6:0] ? rob_payload_88_tsc : _GEN_5981; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5983 = 7'h59 == out_payload_1_rob_idx[6:0] ? rob_payload_89_tsc : _GEN_5982; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5984 = 7'h5a == out_payload_1_rob_idx[6:0] ? rob_payload_90_tsc : _GEN_5983; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5985 = 7'h5b == out_payload_1_rob_idx[6:0] ? rob_payload_91_tsc : _GEN_5984; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5986 = 7'h5c == out_payload_1_rob_idx[6:0] ? rob_payload_92_tsc : _GEN_5985; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5987 = 7'h5d == out_payload_1_rob_idx[6:0] ? rob_payload_93_tsc : _GEN_5986; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5988 = 7'h5e == out_payload_1_rob_idx[6:0] ? rob_payload_94_tsc : _GEN_5987; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5989 = 7'h5f == out_payload_1_rob_idx[6:0] ? rob_payload_95_tsc : _GEN_5988; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5990 = 7'h60 == out_payload_1_rob_idx[6:0] ? rob_payload_96_tsc : _GEN_5989; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5991 = 7'h61 == out_payload_1_rob_idx[6:0] ? rob_payload_97_tsc : _GEN_5990; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5992 = 7'h62 == out_payload_1_rob_idx[6:0] ? rob_payload_98_tsc : _GEN_5991; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5993 = 7'h63 == out_payload_1_rob_idx[6:0] ? rob_payload_99_tsc : _GEN_5992; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5994 = 7'h64 == out_payload_1_rob_idx[6:0] ? rob_payload_100_tsc : _GEN_5993; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5995 = 7'h65 == out_payload_1_rob_idx[6:0] ? rob_payload_101_tsc : _GEN_5994; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5996 = 7'h66 == out_payload_1_rob_idx[6:0] ? rob_payload_102_tsc : _GEN_5995; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5997 = 7'h67 == out_payload_1_rob_idx[6:0] ? rob_payload_103_tsc : _GEN_5996; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5998 = 7'h68 == out_payload_1_rob_idx[6:0] ? rob_payload_104_tsc : _GEN_5997; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_5999 = 7'h69 == out_payload_1_rob_idx[6:0] ? rob_payload_105_tsc : _GEN_5998; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_6000 = 7'h6a == out_payload_1_rob_idx[6:0] ? rob_payload_106_tsc : _GEN_5999; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_6001 = 7'h6b == out_payload_1_rob_idx[6:0] ? rob_payload_107_tsc : _GEN_6000; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_6002 = 7'h6c == out_payload_1_rob_idx[6:0] ? rob_payload_108_tsc : _GEN_6001; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_6003 = 7'h6d == out_payload_1_rob_idx[6:0] ? rob_payload_109_tsc : _GEN_6002; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_6004 = 7'h6e == out_payload_1_rob_idx[6:0] ? rob_payload_110_tsc : _GEN_6003; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_6005 = 7'h6f == out_payload_1_rob_idx[6:0] ? rob_payload_111_tsc : _GEN_6004; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_6006 = 7'h70 == out_payload_1_rob_idx[6:0] ? rob_payload_112_tsc : _GEN_6005; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_6007 = 7'h71 == out_payload_1_rob_idx[6:0] ? rob_payload_113_tsc : _GEN_6006; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_6008 = 7'h72 == out_payload_1_rob_idx[6:0] ? rob_payload_114_tsc : _GEN_6007; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_6009 = 7'h73 == out_payload_1_rob_idx[6:0] ? rob_payload_115_tsc : _GEN_6008; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_6010 = 7'h74 == out_payload_1_rob_idx[6:0] ? rob_payload_116_tsc : _GEN_6009; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_6011 = 7'h75 == out_payload_1_rob_idx[6:0] ? rob_payload_117_tsc : _GEN_6010; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_6012 = 7'h76 == out_payload_1_rob_idx[6:0] ? rob_payload_118_tsc : _GEN_6011; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_6013 = 7'h77 == out_payload_1_rob_idx[6:0] ? rob_payload_119_tsc : _GEN_6012; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_6014 = 7'h78 == out_payload_1_rob_idx[6:0] ? rob_payload_120_tsc : _GEN_6013; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_6015 = 7'h79 == out_payload_1_rob_idx[6:0] ? rob_payload_121_tsc : _GEN_6014; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_6016 = 7'h7a == out_payload_1_rob_idx[6:0] ? rob_payload_122_tsc : _GEN_6015; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_6017 = 7'h7b == out_payload_1_rob_idx[6:0] ? rob_payload_123_tsc : _GEN_6016; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_6018 = 7'h7c == out_payload_1_rob_idx[6:0] ? rob_payload_124_tsc : _GEN_6017; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_6019 = 7'h7d == out_payload_1_rob_idx[6:0] ? rob_payload_125_tsc : _GEN_6018; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_6020 = 7'h7e == out_payload_1_rob_idx[6:0] ? rob_payload_126_tsc : _GEN_6019; // @[TestHarness.scala 202:{35,35}]
  wire [31:0] _GEN_6021 = 7'h7f == out_payload_1_rob_idx[6:0] ? rob_payload_127_tsc : _GEN_6020; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6023 = 7'h1 == out_payload_1_rob_idx[6:0] ? rob_payload_1_rob_idx : rob_payload_0_rob_idx; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6024 = 7'h2 == out_payload_1_rob_idx[6:0] ? rob_payload_2_rob_idx : _GEN_6023; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6025 = 7'h3 == out_payload_1_rob_idx[6:0] ? rob_payload_3_rob_idx : _GEN_6024; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6026 = 7'h4 == out_payload_1_rob_idx[6:0] ? rob_payload_4_rob_idx : _GEN_6025; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6027 = 7'h5 == out_payload_1_rob_idx[6:0] ? rob_payload_5_rob_idx : _GEN_6026; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6028 = 7'h6 == out_payload_1_rob_idx[6:0] ? rob_payload_6_rob_idx : _GEN_6027; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6029 = 7'h7 == out_payload_1_rob_idx[6:0] ? rob_payload_7_rob_idx : _GEN_6028; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6030 = 7'h8 == out_payload_1_rob_idx[6:0] ? rob_payload_8_rob_idx : _GEN_6029; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6031 = 7'h9 == out_payload_1_rob_idx[6:0] ? rob_payload_9_rob_idx : _GEN_6030; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6032 = 7'ha == out_payload_1_rob_idx[6:0] ? rob_payload_10_rob_idx : _GEN_6031; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6033 = 7'hb == out_payload_1_rob_idx[6:0] ? rob_payload_11_rob_idx : _GEN_6032; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6034 = 7'hc == out_payload_1_rob_idx[6:0] ? rob_payload_12_rob_idx : _GEN_6033; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6035 = 7'hd == out_payload_1_rob_idx[6:0] ? rob_payload_13_rob_idx : _GEN_6034; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6036 = 7'he == out_payload_1_rob_idx[6:0] ? rob_payload_14_rob_idx : _GEN_6035; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6037 = 7'hf == out_payload_1_rob_idx[6:0] ? rob_payload_15_rob_idx : _GEN_6036; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6038 = 7'h10 == out_payload_1_rob_idx[6:0] ? rob_payload_16_rob_idx : _GEN_6037; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6039 = 7'h11 == out_payload_1_rob_idx[6:0] ? rob_payload_17_rob_idx : _GEN_6038; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6040 = 7'h12 == out_payload_1_rob_idx[6:0] ? rob_payload_18_rob_idx : _GEN_6039; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6041 = 7'h13 == out_payload_1_rob_idx[6:0] ? rob_payload_19_rob_idx : _GEN_6040; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6042 = 7'h14 == out_payload_1_rob_idx[6:0] ? rob_payload_20_rob_idx : _GEN_6041; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6043 = 7'h15 == out_payload_1_rob_idx[6:0] ? rob_payload_21_rob_idx : _GEN_6042; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6044 = 7'h16 == out_payload_1_rob_idx[6:0] ? rob_payload_22_rob_idx : _GEN_6043; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6045 = 7'h17 == out_payload_1_rob_idx[6:0] ? rob_payload_23_rob_idx : _GEN_6044; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6046 = 7'h18 == out_payload_1_rob_idx[6:0] ? rob_payload_24_rob_idx : _GEN_6045; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6047 = 7'h19 == out_payload_1_rob_idx[6:0] ? rob_payload_25_rob_idx : _GEN_6046; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6048 = 7'h1a == out_payload_1_rob_idx[6:0] ? rob_payload_26_rob_idx : _GEN_6047; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6049 = 7'h1b == out_payload_1_rob_idx[6:0] ? rob_payload_27_rob_idx : _GEN_6048; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6050 = 7'h1c == out_payload_1_rob_idx[6:0] ? rob_payload_28_rob_idx : _GEN_6049; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6051 = 7'h1d == out_payload_1_rob_idx[6:0] ? rob_payload_29_rob_idx : _GEN_6050; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6052 = 7'h1e == out_payload_1_rob_idx[6:0] ? rob_payload_30_rob_idx : _GEN_6051; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6053 = 7'h1f == out_payload_1_rob_idx[6:0] ? rob_payload_31_rob_idx : _GEN_6052; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6054 = 7'h20 == out_payload_1_rob_idx[6:0] ? rob_payload_32_rob_idx : _GEN_6053; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6055 = 7'h21 == out_payload_1_rob_idx[6:0] ? rob_payload_33_rob_idx : _GEN_6054; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6056 = 7'h22 == out_payload_1_rob_idx[6:0] ? rob_payload_34_rob_idx : _GEN_6055; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6057 = 7'h23 == out_payload_1_rob_idx[6:0] ? rob_payload_35_rob_idx : _GEN_6056; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6058 = 7'h24 == out_payload_1_rob_idx[6:0] ? rob_payload_36_rob_idx : _GEN_6057; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6059 = 7'h25 == out_payload_1_rob_idx[6:0] ? rob_payload_37_rob_idx : _GEN_6058; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6060 = 7'h26 == out_payload_1_rob_idx[6:0] ? rob_payload_38_rob_idx : _GEN_6059; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6061 = 7'h27 == out_payload_1_rob_idx[6:0] ? rob_payload_39_rob_idx : _GEN_6060; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6062 = 7'h28 == out_payload_1_rob_idx[6:0] ? rob_payload_40_rob_idx : _GEN_6061; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6063 = 7'h29 == out_payload_1_rob_idx[6:0] ? rob_payload_41_rob_idx : _GEN_6062; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6064 = 7'h2a == out_payload_1_rob_idx[6:0] ? rob_payload_42_rob_idx : _GEN_6063; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6065 = 7'h2b == out_payload_1_rob_idx[6:0] ? rob_payload_43_rob_idx : _GEN_6064; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6066 = 7'h2c == out_payload_1_rob_idx[6:0] ? rob_payload_44_rob_idx : _GEN_6065; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6067 = 7'h2d == out_payload_1_rob_idx[6:0] ? rob_payload_45_rob_idx : _GEN_6066; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6068 = 7'h2e == out_payload_1_rob_idx[6:0] ? rob_payload_46_rob_idx : _GEN_6067; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6069 = 7'h2f == out_payload_1_rob_idx[6:0] ? rob_payload_47_rob_idx : _GEN_6068; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6070 = 7'h30 == out_payload_1_rob_idx[6:0] ? rob_payload_48_rob_idx : _GEN_6069; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6071 = 7'h31 == out_payload_1_rob_idx[6:0] ? rob_payload_49_rob_idx : _GEN_6070; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6072 = 7'h32 == out_payload_1_rob_idx[6:0] ? rob_payload_50_rob_idx : _GEN_6071; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6073 = 7'h33 == out_payload_1_rob_idx[6:0] ? rob_payload_51_rob_idx : _GEN_6072; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6074 = 7'h34 == out_payload_1_rob_idx[6:0] ? rob_payload_52_rob_idx : _GEN_6073; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6075 = 7'h35 == out_payload_1_rob_idx[6:0] ? rob_payload_53_rob_idx : _GEN_6074; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6076 = 7'h36 == out_payload_1_rob_idx[6:0] ? rob_payload_54_rob_idx : _GEN_6075; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6077 = 7'h37 == out_payload_1_rob_idx[6:0] ? rob_payload_55_rob_idx : _GEN_6076; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6078 = 7'h38 == out_payload_1_rob_idx[6:0] ? rob_payload_56_rob_idx : _GEN_6077; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6079 = 7'h39 == out_payload_1_rob_idx[6:0] ? rob_payload_57_rob_idx : _GEN_6078; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6080 = 7'h3a == out_payload_1_rob_idx[6:0] ? rob_payload_58_rob_idx : _GEN_6079; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6081 = 7'h3b == out_payload_1_rob_idx[6:0] ? rob_payload_59_rob_idx : _GEN_6080; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6082 = 7'h3c == out_payload_1_rob_idx[6:0] ? rob_payload_60_rob_idx : _GEN_6081; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6083 = 7'h3d == out_payload_1_rob_idx[6:0] ? rob_payload_61_rob_idx : _GEN_6082; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6084 = 7'h3e == out_payload_1_rob_idx[6:0] ? rob_payload_62_rob_idx : _GEN_6083; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6085 = 7'h3f == out_payload_1_rob_idx[6:0] ? rob_payload_63_rob_idx : _GEN_6084; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6086 = 7'h40 == out_payload_1_rob_idx[6:0] ? rob_payload_64_rob_idx : _GEN_6085; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6087 = 7'h41 == out_payload_1_rob_idx[6:0] ? rob_payload_65_rob_idx : _GEN_6086; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6088 = 7'h42 == out_payload_1_rob_idx[6:0] ? rob_payload_66_rob_idx : _GEN_6087; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6089 = 7'h43 == out_payload_1_rob_idx[6:0] ? rob_payload_67_rob_idx : _GEN_6088; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6090 = 7'h44 == out_payload_1_rob_idx[6:0] ? rob_payload_68_rob_idx : _GEN_6089; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6091 = 7'h45 == out_payload_1_rob_idx[6:0] ? rob_payload_69_rob_idx : _GEN_6090; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6092 = 7'h46 == out_payload_1_rob_idx[6:0] ? rob_payload_70_rob_idx : _GEN_6091; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6093 = 7'h47 == out_payload_1_rob_idx[6:0] ? rob_payload_71_rob_idx : _GEN_6092; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6094 = 7'h48 == out_payload_1_rob_idx[6:0] ? rob_payload_72_rob_idx : _GEN_6093; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6095 = 7'h49 == out_payload_1_rob_idx[6:0] ? rob_payload_73_rob_idx : _GEN_6094; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6096 = 7'h4a == out_payload_1_rob_idx[6:0] ? rob_payload_74_rob_idx : _GEN_6095; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6097 = 7'h4b == out_payload_1_rob_idx[6:0] ? rob_payload_75_rob_idx : _GEN_6096; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6098 = 7'h4c == out_payload_1_rob_idx[6:0] ? rob_payload_76_rob_idx : _GEN_6097; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6099 = 7'h4d == out_payload_1_rob_idx[6:0] ? rob_payload_77_rob_idx : _GEN_6098; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6100 = 7'h4e == out_payload_1_rob_idx[6:0] ? rob_payload_78_rob_idx : _GEN_6099; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6101 = 7'h4f == out_payload_1_rob_idx[6:0] ? rob_payload_79_rob_idx : _GEN_6100; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6102 = 7'h50 == out_payload_1_rob_idx[6:0] ? rob_payload_80_rob_idx : _GEN_6101; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6103 = 7'h51 == out_payload_1_rob_idx[6:0] ? rob_payload_81_rob_idx : _GEN_6102; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6104 = 7'h52 == out_payload_1_rob_idx[6:0] ? rob_payload_82_rob_idx : _GEN_6103; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6105 = 7'h53 == out_payload_1_rob_idx[6:0] ? rob_payload_83_rob_idx : _GEN_6104; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6106 = 7'h54 == out_payload_1_rob_idx[6:0] ? rob_payload_84_rob_idx : _GEN_6105; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6107 = 7'h55 == out_payload_1_rob_idx[6:0] ? rob_payload_85_rob_idx : _GEN_6106; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6108 = 7'h56 == out_payload_1_rob_idx[6:0] ? rob_payload_86_rob_idx : _GEN_6107; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6109 = 7'h57 == out_payload_1_rob_idx[6:0] ? rob_payload_87_rob_idx : _GEN_6108; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6110 = 7'h58 == out_payload_1_rob_idx[6:0] ? rob_payload_88_rob_idx : _GEN_6109; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6111 = 7'h59 == out_payload_1_rob_idx[6:0] ? rob_payload_89_rob_idx : _GEN_6110; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6112 = 7'h5a == out_payload_1_rob_idx[6:0] ? rob_payload_90_rob_idx : _GEN_6111; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6113 = 7'h5b == out_payload_1_rob_idx[6:0] ? rob_payload_91_rob_idx : _GEN_6112; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6114 = 7'h5c == out_payload_1_rob_idx[6:0] ? rob_payload_92_rob_idx : _GEN_6113; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6115 = 7'h5d == out_payload_1_rob_idx[6:0] ? rob_payload_93_rob_idx : _GEN_6114; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6116 = 7'h5e == out_payload_1_rob_idx[6:0] ? rob_payload_94_rob_idx : _GEN_6115; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6117 = 7'h5f == out_payload_1_rob_idx[6:0] ? rob_payload_95_rob_idx : _GEN_6116; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6118 = 7'h60 == out_payload_1_rob_idx[6:0] ? rob_payload_96_rob_idx : _GEN_6117; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6119 = 7'h61 == out_payload_1_rob_idx[6:0] ? rob_payload_97_rob_idx : _GEN_6118; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6120 = 7'h62 == out_payload_1_rob_idx[6:0] ? rob_payload_98_rob_idx : _GEN_6119; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6121 = 7'h63 == out_payload_1_rob_idx[6:0] ? rob_payload_99_rob_idx : _GEN_6120; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6122 = 7'h64 == out_payload_1_rob_idx[6:0] ? rob_payload_100_rob_idx : _GEN_6121; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6123 = 7'h65 == out_payload_1_rob_idx[6:0] ? rob_payload_101_rob_idx : _GEN_6122; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6124 = 7'h66 == out_payload_1_rob_idx[6:0] ? rob_payload_102_rob_idx : _GEN_6123; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6125 = 7'h67 == out_payload_1_rob_idx[6:0] ? rob_payload_103_rob_idx : _GEN_6124; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6126 = 7'h68 == out_payload_1_rob_idx[6:0] ? rob_payload_104_rob_idx : _GEN_6125; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6127 = 7'h69 == out_payload_1_rob_idx[6:0] ? rob_payload_105_rob_idx : _GEN_6126; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6128 = 7'h6a == out_payload_1_rob_idx[6:0] ? rob_payload_106_rob_idx : _GEN_6127; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6129 = 7'h6b == out_payload_1_rob_idx[6:0] ? rob_payload_107_rob_idx : _GEN_6128; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6130 = 7'h6c == out_payload_1_rob_idx[6:0] ? rob_payload_108_rob_idx : _GEN_6129; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6131 = 7'h6d == out_payload_1_rob_idx[6:0] ? rob_payload_109_rob_idx : _GEN_6130; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6132 = 7'h6e == out_payload_1_rob_idx[6:0] ? rob_payload_110_rob_idx : _GEN_6131; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6133 = 7'h6f == out_payload_1_rob_idx[6:0] ? rob_payload_111_rob_idx : _GEN_6132; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6134 = 7'h70 == out_payload_1_rob_idx[6:0] ? rob_payload_112_rob_idx : _GEN_6133; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6135 = 7'h71 == out_payload_1_rob_idx[6:0] ? rob_payload_113_rob_idx : _GEN_6134; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6136 = 7'h72 == out_payload_1_rob_idx[6:0] ? rob_payload_114_rob_idx : _GEN_6135; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6137 = 7'h73 == out_payload_1_rob_idx[6:0] ? rob_payload_115_rob_idx : _GEN_6136; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6138 = 7'h74 == out_payload_1_rob_idx[6:0] ? rob_payload_116_rob_idx : _GEN_6137; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6139 = 7'h75 == out_payload_1_rob_idx[6:0] ? rob_payload_117_rob_idx : _GEN_6138; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6140 = 7'h76 == out_payload_1_rob_idx[6:0] ? rob_payload_118_rob_idx : _GEN_6139; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6141 = 7'h77 == out_payload_1_rob_idx[6:0] ? rob_payload_119_rob_idx : _GEN_6140; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6142 = 7'h78 == out_payload_1_rob_idx[6:0] ? rob_payload_120_rob_idx : _GEN_6141; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6143 = 7'h79 == out_payload_1_rob_idx[6:0] ? rob_payload_121_rob_idx : _GEN_6142; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6144 = 7'h7a == out_payload_1_rob_idx[6:0] ? rob_payload_122_rob_idx : _GEN_6143; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6145 = 7'h7b == out_payload_1_rob_idx[6:0] ? rob_payload_123_rob_idx : _GEN_6144; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6146 = 7'h7c == out_payload_1_rob_idx[6:0] ? rob_payload_124_rob_idx : _GEN_6145; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6147 = 7'h7d == out_payload_1_rob_idx[6:0] ? rob_payload_125_rob_idx : _GEN_6146; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6148 = 7'h7e == out_payload_1_rob_idx[6:0] ? rob_payload_126_rob_idx : _GEN_6147; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6149 = 7'h7f == out_payload_1_rob_idx[6:0] ? rob_payload_127_rob_idx : _GEN_6148; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6151 = 7'h1 == out_payload_1_rob_idx[6:0] ? rob_payload_1_flits_fired : rob_payload_0_flits_fired; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6152 = 7'h2 == out_payload_1_rob_idx[6:0] ? rob_payload_2_flits_fired : _GEN_6151; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6153 = 7'h3 == out_payload_1_rob_idx[6:0] ? rob_payload_3_flits_fired : _GEN_6152; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6154 = 7'h4 == out_payload_1_rob_idx[6:0] ? rob_payload_4_flits_fired : _GEN_6153; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6155 = 7'h5 == out_payload_1_rob_idx[6:0] ? rob_payload_5_flits_fired : _GEN_6154; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6156 = 7'h6 == out_payload_1_rob_idx[6:0] ? rob_payload_6_flits_fired : _GEN_6155; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6157 = 7'h7 == out_payload_1_rob_idx[6:0] ? rob_payload_7_flits_fired : _GEN_6156; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6158 = 7'h8 == out_payload_1_rob_idx[6:0] ? rob_payload_8_flits_fired : _GEN_6157; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6159 = 7'h9 == out_payload_1_rob_idx[6:0] ? rob_payload_9_flits_fired : _GEN_6158; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6160 = 7'ha == out_payload_1_rob_idx[6:0] ? rob_payload_10_flits_fired : _GEN_6159; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6161 = 7'hb == out_payload_1_rob_idx[6:0] ? rob_payload_11_flits_fired : _GEN_6160; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6162 = 7'hc == out_payload_1_rob_idx[6:0] ? rob_payload_12_flits_fired : _GEN_6161; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6163 = 7'hd == out_payload_1_rob_idx[6:0] ? rob_payload_13_flits_fired : _GEN_6162; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6164 = 7'he == out_payload_1_rob_idx[6:0] ? rob_payload_14_flits_fired : _GEN_6163; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6165 = 7'hf == out_payload_1_rob_idx[6:0] ? rob_payload_15_flits_fired : _GEN_6164; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6166 = 7'h10 == out_payload_1_rob_idx[6:0] ? rob_payload_16_flits_fired : _GEN_6165; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6167 = 7'h11 == out_payload_1_rob_idx[6:0] ? rob_payload_17_flits_fired : _GEN_6166; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6168 = 7'h12 == out_payload_1_rob_idx[6:0] ? rob_payload_18_flits_fired : _GEN_6167; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6169 = 7'h13 == out_payload_1_rob_idx[6:0] ? rob_payload_19_flits_fired : _GEN_6168; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6170 = 7'h14 == out_payload_1_rob_idx[6:0] ? rob_payload_20_flits_fired : _GEN_6169; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6171 = 7'h15 == out_payload_1_rob_idx[6:0] ? rob_payload_21_flits_fired : _GEN_6170; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6172 = 7'h16 == out_payload_1_rob_idx[6:0] ? rob_payload_22_flits_fired : _GEN_6171; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6173 = 7'h17 == out_payload_1_rob_idx[6:0] ? rob_payload_23_flits_fired : _GEN_6172; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6174 = 7'h18 == out_payload_1_rob_idx[6:0] ? rob_payload_24_flits_fired : _GEN_6173; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6175 = 7'h19 == out_payload_1_rob_idx[6:0] ? rob_payload_25_flits_fired : _GEN_6174; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6176 = 7'h1a == out_payload_1_rob_idx[6:0] ? rob_payload_26_flits_fired : _GEN_6175; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6177 = 7'h1b == out_payload_1_rob_idx[6:0] ? rob_payload_27_flits_fired : _GEN_6176; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6178 = 7'h1c == out_payload_1_rob_idx[6:0] ? rob_payload_28_flits_fired : _GEN_6177; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6179 = 7'h1d == out_payload_1_rob_idx[6:0] ? rob_payload_29_flits_fired : _GEN_6178; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6180 = 7'h1e == out_payload_1_rob_idx[6:0] ? rob_payload_30_flits_fired : _GEN_6179; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6181 = 7'h1f == out_payload_1_rob_idx[6:0] ? rob_payload_31_flits_fired : _GEN_6180; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6182 = 7'h20 == out_payload_1_rob_idx[6:0] ? rob_payload_32_flits_fired : _GEN_6181; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6183 = 7'h21 == out_payload_1_rob_idx[6:0] ? rob_payload_33_flits_fired : _GEN_6182; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6184 = 7'h22 == out_payload_1_rob_idx[6:0] ? rob_payload_34_flits_fired : _GEN_6183; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6185 = 7'h23 == out_payload_1_rob_idx[6:0] ? rob_payload_35_flits_fired : _GEN_6184; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6186 = 7'h24 == out_payload_1_rob_idx[6:0] ? rob_payload_36_flits_fired : _GEN_6185; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6187 = 7'h25 == out_payload_1_rob_idx[6:0] ? rob_payload_37_flits_fired : _GEN_6186; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6188 = 7'h26 == out_payload_1_rob_idx[6:0] ? rob_payload_38_flits_fired : _GEN_6187; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6189 = 7'h27 == out_payload_1_rob_idx[6:0] ? rob_payload_39_flits_fired : _GEN_6188; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6190 = 7'h28 == out_payload_1_rob_idx[6:0] ? rob_payload_40_flits_fired : _GEN_6189; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6191 = 7'h29 == out_payload_1_rob_idx[6:0] ? rob_payload_41_flits_fired : _GEN_6190; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6192 = 7'h2a == out_payload_1_rob_idx[6:0] ? rob_payload_42_flits_fired : _GEN_6191; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6193 = 7'h2b == out_payload_1_rob_idx[6:0] ? rob_payload_43_flits_fired : _GEN_6192; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6194 = 7'h2c == out_payload_1_rob_idx[6:0] ? rob_payload_44_flits_fired : _GEN_6193; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6195 = 7'h2d == out_payload_1_rob_idx[6:0] ? rob_payload_45_flits_fired : _GEN_6194; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6196 = 7'h2e == out_payload_1_rob_idx[6:0] ? rob_payload_46_flits_fired : _GEN_6195; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6197 = 7'h2f == out_payload_1_rob_idx[6:0] ? rob_payload_47_flits_fired : _GEN_6196; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6198 = 7'h30 == out_payload_1_rob_idx[6:0] ? rob_payload_48_flits_fired : _GEN_6197; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6199 = 7'h31 == out_payload_1_rob_idx[6:0] ? rob_payload_49_flits_fired : _GEN_6198; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6200 = 7'h32 == out_payload_1_rob_idx[6:0] ? rob_payload_50_flits_fired : _GEN_6199; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6201 = 7'h33 == out_payload_1_rob_idx[6:0] ? rob_payload_51_flits_fired : _GEN_6200; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6202 = 7'h34 == out_payload_1_rob_idx[6:0] ? rob_payload_52_flits_fired : _GEN_6201; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6203 = 7'h35 == out_payload_1_rob_idx[6:0] ? rob_payload_53_flits_fired : _GEN_6202; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6204 = 7'h36 == out_payload_1_rob_idx[6:0] ? rob_payload_54_flits_fired : _GEN_6203; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6205 = 7'h37 == out_payload_1_rob_idx[6:0] ? rob_payload_55_flits_fired : _GEN_6204; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6206 = 7'h38 == out_payload_1_rob_idx[6:0] ? rob_payload_56_flits_fired : _GEN_6205; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6207 = 7'h39 == out_payload_1_rob_idx[6:0] ? rob_payload_57_flits_fired : _GEN_6206; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6208 = 7'h3a == out_payload_1_rob_idx[6:0] ? rob_payload_58_flits_fired : _GEN_6207; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6209 = 7'h3b == out_payload_1_rob_idx[6:0] ? rob_payload_59_flits_fired : _GEN_6208; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6210 = 7'h3c == out_payload_1_rob_idx[6:0] ? rob_payload_60_flits_fired : _GEN_6209; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6211 = 7'h3d == out_payload_1_rob_idx[6:0] ? rob_payload_61_flits_fired : _GEN_6210; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6212 = 7'h3e == out_payload_1_rob_idx[6:0] ? rob_payload_62_flits_fired : _GEN_6211; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6213 = 7'h3f == out_payload_1_rob_idx[6:0] ? rob_payload_63_flits_fired : _GEN_6212; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6214 = 7'h40 == out_payload_1_rob_idx[6:0] ? rob_payload_64_flits_fired : _GEN_6213; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6215 = 7'h41 == out_payload_1_rob_idx[6:0] ? rob_payload_65_flits_fired : _GEN_6214; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6216 = 7'h42 == out_payload_1_rob_idx[6:0] ? rob_payload_66_flits_fired : _GEN_6215; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6217 = 7'h43 == out_payload_1_rob_idx[6:0] ? rob_payload_67_flits_fired : _GEN_6216; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6218 = 7'h44 == out_payload_1_rob_idx[6:0] ? rob_payload_68_flits_fired : _GEN_6217; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6219 = 7'h45 == out_payload_1_rob_idx[6:0] ? rob_payload_69_flits_fired : _GEN_6218; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6220 = 7'h46 == out_payload_1_rob_idx[6:0] ? rob_payload_70_flits_fired : _GEN_6219; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6221 = 7'h47 == out_payload_1_rob_idx[6:0] ? rob_payload_71_flits_fired : _GEN_6220; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6222 = 7'h48 == out_payload_1_rob_idx[6:0] ? rob_payload_72_flits_fired : _GEN_6221; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6223 = 7'h49 == out_payload_1_rob_idx[6:0] ? rob_payload_73_flits_fired : _GEN_6222; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6224 = 7'h4a == out_payload_1_rob_idx[6:0] ? rob_payload_74_flits_fired : _GEN_6223; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6225 = 7'h4b == out_payload_1_rob_idx[6:0] ? rob_payload_75_flits_fired : _GEN_6224; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6226 = 7'h4c == out_payload_1_rob_idx[6:0] ? rob_payload_76_flits_fired : _GEN_6225; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6227 = 7'h4d == out_payload_1_rob_idx[6:0] ? rob_payload_77_flits_fired : _GEN_6226; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6228 = 7'h4e == out_payload_1_rob_idx[6:0] ? rob_payload_78_flits_fired : _GEN_6227; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6229 = 7'h4f == out_payload_1_rob_idx[6:0] ? rob_payload_79_flits_fired : _GEN_6228; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6230 = 7'h50 == out_payload_1_rob_idx[6:0] ? rob_payload_80_flits_fired : _GEN_6229; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6231 = 7'h51 == out_payload_1_rob_idx[6:0] ? rob_payload_81_flits_fired : _GEN_6230; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6232 = 7'h52 == out_payload_1_rob_idx[6:0] ? rob_payload_82_flits_fired : _GEN_6231; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6233 = 7'h53 == out_payload_1_rob_idx[6:0] ? rob_payload_83_flits_fired : _GEN_6232; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6234 = 7'h54 == out_payload_1_rob_idx[6:0] ? rob_payload_84_flits_fired : _GEN_6233; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6235 = 7'h55 == out_payload_1_rob_idx[6:0] ? rob_payload_85_flits_fired : _GEN_6234; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6236 = 7'h56 == out_payload_1_rob_idx[6:0] ? rob_payload_86_flits_fired : _GEN_6235; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6237 = 7'h57 == out_payload_1_rob_idx[6:0] ? rob_payload_87_flits_fired : _GEN_6236; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6238 = 7'h58 == out_payload_1_rob_idx[6:0] ? rob_payload_88_flits_fired : _GEN_6237; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6239 = 7'h59 == out_payload_1_rob_idx[6:0] ? rob_payload_89_flits_fired : _GEN_6238; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6240 = 7'h5a == out_payload_1_rob_idx[6:0] ? rob_payload_90_flits_fired : _GEN_6239; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6241 = 7'h5b == out_payload_1_rob_idx[6:0] ? rob_payload_91_flits_fired : _GEN_6240; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6242 = 7'h5c == out_payload_1_rob_idx[6:0] ? rob_payload_92_flits_fired : _GEN_6241; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6243 = 7'h5d == out_payload_1_rob_idx[6:0] ? rob_payload_93_flits_fired : _GEN_6242; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6244 = 7'h5e == out_payload_1_rob_idx[6:0] ? rob_payload_94_flits_fired : _GEN_6243; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6245 = 7'h5f == out_payload_1_rob_idx[6:0] ? rob_payload_95_flits_fired : _GEN_6244; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6246 = 7'h60 == out_payload_1_rob_idx[6:0] ? rob_payload_96_flits_fired : _GEN_6245; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6247 = 7'h61 == out_payload_1_rob_idx[6:0] ? rob_payload_97_flits_fired : _GEN_6246; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6248 = 7'h62 == out_payload_1_rob_idx[6:0] ? rob_payload_98_flits_fired : _GEN_6247; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6249 = 7'h63 == out_payload_1_rob_idx[6:0] ? rob_payload_99_flits_fired : _GEN_6248; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6250 = 7'h64 == out_payload_1_rob_idx[6:0] ? rob_payload_100_flits_fired : _GEN_6249; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6251 = 7'h65 == out_payload_1_rob_idx[6:0] ? rob_payload_101_flits_fired : _GEN_6250; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6252 = 7'h66 == out_payload_1_rob_idx[6:0] ? rob_payload_102_flits_fired : _GEN_6251; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6253 = 7'h67 == out_payload_1_rob_idx[6:0] ? rob_payload_103_flits_fired : _GEN_6252; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6254 = 7'h68 == out_payload_1_rob_idx[6:0] ? rob_payload_104_flits_fired : _GEN_6253; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6255 = 7'h69 == out_payload_1_rob_idx[6:0] ? rob_payload_105_flits_fired : _GEN_6254; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6256 = 7'h6a == out_payload_1_rob_idx[6:0] ? rob_payload_106_flits_fired : _GEN_6255; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6257 = 7'h6b == out_payload_1_rob_idx[6:0] ? rob_payload_107_flits_fired : _GEN_6256; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6258 = 7'h6c == out_payload_1_rob_idx[6:0] ? rob_payload_108_flits_fired : _GEN_6257; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6259 = 7'h6d == out_payload_1_rob_idx[6:0] ? rob_payload_109_flits_fired : _GEN_6258; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6260 = 7'h6e == out_payload_1_rob_idx[6:0] ? rob_payload_110_flits_fired : _GEN_6259; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6261 = 7'h6f == out_payload_1_rob_idx[6:0] ? rob_payload_111_flits_fired : _GEN_6260; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6262 = 7'h70 == out_payload_1_rob_idx[6:0] ? rob_payload_112_flits_fired : _GEN_6261; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6263 = 7'h71 == out_payload_1_rob_idx[6:0] ? rob_payload_113_flits_fired : _GEN_6262; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6264 = 7'h72 == out_payload_1_rob_idx[6:0] ? rob_payload_114_flits_fired : _GEN_6263; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6265 = 7'h73 == out_payload_1_rob_idx[6:0] ? rob_payload_115_flits_fired : _GEN_6264; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6266 = 7'h74 == out_payload_1_rob_idx[6:0] ? rob_payload_116_flits_fired : _GEN_6265; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6267 = 7'h75 == out_payload_1_rob_idx[6:0] ? rob_payload_117_flits_fired : _GEN_6266; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6268 = 7'h76 == out_payload_1_rob_idx[6:0] ? rob_payload_118_flits_fired : _GEN_6267; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6269 = 7'h77 == out_payload_1_rob_idx[6:0] ? rob_payload_119_flits_fired : _GEN_6268; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6270 = 7'h78 == out_payload_1_rob_idx[6:0] ? rob_payload_120_flits_fired : _GEN_6269; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6271 = 7'h79 == out_payload_1_rob_idx[6:0] ? rob_payload_121_flits_fired : _GEN_6270; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6272 = 7'h7a == out_payload_1_rob_idx[6:0] ? rob_payload_122_flits_fired : _GEN_6271; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6273 = 7'h7b == out_payload_1_rob_idx[6:0] ? rob_payload_123_flits_fired : _GEN_6272; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6274 = 7'h7c == out_payload_1_rob_idx[6:0] ? rob_payload_124_flits_fired : _GEN_6273; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6275 = 7'h7d == out_payload_1_rob_idx[6:0] ? rob_payload_125_flits_fired : _GEN_6274; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6276 = 7'h7e == out_payload_1_rob_idx[6:0] ? rob_payload_126_flits_fired : _GEN_6275; // @[TestHarness.scala 202:{35,35}]
  wire [15:0] _GEN_6277 = 7'h7f == out_payload_1_rob_idx[6:0] ? rob_payload_127_flits_fired : _GEN_6276; // @[TestHarness.scala 202:{35,35}]
  wire [63:0] _T_95 = {_GEN_6021,_GEN_6149,_GEN_6277}; // @[TestHarness.scala 202:35]
  wire  _GEN_6279 = 7'h1 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_1 : rob_ingress_id_0; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6280 = 7'h2 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_2 : _GEN_6279; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6281 = 7'h3 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_3 : _GEN_6280; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6282 = 7'h4 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_4 : _GEN_6281; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6283 = 7'h5 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_5 : _GEN_6282; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6284 = 7'h6 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_6 : _GEN_6283; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6285 = 7'h7 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_7 : _GEN_6284; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6286 = 7'h8 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_8 : _GEN_6285; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6287 = 7'h9 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_9 : _GEN_6286; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6288 = 7'ha == out_payload_1_rob_idx[6:0] ? rob_ingress_id_10 : _GEN_6287; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6289 = 7'hb == out_payload_1_rob_idx[6:0] ? rob_ingress_id_11 : _GEN_6288; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6290 = 7'hc == out_payload_1_rob_idx[6:0] ? rob_ingress_id_12 : _GEN_6289; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6291 = 7'hd == out_payload_1_rob_idx[6:0] ? rob_ingress_id_13 : _GEN_6290; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6292 = 7'he == out_payload_1_rob_idx[6:0] ? rob_ingress_id_14 : _GEN_6291; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6293 = 7'hf == out_payload_1_rob_idx[6:0] ? rob_ingress_id_15 : _GEN_6292; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6294 = 7'h10 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_16 : _GEN_6293; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6295 = 7'h11 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_17 : _GEN_6294; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6296 = 7'h12 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_18 : _GEN_6295; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6297 = 7'h13 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_19 : _GEN_6296; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6298 = 7'h14 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_20 : _GEN_6297; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6299 = 7'h15 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_21 : _GEN_6298; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6300 = 7'h16 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_22 : _GEN_6299; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6301 = 7'h17 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_23 : _GEN_6300; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6302 = 7'h18 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_24 : _GEN_6301; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6303 = 7'h19 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_25 : _GEN_6302; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6304 = 7'h1a == out_payload_1_rob_idx[6:0] ? rob_ingress_id_26 : _GEN_6303; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6305 = 7'h1b == out_payload_1_rob_idx[6:0] ? rob_ingress_id_27 : _GEN_6304; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6306 = 7'h1c == out_payload_1_rob_idx[6:0] ? rob_ingress_id_28 : _GEN_6305; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6307 = 7'h1d == out_payload_1_rob_idx[6:0] ? rob_ingress_id_29 : _GEN_6306; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6308 = 7'h1e == out_payload_1_rob_idx[6:0] ? rob_ingress_id_30 : _GEN_6307; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6309 = 7'h1f == out_payload_1_rob_idx[6:0] ? rob_ingress_id_31 : _GEN_6308; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6310 = 7'h20 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_32 : _GEN_6309; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6311 = 7'h21 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_33 : _GEN_6310; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6312 = 7'h22 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_34 : _GEN_6311; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6313 = 7'h23 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_35 : _GEN_6312; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6314 = 7'h24 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_36 : _GEN_6313; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6315 = 7'h25 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_37 : _GEN_6314; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6316 = 7'h26 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_38 : _GEN_6315; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6317 = 7'h27 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_39 : _GEN_6316; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6318 = 7'h28 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_40 : _GEN_6317; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6319 = 7'h29 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_41 : _GEN_6318; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6320 = 7'h2a == out_payload_1_rob_idx[6:0] ? rob_ingress_id_42 : _GEN_6319; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6321 = 7'h2b == out_payload_1_rob_idx[6:0] ? rob_ingress_id_43 : _GEN_6320; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6322 = 7'h2c == out_payload_1_rob_idx[6:0] ? rob_ingress_id_44 : _GEN_6321; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6323 = 7'h2d == out_payload_1_rob_idx[6:0] ? rob_ingress_id_45 : _GEN_6322; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6324 = 7'h2e == out_payload_1_rob_idx[6:0] ? rob_ingress_id_46 : _GEN_6323; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6325 = 7'h2f == out_payload_1_rob_idx[6:0] ? rob_ingress_id_47 : _GEN_6324; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6326 = 7'h30 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_48 : _GEN_6325; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6327 = 7'h31 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_49 : _GEN_6326; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6328 = 7'h32 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_50 : _GEN_6327; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6329 = 7'h33 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_51 : _GEN_6328; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6330 = 7'h34 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_52 : _GEN_6329; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6331 = 7'h35 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_53 : _GEN_6330; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6332 = 7'h36 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_54 : _GEN_6331; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6333 = 7'h37 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_55 : _GEN_6332; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6334 = 7'h38 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_56 : _GEN_6333; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6335 = 7'h39 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_57 : _GEN_6334; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6336 = 7'h3a == out_payload_1_rob_idx[6:0] ? rob_ingress_id_58 : _GEN_6335; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6337 = 7'h3b == out_payload_1_rob_idx[6:0] ? rob_ingress_id_59 : _GEN_6336; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6338 = 7'h3c == out_payload_1_rob_idx[6:0] ? rob_ingress_id_60 : _GEN_6337; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6339 = 7'h3d == out_payload_1_rob_idx[6:0] ? rob_ingress_id_61 : _GEN_6338; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6340 = 7'h3e == out_payload_1_rob_idx[6:0] ? rob_ingress_id_62 : _GEN_6339; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6341 = 7'h3f == out_payload_1_rob_idx[6:0] ? rob_ingress_id_63 : _GEN_6340; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6342 = 7'h40 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_64 : _GEN_6341; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6343 = 7'h41 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_65 : _GEN_6342; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6344 = 7'h42 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_66 : _GEN_6343; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6345 = 7'h43 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_67 : _GEN_6344; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6346 = 7'h44 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_68 : _GEN_6345; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6347 = 7'h45 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_69 : _GEN_6346; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6348 = 7'h46 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_70 : _GEN_6347; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6349 = 7'h47 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_71 : _GEN_6348; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6350 = 7'h48 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_72 : _GEN_6349; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6351 = 7'h49 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_73 : _GEN_6350; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6352 = 7'h4a == out_payload_1_rob_idx[6:0] ? rob_ingress_id_74 : _GEN_6351; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6353 = 7'h4b == out_payload_1_rob_idx[6:0] ? rob_ingress_id_75 : _GEN_6352; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6354 = 7'h4c == out_payload_1_rob_idx[6:0] ? rob_ingress_id_76 : _GEN_6353; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6355 = 7'h4d == out_payload_1_rob_idx[6:0] ? rob_ingress_id_77 : _GEN_6354; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6356 = 7'h4e == out_payload_1_rob_idx[6:0] ? rob_ingress_id_78 : _GEN_6355; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6357 = 7'h4f == out_payload_1_rob_idx[6:0] ? rob_ingress_id_79 : _GEN_6356; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6358 = 7'h50 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_80 : _GEN_6357; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6359 = 7'h51 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_81 : _GEN_6358; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6360 = 7'h52 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_82 : _GEN_6359; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6361 = 7'h53 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_83 : _GEN_6360; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6362 = 7'h54 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_84 : _GEN_6361; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6363 = 7'h55 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_85 : _GEN_6362; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6364 = 7'h56 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_86 : _GEN_6363; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6365 = 7'h57 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_87 : _GEN_6364; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6366 = 7'h58 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_88 : _GEN_6365; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6367 = 7'h59 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_89 : _GEN_6366; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6368 = 7'h5a == out_payload_1_rob_idx[6:0] ? rob_ingress_id_90 : _GEN_6367; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6369 = 7'h5b == out_payload_1_rob_idx[6:0] ? rob_ingress_id_91 : _GEN_6368; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6370 = 7'h5c == out_payload_1_rob_idx[6:0] ? rob_ingress_id_92 : _GEN_6369; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6371 = 7'h5d == out_payload_1_rob_idx[6:0] ? rob_ingress_id_93 : _GEN_6370; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6372 = 7'h5e == out_payload_1_rob_idx[6:0] ? rob_ingress_id_94 : _GEN_6371; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6373 = 7'h5f == out_payload_1_rob_idx[6:0] ? rob_ingress_id_95 : _GEN_6372; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6374 = 7'h60 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_96 : _GEN_6373; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6375 = 7'h61 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_97 : _GEN_6374; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6376 = 7'h62 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_98 : _GEN_6375; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6377 = 7'h63 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_99 : _GEN_6376; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6378 = 7'h64 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_100 : _GEN_6377; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6379 = 7'h65 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_101 : _GEN_6378; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6380 = 7'h66 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_102 : _GEN_6379; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6381 = 7'h67 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_103 : _GEN_6380; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6382 = 7'h68 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_104 : _GEN_6381; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6383 = 7'h69 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_105 : _GEN_6382; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6384 = 7'h6a == out_payload_1_rob_idx[6:0] ? rob_ingress_id_106 : _GEN_6383; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6385 = 7'h6b == out_payload_1_rob_idx[6:0] ? rob_ingress_id_107 : _GEN_6384; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6386 = 7'h6c == out_payload_1_rob_idx[6:0] ? rob_ingress_id_108 : _GEN_6385; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6387 = 7'h6d == out_payload_1_rob_idx[6:0] ? rob_ingress_id_109 : _GEN_6386; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6388 = 7'h6e == out_payload_1_rob_idx[6:0] ? rob_ingress_id_110 : _GEN_6387; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6389 = 7'h6f == out_payload_1_rob_idx[6:0] ? rob_ingress_id_111 : _GEN_6388; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6390 = 7'h70 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_112 : _GEN_6389; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6391 = 7'h71 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_113 : _GEN_6390; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6392 = 7'h72 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_114 : _GEN_6391; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6393 = 7'h73 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_115 : _GEN_6392; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6394 = 7'h74 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_116 : _GEN_6393; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6395 = 7'h75 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_117 : _GEN_6394; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6396 = 7'h76 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_118 : _GEN_6395; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6397 = 7'h77 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_119 : _GEN_6396; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6398 = 7'h78 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_120 : _GEN_6397; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6399 = 7'h79 == out_payload_1_rob_idx[6:0] ? rob_ingress_id_121 : _GEN_6398; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6400 = 7'h7a == out_payload_1_rob_idx[6:0] ? rob_ingress_id_122 : _GEN_6399; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6401 = 7'h7b == out_payload_1_rob_idx[6:0] ? rob_ingress_id_123 : _GEN_6400; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6402 = 7'h7c == out_payload_1_rob_idx[6:0] ? rob_ingress_id_124 : _GEN_6401; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6403 = 7'h7d == out_payload_1_rob_idx[6:0] ? rob_ingress_id_125 : _GEN_6402; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6404 = 7'h7e == out_payload_1_rob_idx[6:0] ? rob_ingress_id_126 : _GEN_6403; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6405 = 7'h7f == out_payload_1_rob_idx[6:0] ? rob_ingress_id_127 : _GEN_6404; // @[TestHarness.scala 203:{37,37}]
  wire  _GEN_6407 = 7'h1 == out_payload_1_rob_idx[6:0] ? rob_egress_id_1 : rob_egress_id_0; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6408 = 7'h2 == out_payload_1_rob_idx[6:0] ? rob_egress_id_2 : _GEN_6407; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6409 = 7'h3 == out_payload_1_rob_idx[6:0] ? rob_egress_id_3 : _GEN_6408; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6410 = 7'h4 == out_payload_1_rob_idx[6:0] ? rob_egress_id_4 : _GEN_6409; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6411 = 7'h5 == out_payload_1_rob_idx[6:0] ? rob_egress_id_5 : _GEN_6410; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6412 = 7'h6 == out_payload_1_rob_idx[6:0] ? rob_egress_id_6 : _GEN_6411; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6413 = 7'h7 == out_payload_1_rob_idx[6:0] ? rob_egress_id_7 : _GEN_6412; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6414 = 7'h8 == out_payload_1_rob_idx[6:0] ? rob_egress_id_8 : _GEN_6413; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6415 = 7'h9 == out_payload_1_rob_idx[6:0] ? rob_egress_id_9 : _GEN_6414; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6416 = 7'ha == out_payload_1_rob_idx[6:0] ? rob_egress_id_10 : _GEN_6415; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6417 = 7'hb == out_payload_1_rob_idx[6:0] ? rob_egress_id_11 : _GEN_6416; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6418 = 7'hc == out_payload_1_rob_idx[6:0] ? rob_egress_id_12 : _GEN_6417; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6419 = 7'hd == out_payload_1_rob_idx[6:0] ? rob_egress_id_13 : _GEN_6418; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6420 = 7'he == out_payload_1_rob_idx[6:0] ? rob_egress_id_14 : _GEN_6419; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6421 = 7'hf == out_payload_1_rob_idx[6:0] ? rob_egress_id_15 : _GEN_6420; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6422 = 7'h10 == out_payload_1_rob_idx[6:0] ? rob_egress_id_16 : _GEN_6421; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6423 = 7'h11 == out_payload_1_rob_idx[6:0] ? rob_egress_id_17 : _GEN_6422; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6424 = 7'h12 == out_payload_1_rob_idx[6:0] ? rob_egress_id_18 : _GEN_6423; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6425 = 7'h13 == out_payload_1_rob_idx[6:0] ? rob_egress_id_19 : _GEN_6424; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6426 = 7'h14 == out_payload_1_rob_idx[6:0] ? rob_egress_id_20 : _GEN_6425; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6427 = 7'h15 == out_payload_1_rob_idx[6:0] ? rob_egress_id_21 : _GEN_6426; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6428 = 7'h16 == out_payload_1_rob_idx[6:0] ? rob_egress_id_22 : _GEN_6427; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6429 = 7'h17 == out_payload_1_rob_idx[6:0] ? rob_egress_id_23 : _GEN_6428; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6430 = 7'h18 == out_payload_1_rob_idx[6:0] ? rob_egress_id_24 : _GEN_6429; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6431 = 7'h19 == out_payload_1_rob_idx[6:0] ? rob_egress_id_25 : _GEN_6430; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6432 = 7'h1a == out_payload_1_rob_idx[6:0] ? rob_egress_id_26 : _GEN_6431; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6433 = 7'h1b == out_payload_1_rob_idx[6:0] ? rob_egress_id_27 : _GEN_6432; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6434 = 7'h1c == out_payload_1_rob_idx[6:0] ? rob_egress_id_28 : _GEN_6433; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6435 = 7'h1d == out_payload_1_rob_idx[6:0] ? rob_egress_id_29 : _GEN_6434; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6436 = 7'h1e == out_payload_1_rob_idx[6:0] ? rob_egress_id_30 : _GEN_6435; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6437 = 7'h1f == out_payload_1_rob_idx[6:0] ? rob_egress_id_31 : _GEN_6436; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6438 = 7'h20 == out_payload_1_rob_idx[6:0] ? rob_egress_id_32 : _GEN_6437; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6439 = 7'h21 == out_payload_1_rob_idx[6:0] ? rob_egress_id_33 : _GEN_6438; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6440 = 7'h22 == out_payload_1_rob_idx[6:0] ? rob_egress_id_34 : _GEN_6439; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6441 = 7'h23 == out_payload_1_rob_idx[6:0] ? rob_egress_id_35 : _GEN_6440; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6442 = 7'h24 == out_payload_1_rob_idx[6:0] ? rob_egress_id_36 : _GEN_6441; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6443 = 7'h25 == out_payload_1_rob_idx[6:0] ? rob_egress_id_37 : _GEN_6442; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6444 = 7'h26 == out_payload_1_rob_idx[6:0] ? rob_egress_id_38 : _GEN_6443; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6445 = 7'h27 == out_payload_1_rob_idx[6:0] ? rob_egress_id_39 : _GEN_6444; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6446 = 7'h28 == out_payload_1_rob_idx[6:0] ? rob_egress_id_40 : _GEN_6445; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6447 = 7'h29 == out_payload_1_rob_idx[6:0] ? rob_egress_id_41 : _GEN_6446; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6448 = 7'h2a == out_payload_1_rob_idx[6:0] ? rob_egress_id_42 : _GEN_6447; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6449 = 7'h2b == out_payload_1_rob_idx[6:0] ? rob_egress_id_43 : _GEN_6448; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6450 = 7'h2c == out_payload_1_rob_idx[6:0] ? rob_egress_id_44 : _GEN_6449; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6451 = 7'h2d == out_payload_1_rob_idx[6:0] ? rob_egress_id_45 : _GEN_6450; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6452 = 7'h2e == out_payload_1_rob_idx[6:0] ? rob_egress_id_46 : _GEN_6451; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6453 = 7'h2f == out_payload_1_rob_idx[6:0] ? rob_egress_id_47 : _GEN_6452; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6454 = 7'h30 == out_payload_1_rob_idx[6:0] ? rob_egress_id_48 : _GEN_6453; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6455 = 7'h31 == out_payload_1_rob_idx[6:0] ? rob_egress_id_49 : _GEN_6454; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6456 = 7'h32 == out_payload_1_rob_idx[6:0] ? rob_egress_id_50 : _GEN_6455; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6457 = 7'h33 == out_payload_1_rob_idx[6:0] ? rob_egress_id_51 : _GEN_6456; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6458 = 7'h34 == out_payload_1_rob_idx[6:0] ? rob_egress_id_52 : _GEN_6457; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6459 = 7'h35 == out_payload_1_rob_idx[6:0] ? rob_egress_id_53 : _GEN_6458; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6460 = 7'h36 == out_payload_1_rob_idx[6:0] ? rob_egress_id_54 : _GEN_6459; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6461 = 7'h37 == out_payload_1_rob_idx[6:0] ? rob_egress_id_55 : _GEN_6460; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6462 = 7'h38 == out_payload_1_rob_idx[6:0] ? rob_egress_id_56 : _GEN_6461; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6463 = 7'h39 == out_payload_1_rob_idx[6:0] ? rob_egress_id_57 : _GEN_6462; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6464 = 7'h3a == out_payload_1_rob_idx[6:0] ? rob_egress_id_58 : _GEN_6463; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6465 = 7'h3b == out_payload_1_rob_idx[6:0] ? rob_egress_id_59 : _GEN_6464; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6466 = 7'h3c == out_payload_1_rob_idx[6:0] ? rob_egress_id_60 : _GEN_6465; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6467 = 7'h3d == out_payload_1_rob_idx[6:0] ? rob_egress_id_61 : _GEN_6466; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6468 = 7'h3e == out_payload_1_rob_idx[6:0] ? rob_egress_id_62 : _GEN_6467; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6469 = 7'h3f == out_payload_1_rob_idx[6:0] ? rob_egress_id_63 : _GEN_6468; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6470 = 7'h40 == out_payload_1_rob_idx[6:0] ? rob_egress_id_64 : _GEN_6469; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6471 = 7'h41 == out_payload_1_rob_idx[6:0] ? rob_egress_id_65 : _GEN_6470; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6472 = 7'h42 == out_payload_1_rob_idx[6:0] ? rob_egress_id_66 : _GEN_6471; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6473 = 7'h43 == out_payload_1_rob_idx[6:0] ? rob_egress_id_67 : _GEN_6472; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6474 = 7'h44 == out_payload_1_rob_idx[6:0] ? rob_egress_id_68 : _GEN_6473; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6475 = 7'h45 == out_payload_1_rob_idx[6:0] ? rob_egress_id_69 : _GEN_6474; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6476 = 7'h46 == out_payload_1_rob_idx[6:0] ? rob_egress_id_70 : _GEN_6475; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6477 = 7'h47 == out_payload_1_rob_idx[6:0] ? rob_egress_id_71 : _GEN_6476; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6478 = 7'h48 == out_payload_1_rob_idx[6:0] ? rob_egress_id_72 : _GEN_6477; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6479 = 7'h49 == out_payload_1_rob_idx[6:0] ? rob_egress_id_73 : _GEN_6478; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6480 = 7'h4a == out_payload_1_rob_idx[6:0] ? rob_egress_id_74 : _GEN_6479; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6481 = 7'h4b == out_payload_1_rob_idx[6:0] ? rob_egress_id_75 : _GEN_6480; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6482 = 7'h4c == out_payload_1_rob_idx[6:0] ? rob_egress_id_76 : _GEN_6481; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6483 = 7'h4d == out_payload_1_rob_idx[6:0] ? rob_egress_id_77 : _GEN_6482; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6484 = 7'h4e == out_payload_1_rob_idx[6:0] ? rob_egress_id_78 : _GEN_6483; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6485 = 7'h4f == out_payload_1_rob_idx[6:0] ? rob_egress_id_79 : _GEN_6484; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6486 = 7'h50 == out_payload_1_rob_idx[6:0] ? rob_egress_id_80 : _GEN_6485; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6487 = 7'h51 == out_payload_1_rob_idx[6:0] ? rob_egress_id_81 : _GEN_6486; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6488 = 7'h52 == out_payload_1_rob_idx[6:0] ? rob_egress_id_82 : _GEN_6487; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6489 = 7'h53 == out_payload_1_rob_idx[6:0] ? rob_egress_id_83 : _GEN_6488; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6490 = 7'h54 == out_payload_1_rob_idx[6:0] ? rob_egress_id_84 : _GEN_6489; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6491 = 7'h55 == out_payload_1_rob_idx[6:0] ? rob_egress_id_85 : _GEN_6490; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6492 = 7'h56 == out_payload_1_rob_idx[6:0] ? rob_egress_id_86 : _GEN_6491; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6493 = 7'h57 == out_payload_1_rob_idx[6:0] ? rob_egress_id_87 : _GEN_6492; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6494 = 7'h58 == out_payload_1_rob_idx[6:0] ? rob_egress_id_88 : _GEN_6493; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6495 = 7'h59 == out_payload_1_rob_idx[6:0] ? rob_egress_id_89 : _GEN_6494; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6496 = 7'h5a == out_payload_1_rob_idx[6:0] ? rob_egress_id_90 : _GEN_6495; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6497 = 7'h5b == out_payload_1_rob_idx[6:0] ? rob_egress_id_91 : _GEN_6496; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6498 = 7'h5c == out_payload_1_rob_idx[6:0] ? rob_egress_id_92 : _GEN_6497; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6499 = 7'h5d == out_payload_1_rob_idx[6:0] ? rob_egress_id_93 : _GEN_6498; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6500 = 7'h5e == out_payload_1_rob_idx[6:0] ? rob_egress_id_94 : _GEN_6499; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6501 = 7'h5f == out_payload_1_rob_idx[6:0] ? rob_egress_id_95 : _GEN_6500; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6502 = 7'h60 == out_payload_1_rob_idx[6:0] ? rob_egress_id_96 : _GEN_6501; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6503 = 7'h61 == out_payload_1_rob_idx[6:0] ? rob_egress_id_97 : _GEN_6502; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6504 = 7'h62 == out_payload_1_rob_idx[6:0] ? rob_egress_id_98 : _GEN_6503; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6505 = 7'h63 == out_payload_1_rob_idx[6:0] ? rob_egress_id_99 : _GEN_6504; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6506 = 7'h64 == out_payload_1_rob_idx[6:0] ? rob_egress_id_100 : _GEN_6505; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6507 = 7'h65 == out_payload_1_rob_idx[6:0] ? rob_egress_id_101 : _GEN_6506; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6508 = 7'h66 == out_payload_1_rob_idx[6:0] ? rob_egress_id_102 : _GEN_6507; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6509 = 7'h67 == out_payload_1_rob_idx[6:0] ? rob_egress_id_103 : _GEN_6508; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6510 = 7'h68 == out_payload_1_rob_idx[6:0] ? rob_egress_id_104 : _GEN_6509; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6511 = 7'h69 == out_payload_1_rob_idx[6:0] ? rob_egress_id_105 : _GEN_6510; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6512 = 7'h6a == out_payload_1_rob_idx[6:0] ? rob_egress_id_106 : _GEN_6511; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6513 = 7'h6b == out_payload_1_rob_idx[6:0] ? rob_egress_id_107 : _GEN_6512; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6514 = 7'h6c == out_payload_1_rob_idx[6:0] ? rob_egress_id_108 : _GEN_6513; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6515 = 7'h6d == out_payload_1_rob_idx[6:0] ? rob_egress_id_109 : _GEN_6514; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6516 = 7'h6e == out_payload_1_rob_idx[6:0] ? rob_egress_id_110 : _GEN_6515; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6517 = 7'h6f == out_payload_1_rob_idx[6:0] ? rob_egress_id_111 : _GEN_6516; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6518 = 7'h70 == out_payload_1_rob_idx[6:0] ? rob_egress_id_112 : _GEN_6517; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6519 = 7'h71 == out_payload_1_rob_idx[6:0] ? rob_egress_id_113 : _GEN_6518; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6520 = 7'h72 == out_payload_1_rob_idx[6:0] ? rob_egress_id_114 : _GEN_6519; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6521 = 7'h73 == out_payload_1_rob_idx[6:0] ? rob_egress_id_115 : _GEN_6520; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6522 = 7'h74 == out_payload_1_rob_idx[6:0] ? rob_egress_id_116 : _GEN_6521; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6523 = 7'h75 == out_payload_1_rob_idx[6:0] ? rob_egress_id_117 : _GEN_6522; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6524 = 7'h76 == out_payload_1_rob_idx[6:0] ? rob_egress_id_118 : _GEN_6523; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6525 = 7'h77 == out_payload_1_rob_idx[6:0] ? rob_egress_id_119 : _GEN_6524; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6526 = 7'h78 == out_payload_1_rob_idx[6:0] ? rob_egress_id_120 : _GEN_6525; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6527 = 7'h79 == out_payload_1_rob_idx[6:0] ? rob_egress_id_121 : _GEN_6526; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6528 = 7'h7a == out_payload_1_rob_idx[6:0] ? rob_egress_id_122 : _GEN_6527; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6529 = 7'h7b == out_payload_1_rob_idx[6:0] ? rob_egress_id_123 : _GEN_6528; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6530 = 7'h7c == out_payload_1_rob_idx[6:0] ? rob_egress_id_124 : _GEN_6529; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6531 = 7'h7d == out_payload_1_rob_idx[6:0] ? rob_egress_id_125 : _GEN_6530; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6532 = 7'h7e == out_payload_1_rob_idx[6:0] ? rob_egress_id_126 : _GEN_6531; // @[TestHarness.scala 204:{18,18}]
  wire  _GEN_6533 = 7'h7f == out_payload_1_rob_idx[6:0] ? rob_egress_id_127 : _GEN_6532; // @[TestHarness.scala 204:{18,18}]
  wire [3:0] _GEN_6535 = 7'h1 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_1 : rob_flits_returned_0; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6536 = 7'h2 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_2 : _GEN_6535; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6537 = 7'h3 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_3 : _GEN_6536; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6538 = 7'h4 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_4 : _GEN_6537; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6539 = 7'h5 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_5 : _GEN_6538; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6540 = 7'h6 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_6 : _GEN_6539; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6541 = 7'h7 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_7 : _GEN_6540; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6542 = 7'h8 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_8 : _GEN_6541; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6543 = 7'h9 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_9 : _GEN_6542; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6544 = 7'ha == out_payload_1_rob_idx[6:0] ? rob_flits_returned_10 : _GEN_6543; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6545 = 7'hb == out_payload_1_rob_idx[6:0] ? rob_flits_returned_11 : _GEN_6544; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6546 = 7'hc == out_payload_1_rob_idx[6:0] ? rob_flits_returned_12 : _GEN_6545; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6547 = 7'hd == out_payload_1_rob_idx[6:0] ? rob_flits_returned_13 : _GEN_6546; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6548 = 7'he == out_payload_1_rob_idx[6:0] ? rob_flits_returned_14 : _GEN_6547; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6549 = 7'hf == out_payload_1_rob_idx[6:0] ? rob_flits_returned_15 : _GEN_6548; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6550 = 7'h10 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_16 : _GEN_6549; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6551 = 7'h11 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_17 : _GEN_6550; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6552 = 7'h12 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_18 : _GEN_6551; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6553 = 7'h13 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_19 : _GEN_6552; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6554 = 7'h14 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_20 : _GEN_6553; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6555 = 7'h15 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_21 : _GEN_6554; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6556 = 7'h16 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_22 : _GEN_6555; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6557 = 7'h17 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_23 : _GEN_6556; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6558 = 7'h18 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_24 : _GEN_6557; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6559 = 7'h19 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_25 : _GEN_6558; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6560 = 7'h1a == out_payload_1_rob_idx[6:0] ? rob_flits_returned_26 : _GEN_6559; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6561 = 7'h1b == out_payload_1_rob_idx[6:0] ? rob_flits_returned_27 : _GEN_6560; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6562 = 7'h1c == out_payload_1_rob_idx[6:0] ? rob_flits_returned_28 : _GEN_6561; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6563 = 7'h1d == out_payload_1_rob_idx[6:0] ? rob_flits_returned_29 : _GEN_6562; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6564 = 7'h1e == out_payload_1_rob_idx[6:0] ? rob_flits_returned_30 : _GEN_6563; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6565 = 7'h1f == out_payload_1_rob_idx[6:0] ? rob_flits_returned_31 : _GEN_6564; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6566 = 7'h20 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_32 : _GEN_6565; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6567 = 7'h21 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_33 : _GEN_6566; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6568 = 7'h22 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_34 : _GEN_6567; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6569 = 7'h23 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_35 : _GEN_6568; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6570 = 7'h24 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_36 : _GEN_6569; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6571 = 7'h25 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_37 : _GEN_6570; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6572 = 7'h26 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_38 : _GEN_6571; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6573 = 7'h27 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_39 : _GEN_6572; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6574 = 7'h28 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_40 : _GEN_6573; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6575 = 7'h29 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_41 : _GEN_6574; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6576 = 7'h2a == out_payload_1_rob_idx[6:0] ? rob_flits_returned_42 : _GEN_6575; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6577 = 7'h2b == out_payload_1_rob_idx[6:0] ? rob_flits_returned_43 : _GEN_6576; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6578 = 7'h2c == out_payload_1_rob_idx[6:0] ? rob_flits_returned_44 : _GEN_6577; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6579 = 7'h2d == out_payload_1_rob_idx[6:0] ? rob_flits_returned_45 : _GEN_6578; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6580 = 7'h2e == out_payload_1_rob_idx[6:0] ? rob_flits_returned_46 : _GEN_6579; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6581 = 7'h2f == out_payload_1_rob_idx[6:0] ? rob_flits_returned_47 : _GEN_6580; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6582 = 7'h30 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_48 : _GEN_6581; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6583 = 7'h31 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_49 : _GEN_6582; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6584 = 7'h32 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_50 : _GEN_6583; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6585 = 7'h33 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_51 : _GEN_6584; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6586 = 7'h34 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_52 : _GEN_6585; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6587 = 7'h35 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_53 : _GEN_6586; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6588 = 7'h36 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_54 : _GEN_6587; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6589 = 7'h37 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_55 : _GEN_6588; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6590 = 7'h38 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_56 : _GEN_6589; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6591 = 7'h39 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_57 : _GEN_6590; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6592 = 7'h3a == out_payload_1_rob_idx[6:0] ? rob_flits_returned_58 : _GEN_6591; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6593 = 7'h3b == out_payload_1_rob_idx[6:0] ? rob_flits_returned_59 : _GEN_6592; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6594 = 7'h3c == out_payload_1_rob_idx[6:0] ? rob_flits_returned_60 : _GEN_6593; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6595 = 7'h3d == out_payload_1_rob_idx[6:0] ? rob_flits_returned_61 : _GEN_6594; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6596 = 7'h3e == out_payload_1_rob_idx[6:0] ? rob_flits_returned_62 : _GEN_6595; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6597 = 7'h3f == out_payload_1_rob_idx[6:0] ? rob_flits_returned_63 : _GEN_6596; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6598 = 7'h40 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_64 : _GEN_6597; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6599 = 7'h41 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_65 : _GEN_6598; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6600 = 7'h42 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_66 : _GEN_6599; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6601 = 7'h43 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_67 : _GEN_6600; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6602 = 7'h44 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_68 : _GEN_6601; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6603 = 7'h45 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_69 : _GEN_6602; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6604 = 7'h46 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_70 : _GEN_6603; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6605 = 7'h47 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_71 : _GEN_6604; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6606 = 7'h48 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_72 : _GEN_6605; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6607 = 7'h49 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_73 : _GEN_6606; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6608 = 7'h4a == out_payload_1_rob_idx[6:0] ? rob_flits_returned_74 : _GEN_6607; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6609 = 7'h4b == out_payload_1_rob_idx[6:0] ? rob_flits_returned_75 : _GEN_6608; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6610 = 7'h4c == out_payload_1_rob_idx[6:0] ? rob_flits_returned_76 : _GEN_6609; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6611 = 7'h4d == out_payload_1_rob_idx[6:0] ? rob_flits_returned_77 : _GEN_6610; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6612 = 7'h4e == out_payload_1_rob_idx[6:0] ? rob_flits_returned_78 : _GEN_6611; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6613 = 7'h4f == out_payload_1_rob_idx[6:0] ? rob_flits_returned_79 : _GEN_6612; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6614 = 7'h50 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_80 : _GEN_6613; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6615 = 7'h51 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_81 : _GEN_6614; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6616 = 7'h52 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_82 : _GEN_6615; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6617 = 7'h53 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_83 : _GEN_6616; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6618 = 7'h54 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_84 : _GEN_6617; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6619 = 7'h55 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_85 : _GEN_6618; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6620 = 7'h56 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_86 : _GEN_6619; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6621 = 7'h57 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_87 : _GEN_6620; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6622 = 7'h58 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_88 : _GEN_6621; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6623 = 7'h59 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_89 : _GEN_6622; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6624 = 7'h5a == out_payload_1_rob_idx[6:0] ? rob_flits_returned_90 : _GEN_6623; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6625 = 7'h5b == out_payload_1_rob_idx[6:0] ? rob_flits_returned_91 : _GEN_6624; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6626 = 7'h5c == out_payload_1_rob_idx[6:0] ? rob_flits_returned_92 : _GEN_6625; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6627 = 7'h5d == out_payload_1_rob_idx[6:0] ? rob_flits_returned_93 : _GEN_6626; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6628 = 7'h5e == out_payload_1_rob_idx[6:0] ? rob_flits_returned_94 : _GEN_6627; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6629 = 7'h5f == out_payload_1_rob_idx[6:0] ? rob_flits_returned_95 : _GEN_6628; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6630 = 7'h60 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_96 : _GEN_6629; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6631 = 7'h61 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_97 : _GEN_6630; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6632 = 7'h62 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_98 : _GEN_6631; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6633 = 7'h63 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_99 : _GEN_6632; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6634 = 7'h64 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_100 : _GEN_6633; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6635 = 7'h65 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_101 : _GEN_6634; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6636 = 7'h66 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_102 : _GEN_6635; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6637 = 7'h67 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_103 : _GEN_6636; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6638 = 7'h68 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_104 : _GEN_6637; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6639 = 7'h69 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_105 : _GEN_6638; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6640 = 7'h6a == out_payload_1_rob_idx[6:0] ? rob_flits_returned_106 : _GEN_6639; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6641 = 7'h6b == out_payload_1_rob_idx[6:0] ? rob_flits_returned_107 : _GEN_6640; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6642 = 7'h6c == out_payload_1_rob_idx[6:0] ? rob_flits_returned_108 : _GEN_6641; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6643 = 7'h6d == out_payload_1_rob_idx[6:0] ? rob_flits_returned_109 : _GEN_6642; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6644 = 7'h6e == out_payload_1_rob_idx[6:0] ? rob_flits_returned_110 : _GEN_6643; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6645 = 7'h6f == out_payload_1_rob_idx[6:0] ? rob_flits_returned_111 : _GEN_6644; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6646 = 7'h70 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_112 : _GEN_6645; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6647 = 7'h71 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_113 : _GEN_6646; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6648 = 7'h72 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_114 : _GEN_6647; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6649 = 7'h73 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_115 : _GEN_6648; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6650 = 7'h74 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_116 : _GEN_6649; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6651 = 7'h75 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_117 : _GEN_6650; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6652 = 7'h76 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_118 : _GEN_6651; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6653 = 7'h77 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_119 : _GEN_6652; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6654 = 7'h78 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_120 : _GEN_6653; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6655 = 7'h79 == out_payload_1_rob_idx[6:0] ? rob_flits_returned_121 : _GEN_6654; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6656 = 7'h7a == out_payload_1_rob_idx[6:0] ? rob_flits_returned_122 : _GEN_6655; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6657 = 7'h7b == out_payload_1_rob_idx[6:0] ? rob_flits_returned_123 : _GEN_6656; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6658 = 7'h7c == out_payload_1_rob_idx[6:0] ? rob_flits_returned_124 : _GEN_6657; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6659 = 7'h7d == out_payload_1_rob_idx[6:0] ? rob_flits_returned_125 : _GEN_6658; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6660 = 7'h7e == out_payload_1_rob_idx[6:0] ? rob_flits_returned_126 : _GEN_6659; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6661 = 7'h7f == out_payload_1_rob_idx[6:0] ? rob_flits_returned_127 : _GEN_6660; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6663 = 7'h1 == out_payload_1_rob_idx[6:0] ? rob_n_flits_1 : rob_n_flits_0; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6664 = 7'h2 == out_payload_1_rob_idx[6:0] ? rob_n_flits_2 : _GEN_6663; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6665 = 7'h3 == out_payload_1_rob_idx[6:0] ? rob_n_flits_3 : _GEN_6664; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6666 = 7'h4 == out_payload_1_rob_idx[6:0] ? rob_n_flits_4 : _GEN_6665; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6667 = 7'h5 == out_payload_1_rob_idx[6:0] ? rob_n_flits_5 : _GEN_6666; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6668 = 7'h6 == out_payload_1_rob_idx[6:0] ? rob_n_flits_6 : _GEN_6667; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6669 = 7'h7 == out_payload_1_rob_idx[6:0] ? rob_n_flits_7 : _GEN_6668; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6670 = 7'h8 == out_payload_1_rob_idx[6:0] ? rob_n_flits_8 : _GEN_6669; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6671 = 7'h9 == out_payload_1_rob_idx[6:0] ? rob_n_flits_9 : _GEN_6670; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6672 = 7'ha == out_payload_1_rob_idx[6:0] ? rob_n_flits_10 : _GEN_6671; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6673 = 7'hb == out_payload_1_rob_idx[6:0] ? rob_n_flits_11 : _GEN_6672; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6674 = 7'hc == out_payload_1_rob_idx[6:0] ? rob_n_flits_12 : _GEN_6673; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6675 = 7'hd == out_payload_1_rob_idx[6:0] ? rob_n_flits_13 : _GEN_6674; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6676 = 7'he == out_payload_1_rob_idx[6:0] ? rob_n_flits_14 : _GEN_6675; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6677 = 7'hf == out_payload_1_rob_idx[6:0] ? rob_n_flits_15 : _GEN_6676; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6678 = 7'h10 == out_payload_1_rob_idx[6:0] ? rob_n_flits_16 : _GEN_6677; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6679 = 7'h11 == out_payload_1_rob_idx[6:0] ? rob_n_flits_17 : _GEN_6678; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6680 = 7'h12 == out_payload_1_rob_idx[6:0] ? rob_n_flits_18 : _GEN_6679; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6681 = 7'h13 == out_payload_1_rob_idx[6:0] ? rob_n_flits_19 : _GEN_6680; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6682 = 7'h14 == out_payload_1_rob_idx[6:0] ? rob_n_flits_20 : _GEN_6681; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6683 = 7'h15 == out_payload_1_rob_idx[6:0] ? rob_n_flits_21 : _GEN_6682; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6684 = 7'h16 == out_payload_1_rob_idx[6:0] ? rob_n_flits_22 : _GEN_6683; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6685 = 7'h17 == out_payload_1_rob_idx[6:0] ? rob_n_flits_23 : _GEN_6684; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6686 = 7'h18 == out_payload_1_rob_idx[6:0] ? rob_n_flits_24 : _GEN_6685; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6687 = 7'h19 == out_payload_1_rob_idx[6:0] ? rob_n_flits_25 : _GEN_6686; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6688 = 7'h1a == out_payload_1_rob_idx[6:0] ? rob_n_flits_26 : _GEN_6687; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6689 = 7'h1b == out_payload_1_rob_idx[6:0] ? rob_n_flits_27 : _GEN_6688; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6690 = 7'h1c == out_payload_1_rob_idx[6:0] ? rob_n_flits_28 : _GEN_6689; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6691 = 7'h1d == out_payload_1_rob_idx[6:0] ? rob_n_flits_29 : _GEN_6690; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6692 = 7'h1e == out_payload_1_rob_idx[6:0] ? rob_n_flits_30 : _GEN_6691; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6693 = 7'h1f == out_payload_1_rob_idx[6:0] ? rob_n_flits_31 : _GEN_6692; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6694 = 7'h20 == out_payload_1_rob_idx[6:0] ? rob_n_flits_32 : _GEN_6693; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6695 = 7'h21 == out_payload_1_rob_idx[6:0] ? rob_n_flits_33 : _GEN_6694; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6696 = 7'h22 == out_payload_1_rob_idx[6:0] ? rob_n_flits_34 : _GEN_6695; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6697 = 7'h23 == out_payload_1_rob_idx[6:0] ? rob_n_flits_35 : _GEN_6696; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6698 = 7'h24 == out_payload_1_rob_idx[6:0] ? rob_n_flits_36 : _GEN_6697; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6699 = 7'h25 == out_payload_1_rob_idx[6:0] ? rob_n_flits_37 : _GEN_6698; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6700 = 7'h26 == out_payload_1_rob_idx[6:0] ? rob_n_flits_38 : _GEN_6699; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6701 = 7'h27 == out_payload_1_rob_idx[6:0] ? rob_n_flits_39 : _GEN_6700; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6702 = 7'h28 == out_payload_1_rob_idx[6:0] ? rob_n_flits_40 : _GEN_6701; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6703 = 7'h29 == out_payload_1_rob_idx[6:0] ? rob_n_flits_41 : _GEN_6702; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6704 = 7'h2a == out_payload_1_rob_idx[6:0] ? rob_n_flits_42 : _GEN_6703; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6705 = 7'h2b == out_payload_1_rob_idx[6:0] ? rob_n_flits_43 : _GEN_6704; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6706 = 7'h2c == out_payload_1_rob_idx[6:0] ? rob_n_flits_44 : _GEN_6705; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6707 = 7'h2d == out_payload_1_rob_idx[6:0] ? rob_n_flits_45 : _GEN_6706; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6708 = 7'h2e == out_payload_1_rob_idx[6:0] ? rob_n_flits_46 : _GEN_6707; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6709 = 7'h2f == out_payload_1_rob_idx[6:0] ? rob_n_flits_47 : _GEN_6708; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6710 = 7'h30 == out_payload_1_rob_idx[6:0] ? rob_n_flits_48 : _GEN_6709; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6711 = 7'h31 == out_payload_1_rob_idx[6:0] ? rob_n_flits_49 : _GEN_6710; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6712 = 7'h32 == out_payload_1_rob_idx[6:0] ? rob_n_flits_50 : _GEN_6711; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6713 = 7'h33 == out_payload_1_rob_idx[6:0] ? rob_n_flits_51 : _GEN_6712; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6714 = 7'h34 == out_payload_1_rob_idx[6:0] ? rob_n_flits_52 : _GEN_6713; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6715 = 7'h35 == out_payload_1_rob_idx[6:0] ? rob_n_flits_53 : _GEN_6714; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6716 = 7'h36 == out_payload_1_rob_idx[6:0] ? rob_n_flits_54 : _GEN_6715; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6717 = 7'h37 == out_payload_1_rob_idx[6:0] ? rob_n_flits_55 : _GEN_6716; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6718 = 7'h38 == out_payload_1_rob_idx[6:0] ? rob_n_flits_56 : _GEN_6717; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6719 = 7'h39 == out_payload_1_rob_idx[6:0] ? rob_n_flits_57 : _GEN_6718; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6720 = 7'h3a == out_payload_1_rob_idx[6:0] ? rob_n_flits_58 : _GEN_6719; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6721 = 7'h3b == out_payload_1_rob_idx[6:0] ? rob_n_flits_59 : _GEN_6720; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6722 = 7'h3c == out_payload_1_rob_idx[6:0] ? rob_n_flits_60 : _GEN_6721; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6723 = 7'h3d == out_payload_1_rob_idx[6:0] ? rob_n_flits_61 : _GEN_6722; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6724 = 7'h3e == out_payload_1_rob_idx[6:0] ? rob_n_flits_62 : _GEN_6723; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6725 = 7'h3f == out_payload_1_rob_idx[6:0] ? rob_n_flits_63 : _GEN_6724; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6726 = 7'h40 == out_payload_1_rob_idx[6:0] ? rob_n_flits_64 : _GEN_6725; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6727 = 7'h41 == out_payload_1_rob_idx[6:0] ? rob_n_flits_65 : _GEN_6726; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6728 = 7'h42 == out_payload_1_rob_idx[6:0] ? rob_n_flits_66 : _GEN_6727; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6729 = 7'h43 == out_payload_1_rob_idx[6:0] ? rob_n_flits_67 : _GEN_6728; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6730 = 7'h44 == out_payload_1_rob_idx[6:0] ? rob_n_flits_68 : _GEN_6729; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6731 = 7'h45 == out_payload_1_rob_idx[6:0] ? rob_n_flits_69 : _GEN_6730; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6732 = 7'h46 == out_payload_1_rob_idx[6:0] ? rob_n_flits_70 : _GEN_6731; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6733 = 7'h47 == out_payload_1_rob_idx[6:0] ? rob_n_flits_71 : _GEN_6732; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6734 = 7'h48 == out_payload_1_rob_idx[6:0] ? rob_n_flits_72 : _GEN_6733; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6735 = 7'h49 == out_payload_1_rob_idx[6:0] ? rob_n_flits_73 : _GEN_6734; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6736 = 7'h4a == out_payload_1_rob_idx[6:0] ? rob_n_flits_74 : _GEN_6735; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6737 = 7'h4b == out_payload_1_rob_idx[6:0] ? rob_n_flits_75 : _GEN_6736; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6738 = 7'h4c == out_payload_1_rob_idx[6:0] ? rob_n_flits_76 : _GEN_6737; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6739 = 7'h4d == out_payload_1_rob_idx[6:0] ? rob_n_flits_77 : _GEN_6738; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6740 = 7'h4e == out_payload_1_rob_idx[6:0] ? rob_n_flits_78 : _GEN_6739; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6741 = 7'h4f == out_payload_1_rob_idx[6:0] ? rob_n_flits_79 : _GEN_6740; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6742 = 7'h50 == out_payload_1_rob_idx[6:0] ? rob_n_flits_80 : _GEN_6741; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6743 = 7'h51 == out_payload_1_rob_idx[6:0] ? rob_n_flits_81 : _GEN_6742; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6744 = 7'h52 == out_payload_1_rob_idx[6:0] ? rob_n_flits_82 : _GEN_6743; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6745 = 7'h53 == out_payload_1_rob_idx[6:0] ? rob_n_flits_83 : _GEN_6744; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6746 = 7'h54 == out_payload_1_rob_idx[6:0] ? rob_n_flits_84 : _GEN_6745; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6747 = 7'h55 == out_payload_1_rob_idx[6:0] ? rob_n_flits_85 : _GEN_6746; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6748 = 7'h56 == out_payload_1_rob_idx[6:0] ? rob_n_flits_86 : _GEN_6747; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6749 = 7'h57 == out_payload_1_rob_idx[6:0] ? rob_n_flits_87 : _GEN_6748; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6750 = 7'h58 == out_payload_1_rob_idx[6:0] ? rob_n_flits_88 : _GEN_6749; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6751 = 7'h59 == out_payload_1_rob_idx[6:0] ? rob_n_flits_89 : _GEN_6750; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6752 = 7'h5a == out_payload_1_rob_idx[6:0] ? rob_n_flits_90 : _GEN_6751; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6753 = 7'h5b == out_payload_1_rob_idx[6:0] ? rob_n_flits_91 : _GEN_6752; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6754 = 7'h5c == out_payload_1_rob_idx[6:0] ? rob_n_flits_92 : _GEN_6753; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6755 = 7'h5d == out_payload_1_rob_idx[6:0] ? rob_n_flits_93 : _GEN_6754; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6756 = 7'h5e == out_payload_1_rob_idx[6:0] ? rob_n_flits_94 : _GEN_6755; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6757 = 7'h5f == out_payload_1_rob_idx[6:0] ? rob_n_flits_95 : _GEN_6756; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6758 = 7'h60 == out_payload_1_rob_idx[6:0] ? rob_n_flits_96 : _GEN_6757; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6759 = 7'h61 == out_payload_1_rob_idx[6:0] ? rob_n_flits_97 : _GEN_6758; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6760 = 7'h62 == out_payload_1_rob_idx[6:0] ? rob_n_flits_98 : _GEN_6759; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6761 = 7'h63 == out_payload_1_rob_idx[6:0] ? rob_n_flits_99 : _GEN_6760; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6762 = 7'h64 == out_payload_1_rob_idx[6:0] ? rob_n_flits_100 : _GEN_6761; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6763 = 7'h65 == out_payload_1_rob_idx[6:0] ? rob_n_flits_101 : _GEN_6762; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6764 = 7'h66 == out_payload_1_rob_idx[6:0] ? rob_n_flits_102 : _GEN_6763; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6765 = 7'h67 == out_payload_1_rob_idx[6:0] ? rob_n_flits_103 : _GEN_6764; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6766 = 7'h68 == out_payload_1_rob_idx[6:0] ? rob_n_flits_104 : _GEN_6765; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6767 = 7'h69 == out_payload_1_rob_idx[6:0] ? rob_n_flits_105 : _GEN_6766; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6768 = 7'h6a == out_payload_1_rob_idx[6:0] ? rob_n_flits_106 : _GEN_6767; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6769 = 7'h6b == out_payload_1_rob_idx[6:0] ? rob_n_flits_107 : _GEN_6768; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6770 = 7'h6c == out_payload_1_rob_idx[6:0] ? rob_n_flits_108 : _GEN_6769; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6771 = 7'h6d == out_payload_1_rob_idx[6:0] ? rob_n_flits_109 : _GEN_6770; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6772 = 7'h6e == out_payload_1_rob_idx[6:0] ? rob_n_flits_110 : _GEN_6771; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6773 = 7'h6f == out_payload_1_rob_idx[6:0] ? rob_n_flits_111 : _GEN_6772; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6774 = 7'h70 == out_payload_1_rob_idx[6:0] ? rob_n_flits_112 : _GEN_6773; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6775 = 7'h71 == out_payload_1_rob_idx[6:0] ? rob_n_flits_113 : _GEN_6774; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6776 = 7'h72 == out_payload_1_rob_idx[6:0] ? rob_n_flits_114 : _GEN_6775; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6777 = 7'h73 == out_payload_1_rob_idx[6:0] ? rob_n_flits_115 : _GEN_6776; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6778 = 7'h74 == out_payload_1_rob_idx[6:0] ? rob_n_flits_116 : _GEN_6777; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6779 = 7'h75 == out_payload_1_rob_idx[6:0] ? rob_n_flits_117 : _GEN_6778; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6780 = 7'h76 == out_payload_1_rob_idx[6:0] ? rob_n_flits_118 : _GEN_6779; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6781 = 7'h77 == out_payload_1_rob_idx[6:0] ? rob_n_flits_119 : _GEN_6780; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6782 = 7'h78 == out_payload_1_rob_idx[6:0] ? rob_n_flits_120 : _GEN_6781; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6783 = 7'h79 == out_payload_1_rob_idx[6:0] ? rob_n_flits_121 : _GEN_6782; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6784 = 7'h7a == out_payload_1_rob_idx[6:0] ? rob_n_flits_122 : _GEN_6783; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6785 = 7'h7b == out_payload_1_rob_idx[6:0] ? rob_n_flits_123 : _GEN_6784; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6786 = 7'h7c == out_payload_1_rob_idx[6:0] ? rob_n_flits_124 : _GEN_6785; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6787 = 7'h7d == out_payload_1_rob_idx[6:0] ? rob_n_flits_125 : _GEN_6786; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6788 = 7'h7e == out_payload_1_rob_idx[6:0] ? rob_n_flits_126 : _GEN_6787; // @[TestHarness.scala 205:{42,42}]
  wire [3:0] _GEN_6789 = 7'h7f == out_payload_1_rob_idx[6:0] ? rob_n_flits_127 : _GEN_6788; // @[TestHarness.scala 205:{42,42}]
  wire [15:0] _GEN_7820 = {{9'd0}, packet_rob_idx_1}; // @[TestHarness.scala 206:61]
  wire  _T_123 = io_from_noc_1_flit_bits_head & enable_print_latency; // @[TestHarness.scala 208:30]
  wire [3:0] _rob_flits_returned_T_5 = _GEN_6661 + 4'h1; // @[TestHarness.scala 213:66]
  wire [15:0] _rob_payload_flits_fired_T_5 = _GEN_6277 + 16'h1; // @[TestHarness.scala 214:76]
  wire  _GEN_7430 = io_from_noc_1_flit_bits_head | packet_valid_1; // @[TestHarness.scala 196:31 215:{31,46}]
  wire [15:0] _GEN_7431 = io_from_noc_1_flit_bits_head ? out_payload_1_rob_idx : {{9'd0}, packet_rob_idx_1}; // @[TestHarness.scala 197:29 215:{31,72}]
  wire [15:0] _GEN_7690 = _T_131 ? _GEN_7431 : {{9'd0}, packet_rob_idx_1}; // @[TestHarness.scala 199:26 197:29]
  wire [127:0] _rob_valids_T = rob_valids | rob_allocs; // @[TestHarness.scala 222:29]
  wire [65535:0] _rob_valids_T_1 = ~rob_frees; // @[TestHarness.scala 222:45]
  wire [65535:0] _GEN_7821 = {{65408'd0}, _rob_valids_T}; // @[TestHarness.scala 222:43]
  wire [65535:0] _rob_valids_T_2 = _GEN_7821 & _rob_valids_T_1; // @[TestHarness.scala 222:43]
  wire [1:0] _flits_T_2 = _T_84 + _T_131; // @[TestHarness.scala 224:66]
  wire [31:0] _GEN_7822 = {{30'd0}, _flits_T_2}; // @[TestHarness.scala 224:18]
  wire [31:0] _flits_T_4 = flits + _GEN_7822; // @[TestHarness.scala 224:18]
  wire  tx_fire_0 = igen_io_fire; // @[TestHarness.scala 169:21 186:18]
  wire  tx_fire_1 = igen_1_io_fire; // @[TestHarness.scala 169:21 186:18]
  wire [1:0] _txs_T = tx_fire_0 + tx_fire_1; // @[Bitwise.scala 51:90]
  wire [31:0] _GEN_7823 = {{30'd0}, _txs_T}; // @[TestHarness.scala 225:14]
  wire [31:0] _txs_T_3 = txs + _GEN_7823; // @[TestHarness.scala 225:14]
  wire [63:0] _T_136 = _rob_tscs_T_25 - rob_tscs_0; // @[TestHarness.scala 229:18]
  wire [63:0] _T_143 = _rob_tscs_T_25 - rob_tscs_1; // @[TestHarness.scala 229:18]
  wire [63:0] _T_150 = _rob_tscs_T_25 - rob_tscs_2; // @[TestHarness.scala 229:18]
  wire [63:0] _T_157 = _rob_tscs_T_25 - rob_tscs_3; // @[TestHarness.scala 229:18]
  wire [63:0] _T_164 = _rob_tscs_T_25 - rob_tscs_4; // @[TestHarness.scala 229:18]
  wire [63:0] _T_171 = _rob_tscs_T_25 - rob_tscs_5; // @[TestHarness.scala 229:18]
  wire [63:0] _T_178 = _rob_tscs_T_25 - rob_tscs_6; // @[TestHarness.scala 229:18]
  wire [63:0] _T_185 = _rob_tscs_T_25 - rob_tscs_7; // @[TestHarness.scala 229:18]
  wire [63:0] _T_192 = _rob_tscs_T_25 - rob_tscs_8; // @[TestHarness.scala 229:18]
  wire [63:0] _T_199 = _rob_tscs_T_25 - rob_tscs_9; // @[TestHarness.scala 229:18]
  wire [63:0] _T_206 = _rob_tscs_T_25 - rob_tscs_10; // @[TestHarness.scala 229:18]
  wire [63:0] _T_213 = _rob_tscs_T_25 - rob_tscs_11; // @[TestHarness.scala 229:18]
  wire [63:0] _T_220 = _rob_tscs_T_25 - rob_tscs_12; // @[TestHarness.scala 229:18]
  wire [63:0] _T_227 = _rob_tscs_T_25 - rob_tscs_13; // @[TestHarness.scala 229:18]
  wire [63:0] _T_234 = _rob_tscs_T_25 - rob_tscs_14; // @[TestHarness.scala 229:18]
  wire [63:0] _T_241 = _rob_tscs_T_25 - rob_tscs_15; // @[TestHarness.scala 229:18]
  wire [63:0] _T_248 = _rob_tscs_T_25 - rob_tscs_16; // @[TestHarness.scala 229:18]
  wire [63:0] _T_255 = _rob_tscs_T_25 - rob_tscs_17; // @[TestHarness.scala 229:18]
  wire [63:0] _T_262 = _rob_tscs_T_25 - rob_tscs_18; // @[TestHarness.scala 229:18]
  wire [63:0] _T_269 = _rob_tscs_T_25 - rob_tscs_19; // @[TestHarness.scala 229:18]
  wire [63:0] _T_276 = _rob_tscs_T_25 - rob_tscs_20; // @[TestHarness.scala 229:18]
  wire [63:0] _T_283 = _rob_tscs_T_25 - rob_tscs_21; // @[TestHarness.scala 229:18]
  wire [63:0] _T_290 = _rob_tscs_T_25 - rob_tscs_22; // @[TestHarness.scala 229:18]
  wire [63:0] _T_297 = _rob_tscs_T_25 - rob_tscs_23; // @[TestHarness.scala 229:18]
  wire [63:0] _T_304 = _rob_tscs_T_25 - rob_tscs_24; // @[TestHarness.scala 229:18]
  wire [63:0] _T_311 = _rob_tscs_T_25 - rob_tscs_25; // @[TestHarness.scala 229:18]
  wire [63:0] _T_318 = _rob_tscs_T_25 - rob_tscs_26; // @[TestHarness.scala 229:18]
  wire [63:0] _T_325 = _rob_tscs_T_25 - rob_tscs_27; // @[TestHarness.scala 229:18]
  wire [63:0] _T_332 = _rob_tscs_T_25 - rob_tscs_28; // @[TestHarness.scala 229:18]
  wire [63:0] _T_339 = _rob_tscs_T_25 - rob_tscs_29; // @[TestHarness.scala 229:18]
  wire [63:0] _T_346 = _rob_tscs_T_25 - rob_tscs_30; // @[TestHarness.scala 229:18]
  wire [63:0] _T_353 = _rob_tscs_T_25 - rob_tscs_31; // @[TestHarness.scala 229:18]
  wire [63:0] _T_360 = _rob_tscs_T_25 - rob_tscs_32; // @[TestHarness.scala 229:18]
  wire [63:0] _T_367 = _rob_tscs_T_25 - rob_tscs_33; // @[TestHarness.scala 229:18]
  wire [63:0] _T_374 = _rob_tscs_T_25 - rob_tscs_34; // @[TestHarness.scala 229:18]
  wire [63:0] _T_381 = _rob_tscs_T_25 - rob_tscs_35; // @[TestHarness.scala 229:18]
  wire [63:0] _T_388 = _rob_tscs_T_25 - rob_tscs_36; // @[TestHarness.scala 229:18]
  wire [63:0] _T_395 = _rob_tscs_T_25 - rob_tscs_37; // @[TestHarness.scala 229:18]
  wire [63:0] _T_402 = _rob_tscs_T_25 - rob_tscs_38; // @[TestHarness.scala 229:18]
  wire [63:0] _T_409 = _rob_tscs_T_25 - rob_tscs_39; // @[TestHarness.scala 229:18]
  wire [63:0] _T_416 = _rob_tscs_T_25 - rob_tscs_40; // @[TestHarness.scala 229:18]
  wire [63:0] _T_423 = _rob_tscs_T_25 - rob_tscs_41; // @[TestHarness.scala 229:18]
  wire [63:0] _T_430 = _rob_tscs_T_25 - rob_tscs_42; // @[TestHarness.scala 229:18]
  wire [63:0] _T_437 = _rob_tscs_T_25 - rob_tscs_43; // @[TestHarness.scala 229:18]
  wire [63:0] _T_444 = _rob_tscs_T_25 - rob_tscs_44; // @[TestHarness.scala 229:18]
  wire [63:0] _T_451 = _rob_tscs_T_25 - rob_tscs_45; // @[TestHarness.scala 229:18]
  wire [63:0] _T_458 = _rob_tscs_T_25 - rob_tscs_46; // @[TestHarness.scala 229:18]
  wire [63:0] _T_465 = _rob_tscs_T_25 - rob_tscs_47; // @[TestHarness.scala 229:18]
  wire [63:0] _T_472 = _rob_tscs_T_25 - rob_tscs_48; // @[TestHarness.scala 229:18]
  wire [63:0] _T_479 = _rob_tscs_T_25 - rob_tscs_49; // @[TestHarness.scala 229:18]
  wire [63:0] _T_486 = _rob_tscs_T_25 - rob_tscs_50; // @[TestHarness.scala 229:18]
  wire [63:0] _T_493 = _rob_tscs_T_25 - rob_tscs_51; // @[TestHarness.scala 229:18]
  wire [63:0] _T_500 = _rob_tscs_T_25 - rob_tscs_52; // @[TestHarness.scala 229:18]
  wire [63:0] _T_507 = _rob_tscs_T_25 - rob_tscs_53; // @[TestHarness.scala 229:18]
  wire [63:0] _T_514 = _rob_tscs_T_25 - rob_tscs_54; // @[TestHarness.scala 229:18]
  wire [63:0] _T_521 = _rob_tscs_T_25 - rob_tscs_55; // @[TestHarness.scala 229:18]
  wire [63:0] _T_528 = _rob_tscs_T_25 - rob_tscs_56; // @[TestHarness.scala 229:18]
  wire [63:0] _T_535 = _rob_tscs_T_25 - rob_tscs_57; // @[TestHarness.scala 229:18]
  wire [63:0] _T_542 = _rob_tscs_T_25 - rob_tscs_58; // @[TestHarness.scala 229:18]
  wire [63:0] _T_549 = _rob_tscs_T_25 - rob_tscs_59; // @[TestHarness.scala 229:18]
  wire [63:0] _T_556 = _rob_tscs_T_25 - rob_tscs_60; // @[TestHarness.scala 229:18]
  wire [63:0] _T_563 = _rob_tscs_T_25 - rob_tscs_61; // @[TestHarness.scala 229:18]
  wire [63:0] _T_570 = _rob_tscs_T_25 - rob_tscs_62; // @[TestHarness.scala 229:18]
  wire [63:0] _T_577 = _rob_tscs_T_25 - rob_tscs_63; // @[TestHarness.scala 229:18]
  wire [63:0] _T_584 = _rob_tscs_T_25 - rob_tscs_64; // @[TestHarness.scala 229:18]
  wire [63:0] _T_591 = _rob_tscs_T_25 - rob_tscs_65; // @[TestHarness.scala 229:18]
  wire [63:0] _T_598 = _rob_tscs_T_25 - rob_tscs_66; // @[TestHarness.scala 229:18]
  wire [63:0] _T_605 = _rob_tscs_T_25 - rob_tscs_67; // @[TestHarness.scala 229:18]
  wire [63:0] _T_612 = _rob_tscs_T_25 - rob_tscs_68; // @[TestHarness.scala 229:18]
  wire [63:0] _T_619 = _rob_tscs_T_25 - rob_tscs_69; // @[TestHarness.scala 229:18]
  wire [63:0] _T_626 = _rob_tscs_T_25 - rob_tscs_70; // @[TestHarness.scala 229:18]
  wire [63:0] _T_633 = _rob_tscs_T_25 - rob_tscs_71; // @[TestHarness.scala 229:18]
  wire [63:0] _T_640 = _rob_tscs_T_25 - rob_tscs_72; // @[TestHarness.scala 229:18]
  wire [63:0] _T_647 = _rob_tscs_T_25 - rob_tscs_73; // @[TestHarness.scala 229:18]
  wire [63:0] _T_654 = _rob_tscs_T_25 - rob_tscs_74; // @[TestHarness.scala 229:18]
  wire [63:0] _T_661 = _rob_tscs_T_25 - rob_tscs_75; // @[TestHarness.scala 229:18]
  wire [63:0] _T_668 = _rob_tscs_T_25 - rob_tscs_76; // @[TestHarness.scala 229:18]
  wire [63:0] _T_675 = _rob_tscs_T_25 - rob_tscs_77; // @[TestHarness.scala 229:18]
  wire [63:0] _T_682 = _rob_tscs_T_25 - rob_tscs_78; // @[TestHarness.scala 229:18]
  wire [63:0] _T_689 = _rob_tscs_T_25 - rob_tscs_79; // @[TestHarness.scala 229:18]
  wire [63:0] _T_696 = _rob_tscs_T_25 - rob_tscs_80; // @[TestHarness.scala 229:18]
  wire [63:0] _T_703 = _rob_tscs_T_25 - rob_tscs_81; // @[TestHarness.scala 229:18]
  wire [63:0] _T_710 = _rob_tscs_T_25 - rob_tscs_82; // @[TestHarness.scala 229:18]
  wire [63:0] _T_717 = _rob_tscs_T_25 - rob_tscs_83; // @[TestHarness.scala 229:18]
  wire [63:0] _T_724 = _rob_tscs_T_25 - rob_tscs_84; // @[TestHarness.scala 229:18]
  wire [63:0] _T_731 = _rob_tscs_T_25 - rob_tscs_85; // @[TestHarness.scala 229:18]
  wire [63:0] _T_738 = _rob_tscs_T_25 - rob_tscs_86; // @[TestHarness.scala 229:18]
  wire [63:0] _T_745 = _rob_tscs_T_25 - rob_tscs_87; // @[TestHarness.scala 229:18]
  wire [63:0] _T_752 = _rob_tscs_T_25 - rob_tscs_88; // @[TestHarness.scala 229:18]
  wire [63:0] _T_759 = _rob_tscs_T_25 - rob_tscs_89; // @[TestHarness.scala 229:18]
  wire [63:0] _T_766 = _rob_tscs_T_25 - rob_tscs_90; // @[TestHarness.scala 229:18]
  wire [63:0] _T_773 = _rob_tscs_T_25 - rob_tscs_91; // @[TestHarness.scala 229:18]
  wire [63:0] _T_780 = _rob_tscs_T_25 - rob_tscs_92; // @[TestHarness.scala 229:18]
  wire [63:0] _T_787 = _rob_tscs_T_25 - rob_tscs_93; // @[TestHarness.scala 229:18]
  wire [63:0] _T_794 = _rob_tscs_T_25 - rob_tscs_94; // @[TestHarness.scala 229:18]
  wire [63:0] _T_801 = _rob_tscs_T_25 - rob_tscs_95; // @[TestHarness.scala 229:18]
  wire [63:0] _T_808 = _rob_tscs_T_25 - rob_tscs_96; // @[TestHarness.scala 229:18]
  wire [63:0] _T_815 = _rob_tscs_T_25 - rob_tscs_97; // @[TestHarness.scala 229:18]
  wire [63:0] _T_822 = _rob_tscs_T_25 - rob_tscs_98; // @[TestHarness.scala 229:18]
  wire [63:0] _T_829 = _rob_tscs_T_25 - rob_tscs_99; // @[TestHarness.scala 229:18]
  wire [63:0] _T_836 = _rob_tscs_T_25 - rob_tscs_100; // @[TestHarness.scala 229:18]
  wire [63:0] _T_843 = _rob_tscs_T_25 - rob_tscs_101; // @[TestHarness.scala 229:18]
  wire [63:0] _T_850 = _rob_tscs_T_25 - rob_tscs_102; // @[TestHarness.scala 229:18]
  wire [63:0] _T_857 = _rob_tscs_T_25 - rob_tscs_103; // @[TestHarness.scala 229:18]
  wire [63:0] _T_864 = _rob_tscs_T_25 - rob_tscs_104; // @[TestHarness.scala 229:18]
  wire [63:0] _T_871 = _rob_tscs_T_25 - rob_tscs_105; // @[TestHarness.scala 229:18]
  wire [63:0] _T_878 = _rob_tscs_T_25 - rob_tscs_106; // @[TestHarness.scala 229:18]
  wire [63:0] _T_885 = _rob_tscs_T_25 - rob_tscs_107; // @[TestHarness.scala 229:18]
  wire [63:0] _T_892 = _rob_tscs_T_25 - rob_tscs_108; // @[TestHarness.scala 229:18]
  wire [63:0] _T_899 = _rob_tscs_T_25 - rob_tscs_109; // @[TestHarness.scala 229:18]
  wire [63:0] _T_906 = _rob_tscs_T_25 - rob_tscs_110; // @[TestHarness.scala 229:18]
  wire [63:0] _T_913 = _rob_tscs_T_25 - rob_tscs_111; // @[TestHarness.scala 229:18]
  wire [63:0] _T_920 = _rob_tscs_T_25 - rob_tscs_112; // @[TestHarness.scala 229:18]
  wire [63:0] _T_927 = _rob_tscs_T_25 - rob_tscs_113; // @[TestHarness.scala 229:18]
  wire [63:0] _T_934 = _rob_tscs_T_25 - rob_tscs_114; // @[TestHarness.scala 229:18]
  wire [63:0] _T_941 = _rob_tscs_T_25 - rob_tscs_115; // @[TestHarness.scala 229:18]
  wire [63:0] _T_948 = _rob_tscs_T_25 - rob_tscs_116; // @[TestHarness.scala 229:18]
  wire [63:0] _T_955 = _rob_tscs_T_25 - rob_tscs_117; // @[TestHarness.scala 229:18]
  wire [63:0] _T_962 = _rob_tscs_T_25 - rob_tscs_118; // @[TestHarness.scala 229:18]
  wire [63:0] _T_969 = _rob_tscs_T_25 - rob_tscs_119; // @[TestHarness.scala 229:18]
  wire [63:0] _T_976 = _rob_tscs_T_25 - rob_tscs_120; // @[TestHarness.scala 229:18]
  wire [63:0] _T_983 = _rob_tscs_T_25 - rob_tscs_121; // @[TestHarness.scala 229:18]
  wire [63:0] _T_990 = _rob_tscs_T_25 - rob_tscs_122; // @[TestHarness.scala 229:18]
  wire [63:0] _T_997 = _rob_tscs_T_25 - rob_tscs_123; // @[TestHarness.scala 229:18]
  wire [63:0] _T_1004 = _rob_tscs_T_25 - rob_tscs_124; // @[TestHarness.scala 229:18]
  wire [63:0] _T_1011 = _rob_tscs_T_25 - rob_tscs_125; // @[TestHarness.scala 229:18]
  wire [63:0] _T_1018 = _rob_tscs_T_25 - rob_tscs_126; // @[TestHarness.scala 229:18]
  wire [63:0] _T_1025 = _rob_tscs_T_25 - rob_tscs_127; // @[TestHarness.scala 229:18]
  wire [65535:0] _GEN_7952 = reset ? 65536'h0 : _rob_valids_T_2; // @[TestHarness.scala 156:{27,27} 222:14]
  wire  _GEN_7953 = _T_84 & _T_3; // @[TestHarness.scala 201:13]
  wire  _GEN_7960 = _T_131 & _T_3; // @[TestHarness.scala 201:13]
  InputGen igen ( // @[TestHarness.scala 171:22]
    .clock(igen_clock),
    .reset(igen_reset),
    .io_out_ready(igen_io_out_ready),
    .io_out_valid(igen_io_out_valid),
    .io_out_bits_head(igen_io_out_bits_head),
    .io_out_bits_tail(igen_io_out_bits_tail),
    .io_out_bits_payload(igen_io_out_bits_payload),
    .io_out_bits_egress_id(igen_io_out_bits_egress_id),
    .io_rob_ready(igen_io_rob_ready),
    .io_rob_idx(igen_io_rob_idx),
    .io_tsc(igen_io_tsc),
    .io_fire(igen_io_fire),
    .io_n_flits(igen_io_n_flits)
  );
  Queue_26 io_to_noc_0_flit_q ( // @[Decoupled.scala 375:21]
    .clock(io_to_noc_0_flit_q_clock),
    .reset(io_to_noc_0_flit_q_reset),
    .io_enq_ready(io_to_noc_0_flit_q_io_enq_ready),
    .io_enq_valid(io_to_noc_0_flit_q_io_enq_valid),
    .io_enq_bits_head(io_to_noc_0_flit_q_io_enq_bits_head),
    .io_enq_bits_tail(io_to_noc_0_flit_q_io_enq_bits_tail),
    .io_enq_bits_payload(io_to_noc_0_flit_q_io_enq_bits_payload),
    .io_enq_bits_egress_id(io_to_noc_0_flit_q_io_enq_bits_egress_id),
    .io_deq_ready(io_to_noc_0_flit_q_io_deq_ready),
    .io_deq_valid(io_to_noc_0_flit_q_io_deq_valid),
    .io_deq_bits_head(io_to_noc_0_flit_q_io_deq_bits_head),
    .io_deq_bits_tail(io_to_noc_0_flit_q_io_deq_bits_tail),
    .io_deq_bits_payload(io_to_noc_0_flit_q_io_deq_bits_payload),
    .io_deq_bits_egress_id(io_to_noc_0_flit_q_io_deq_bits_egress_id)
  );
  InputGen igen_1 ( // @[TestHarness.scala 171:22]
    .clock(igen_1_clock),
    .reset(igen_1_reset),
    .io_out_ready(igen_1_io_out_ready),
    .io_out_valid(igen_1_io_out_valid),
    .io_out_bits_head(igen_1_io_out_bits_head),
    .io_out_bits_tail(igen_1_io_out_bits_tail),
    .io_out_bits_payload(igen_1_io_out_bits_payload),
    .io_out_bits_egress_id(igen_1_io_out_bits_egress_id),
    .io_rob_ready(igen_1_io_rob_ready),
    .io_rob_idx(igen_1_io_rob_idx),
    .io_tsc(igen_1_io_tsc),
    .io_fire(igen_1_io_fire),
    .io_n_flits(igen_1_io_n_flits)
  );
  Queue_26 io_to_noc_1_flit_q ( // @[Decoupled.scala 375:21]
    .clock(io_to_noc_1_flit_q_clock),
    .reset(io_to_noc_1_flit_q_reset),
    .io_enq_ready(io_to_noc_1_flit_q_io_enq_ready),
    .io_enq_valid(io_to_noc_1_flit_q_io_enq_valid),
    .io_enq_bits_head(io_to_noc_1_flit_q_io_enq_bits_head),
    .io_enq_bits_tail(io_to_noc_1_flit_q_io_enq_bits_tail),
    .io_enq_bits_payload(io_to_noc_1_flit_q_io_enq_bits_payload),
    .io_enq_bits_egress_id(io_to_noc_1_flit_q_io_enq_bits_egress_id),
    .io_deq_ready(io_to_noc_1_flit_q_io_deq_ready),
    .io_deq_valid(io_to_noc_1_flit_q_io_deq_valid),
    .io_deq_bits_head(io_to_noc_1_flit_q_io_deq_bits_head),
    .io_deq_bits_tail(io_to_noc_1_flit_q_io_deq_bits_tail),
    .io_deq_bits_payload(io_to_noc_1_flit_q_io_deq_bits_payload),
    .io_deq_bits_egress_id(io_to_noc_1_flit_q_io_deq_bits_egress_id)
  );
  plusarg_reader #(.FORMAT("noctest_enable_print=%d"), .DEFAULT(0), .WIDTH(1)) plusarg_reader ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_out)
  );
  MaxPeriodFibonacciLFSR io_from_noc_0_flit_ready_prng ( // @[PRNG.scala 91:22]
    .clock(io_from_noc_0_flit_ready_prng_clock),
    .reset(io_from_noc_0_flit_ready_prng_reset),
    .io_out_0(io_from_noc_0_flit_ready_prng_io_out_0),
    .io_out_1(io_from_noc_0_flit_ready_prng_io_out_1),
    .io_out_2(io_from_noc_0_flit_ready_prng_io_out_2),
    .io_out_3(io_from_noc_0_flit_ready_prng_io_out_3),
    .io_out_4(io_from_noc_0_flit_ready_prng_io_out_4),
    .io_out_5(io_from_noc_0_flit_ready_prng_io_out_5),
    .io_out_6(io_from_noc_0_flit_ready_prng_io_out_6),
    .io_out_7(io_from_noc_0_flit_ready_prng_io_out_7),
    .io_out_8(io_from_noc_0_flit_ready_prng_io_out_8),
    .io_out_9(io_from_noc_0_flit_ready_prng_io_out_9),
    .io_out_10(io_from_noc_0_flit_ready_prng_io_out_10),
    .io_out_11(io_from_noc_0_flit_ready_prng_io_out_11),
    .io_out_12(io_from_noc_0_flit_ready_prng_io_out_12),
    .io_out_13(io_from_noc_0_flit_ready_prng_io_out_13),
    .io_out_14(io_from_noc_0_flit_ready_prng_io_out_14),
    .io_out_15(io_from_noc_0_flit_ready_prng_io_out_15),
    .io_out_16(io_from_noc_0_flit_ready_prng_io_out_16),
    .io_out_17(io_from_noc_0_flit_ready_prng_io_out_17),
    .io_out_18(io_from_noc_0_flit_ready_prng_io_out_18),
    .io_out_19(io_from_noc_0_flit_ready_prng_io_out_19)
  );
  MaxPeriodFibonacciLFSR io_from_noc_1_flit_ready_prng ( // @[PRNG.scala 91:22]
    .clock(io_from_noc_1_flit_ready_prng_clock),
    .reset(io_from_noc_1_flit_ready_prng_reset),
    .io_out_0(io_from_noc_1_flit_ready_prng_io_out_0),
    .io_out_1(io_from_noc_1_flit_ready_prng_io_out_1),
    .io_out_2(io_from_noc_1_flit_ready_prng_io_out_2),
    .io_out_3(io_from_noc_1_flit_ready_prng_io_out_3),
    .io_out_4(io_from_noc_1_flit_ready_prng_io_out_4),
    .io_out_5(io_from_noc_1_flit_ready_prng_io_out_5),
    .io_out_6(io_from_noc_1_flit_ready_prng_io_out_6),
    .io_out_7(io_from_noc_1_flit_ready_prng_io_out_7),
    .io_out_8(io_from_noc_1_flit_ready_prng_io_out_8),
    .io_out_9(io_from_noc_1_flit_ready_prng_io_out_9),
    .io_out_10(io_from_noc_1_flit_ready_prng_io_out_10),
    .io_out_11(io_from_noc_1_flit_ready_prng_io_out_11),
    .io_out_12(io_from_noc_1_flit_ready_prng_io_out_12),
    .io_out_13(io_from_noc_1_flit_ready_prng_io_out_13),
    .io_out_14(io_from_noc_1_flit_ready_prng_io_out_14),
    .io_out_15(io_from_noc_1_flit_ready_prng_io_out_15),
    .io_out_16(io_from_noc_1_flit_ready_prng_io_out_16),
    .io_out_17(io_from_noc_1_flit_ready_prng_io_out_17),
    .io_out_18(io_from_noc_1_flit_ready_prng_io_out_18),
    .io_out_19(io_from_noc_1_flit_ready_prng_io_out_19)
  );
  assign io_to_noc_1_flit_valid = io_to_noc_1_flit_q_io_deq_valid; // @[TestHarness.scala 177:12]
  assign io_to_noc_1_flit_bits_head = io_to_noc_1_flit_q_io_deq_bits_head; // @[TestHarness.scala 177:12]
  assign io_to_noc_1_flit_bits_tail = io_to_noc_1_flit_q_io_deq_bits_tail; // @[TestHarness.scala 177:12]
  assign io_to_noc_1_flit_bits_payload = io_to_noc_1_flit_q_io_deq_bits_payload; // @[TestHarness.scala 177:12]
  assign io_to_noc_1_flit_bits_egress_id = io_to_noc_1_flit_q_io_deq_bits_egress_id; // @[TestHarness.scala 177:12]
  assign io_to_noc_0_flit_valid = io_to_noc_0_flit_q_io_deq_valid; // @[TestHarness.scala 177:12]
  assign io_to_noc_0_flit_bits_head = io_to_noc_0_flit_q_io_deq_bits_head; // @[TestHarness.scala 177:12]
  assign io_to_noc_0_flit_bits_tail = io_to_noc_0_flit_q_io_deq_bits_tail; // @[TestHarness.scala 177:12]
  assign io_to_noc_0_flit_bits_payload = io_to_noc_0_flit_q_io_deq_bits_payload; // @[TestHarness.scala 177:12]
  assign io_to_noc_0_flit_bits_egress_id = io_to_noc_0_flit_q_io_deq_bits_egress_id; // @[TestHarness.scala 177:12]
  assign io_from_noc_1_flit_ready = 1'h1; // @[TestHarness.scala 193:30]
  assign io_from_noc_0_flit_ready = 1'h1; // @[TestHarness.scala 193:30]
  assign io_success = io_success_REG; // @[TestHarness.scala 164:14]
  assign igen_clock = clock;
  assign igen_reset = reset;
  assign igen_io_out_ready = io_to_noc_0_flit_q_io_enq_ready; // @[Decoupled.scala 379:17]
  assign igen_io_rob_ready = _igen_io_rob_ready_T_2 & txs < 32'hc350; // @[TestHarness.scala 175:19]
  assign igen_io_rob_idx = _T_5[0] ? 7'h0 : _sels_0_T_253; // @[Mux.scala 47:70]
  assign igen_io_tsc = tsc; // @[TestHarness.scala 176:17]
  assign io_to_noc_0_flit_q_clock = clock;
  assign io_to_noc_0_flit_q_reset = reset;
  assign io_to_noc_0_flit_q_io_enq_valid = igen_io_out_valid; // @[Decoupled.scala 377:22]
  assign io_to_noc_0_flit_q_io_enq_bits_head = igen_io_out_bits_head; // @[Decoupled.scala 378:21]
  assign io_to_noc_0_flit_q_io_enq_bits_tail = igen_io_out_bits_tail; // @[Decoupled.scala 378:21]
  assign io_to_noc_0_flit_q_io_enq_bits_payload = igen_io_out_bits_payload; // @[Decoupled.scala 378:21]
  assign io_to_noc_0_flit_q_io_enq_bits_egress_id = igen_io_out_bits_egress_id; // @[Decoupled.scala 378:21]
  assign io_to_noc_0_flit_q_io_deq_ready = io_to_noc_0_flit_ready; // @[TestHarness.scala 177:12]
  assign igen_1_clock = clock;
  assign igen_1_reset = reset;
  assign igen_1_io_out_ready = io_to_noc_1_flit_q_io_enq_ready; // @[Decoupled.scala 379:17]
  assign igen_1_io_rob_ready = _igen_io_rob_ready_T_7 & txs < 32'hc350; // @[TestHarness.scala 175:19]
  assign igen_1_io_rob_idx = _T_8[0] ? 7'h0 : _sels_1_T_253; // @[Mux.scala 47:70]
  assign igen_1_io_tsc = tsc; // @[TestHarness.scala 176:17]
  assign io_to_noc_1_flit_q_clock = clock;
  assign io_to_noc_1_flit_q_reset = reset;
  assign io_to_noc_1_flit_q_io_enq_valid = igen_1_io_out_valid; // @[Decoupled.scala 377:22]
  assign io_to_noc_1_flit_q_io_enq_bits_head = igen_1_io_out_bits_head; // @[Decoupled.scala 378:21]
  assign io_to_noc_1_flit_q_io_enq_bits_tail = igen_1_io_out_bits_tail; // @[Decoupled.scala 378:21]
  assign io_to_noc_1_flit_q_io_enq_bits_payload = igen_1_io_out_bits_payload; // @[Decoupled.scala 378:21]
  assign io_to_noc_1_flit_q_io_enq_bits_egress_id = igen_1_io_out_bits_egress_id; // @[Decoupled.scala 378:21]
  assign io_to_noc_1_flit_q_io_deq_ready = io_to_noc_1_flit_ready; // @[TestHarness.scala 177:12]
  assign io_from_noc_0_flit_ready_prng_clock = clock;
  assign io_from_noc_0_flit_ready_prng_reset = reset;
  assign io_from_noc_1_flit_ready_prng_clock = clock;
  assign io_from_noc_1_flit_ready_prng_reset = reset;
  always @(posedge clock) begin
    if (reset) begin // @[TestHarness.scala 136:20]
      txs <= 32'h0; // @[TestHarness.scala 136:20]
    end else begin
      txs <= _txs_T_3; // @[TestHarness.scala 225:7]
    end
    if (reset) begin // @[TestHarness.scala 137:22]
      flits <= 32'h0; // @[TestHarness.scala 137:22]
    end else begin
      flits <= _flits_T_4; // @[TestHarness.scala 224:9]
    end
    if (reset) begin // @[TestHarness.scala 141:20]
      tsc <= 32'h0; // @[TestHarness.scala 141:20]
    end else begin
      tsc <= _tsc_T_1; // @[TestHarness.scala 142:7]
    end
    if (reset) begin // @[TestHarness.scala 144:29]
      idle_counter <= 11'h0; // @[TestHarness.scala 144:29]
    end else if (idle) begin // @[TestHarness.scala 146:15]
      idle_counter <= _idle_counter_T_1; // @[TestHarness.scala 146:30]
    end else begin
      idle_counter <= 11'h0; // @[TestHarness.scala 147:31]
    end
    rob_valids <= _GEN_7952[127:0]; // @[TestHarness.scala 156:{27,27} 222:14]
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h0 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_0_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_0_tsc <= _GEN_1025;
      end
    end else begin
      rob_payload_0_tsc <= _GEN_1025;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h0 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_0_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_0_rob_idx <= _GEN_1153;
      end
    end else begin
      rob_payload_0_rob_idx <= _GEN_1153;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h0 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_0_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_0_flits_fired <= _GEN_5764;
      end
    end else begin
      rob_payload_0_flits_fired <= _GEN_5764;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_1_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_1_tsc <= _GEN_1026;
      end
    end else begin
      rob_payload_1_tsc <= _GEN_1026;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_1_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_1_rob_idx <= _GEN_1154;
      end
    end else begin
      rob_payload_1_rob_idx <= _GEN_1154;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h1 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_1_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_1_flits_fired <= _GEN_5765;
      end
    end else begin
      rob_payload_1_flits_fired <= _GEN_5765;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_2_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_2_tsc <= _GEN_1027;
      end
    end else begin
      rob_payload_2_tsc <= _GEN_1027;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_2_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_2_rob_idx <= _GEN_1155;
      end
    end else begin
      rob_payload_2_rob_idx <= _GEN_1155;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h2 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_2_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_2_flits_fired <= _GEN_5766;
      end
    end else begin
      rob_payload_2_flits_fired <= _GEN_5766;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_3_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_3_tsc <= _GEN_1028;
      end
    end else begin
      rob_payload_3_tsc <= _GEN_1028;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_3_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_3_rob_idx <= _GEN_1156;
      end
    end else begin
      rob_payload_3_rob_idx <= _GEN_1156;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h3 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_3_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_3_flits_fired <= _GEN_5767;
      end
    end else begin
      rob_payload_3_flits_fired <= _GEN_5767;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_4_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_4_tsc <= _GEN_1029;
      end
    end else begin
      rob_payload_4_tsc <= _GEN_1029;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_4_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_4_rob_idx <= _GEN_1157;
      end
    end else begin
      rob_payload_4_rob_idx <= _GEN_1157;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h4 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_4_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_4_flits_fired <= _GEN_5768;
      end
    end else begin
      rob_payload_4_flits_fired <= _GEN_5768;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_5_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_5_tsc <= _GEN_1030;
      end
    end else begin
      rob_payload_5_tsc <= _GEN_1030;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_5_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_5_rob_idx <= _GEN_1158;
      end
    end else begin
      rob_payload_5_rob_idx <= _GEN_1158;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h5 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_5_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_5_flits_fired <= _GEN_5769;
      end
    end else begin
      rob_payload_5_flits_fired <= _GEN_5769;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_6_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_6_tsc <= _GEN_1031;
      end
    end else begin
      rob_payload_6_tsc <= _GEN_1031;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_6_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_6_rob_idx <= _GEN_1159;
      end
    end else begin
      rob_payload_6_rob_idx <= _GEN_1159;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h6 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_6_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_6_flits_fired <= _GEN_5770;
      end
    end else begin
      rob_payload_6_flits_fired <= _GEN_5770;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_7_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_7_tsc <= _GEN_1032;
      end
    end else begin
      rob_payload_7_tsc <= _GEN_1032;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_7_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_7_rob_idx <= _GEN_1160;
      end
    end else begin
      rob_payload_7_rob_idx <= _GEN_1160;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h7 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_7_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_7_flits_fired <= _GEN_5771;
      end
    end else begin
      rob_payload_7_flits_fired <= _GEN_5771;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h8 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_8_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_8_tsc <= _GEN_1033;
      end
    end else begin
      rob_payload_8_tsc <= _GEN_1033;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h8 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_8_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_8_rob_idx <= _GEN_1161;
      end
    end else begin
      rob_payload_8_rob_idx <= _GEN_1161;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h8 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_8_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_8_flits_fired <= _GEN_5772;
      end
    end else begin
      rob_payload_8_flits_fired <= _GEN_5772;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h9 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_9_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_9_tsc <= _GEN_1034;
      end
    end else begin
      rob_payload_9_tsc <= _GEN_1034;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h9 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_9_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_9_rob_idx <= _GEN_1162;
      end
    end else begin
      rob_payload_9_rob_idx <= _GEN_1162;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h9 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_9_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_9_flits_fired <= _GEN_5773;
      end
    end else begin
      rob_payload_9_flits_fired <= _GEN_5773;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'ha == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_10_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_10_tsc <= _GEN_1035;
      end
    end else begin
      rob_payload_10_tsc <= _GEN_1035;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'ha == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_10_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_10_rob_idx <= _GEN_1163;
      end
    end else begin
      rob_payload_10_rob_idx <= _GEN_1163;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'ha == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_10_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_10_flits_fired <= _GEN_5774;
      end
    end else begin
      rob_payload_10_flits_fired <= _GEN_5774;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hb == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_11_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_11_tsc <= _GEN_1036;
      end
    end else begin
      rob_payload_11_tsc <= _GEN_1036;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hb == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_11_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_11_rob_idx <= _GEN_1164;
      end
    end else begin
      rob_payload_11_rob_idx <= _GEN_1164;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'hb == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_11_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_11_flits_fired <= _GEN_5775;
      end
    end else begin
      rob_payload_11_flits_fired <= _GEN_5775;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hc == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_12_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_12_tsc <= _GEN_1037;
      end
    end else begin
      rob_payload_12_tsc <= _GEN_1037;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hc == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_12_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_12_rob_idx <= _GEN_1165;
      end
    end else begin
      rob_payload_12_rob_idx <= _GEN_1165;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'hc == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_12_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_12_flits_fired <= _GEN_5776;
      end
    end else begin
      rob_payload_12_flits_fired <= _GEN_5776;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hd == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_13_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_13_tsc <= _GEN_1038;
      end
    end else begin
      rob_payload_13_tsc <= _GEN_1038;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hd == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_13_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_13_rob_idx <= _GEN_1166;
      end
    end else begin
      rob_payload_13_rob_idx <= _GEN_1166;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'hd == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_13_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_13_flits_fired <= _GEN_5777;
      end
    end else begin
      rob_payload_13_flits_fired <= _GEN_5777;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'he == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_14_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_14_tsc <= _GEN_1039;
      end
    end else begin
      rob_payload_14_tsc <= _GEN_1039;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'he == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_14_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_14_rob_idx <= _GEN_1167;
      end
    end else begin
      rob_payload_14_rob_idx <= _GEN_1167;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'he == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_14_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_14_flits_fired <= _GEN_5778;
      end
    end else begin
      rob_payload_14_flits_fired <= _GEN_5778;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hf == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_15_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_15_tsc <= _GEN_1040;
      end
    end else begin
      rob_payload_15_tsc <= _GEN_1040;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hf == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_15_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_15_rob_idx <= _GEN_1168;
      end
    end else begin
      rob_payload_15_rob_idx <= _GEN_1168;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'hf == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_15_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_15_flits_fired <= _GEN_5779;
      end
    end else begin
      rob_payload_15_flits_fired <= _GEN_5779;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h10 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_16_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_16_tsc <= _GEN_1041;
      end
    end else begin
      rob_payload_16_tsc <= _GEN_1041;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h10 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_16_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_16_rob_idx <= _GEN_1169;
      end
    end else begin
      rob_payload_16_rob_idx <= _GEN_1169;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h10 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_16_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_16_flits_fired <= _GEN_5780;
      end
    end else begin
      rob_payload_16_flits_fired <= _GEN_5780;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h11 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_17_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_17_tsc <= _GEN_1042;
      end
    end else begin
      rob_payload_17_tsc <= _GEN_1042;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h11 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_17_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_17_rob_idx <= _GEN_1170;
      end
    end else begin
      rob_payload_17_rob_idx <= _GEN_1170;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h11 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_17_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_17_flits_fired <= _GEN_5781;
      end
    end else begin
      rob_payload_17_flits_fired <= _GEN_5781;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h12 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_18_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_18_tsc <= _GEN_1043;
      end
    end else begin
      rob_payload_18_tsc <= _GEN_1043;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h12 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_18_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_18_rob_idx <= _GEN_1171;
      end
    end else begin
      rob_payload_18_rob_idx <= _GEN_1171;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h12 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_18_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_18_flits_fired <= _GEN_5782;
      end
    end else begin
      rob_payload_18_flits_fired <= _GEN_5782;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h13 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_19_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_19_tsc <= _GEN_1044;
      end
    end else begin
      rob_payload_19_tsc <= _GEN_1044;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h13 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_19_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_19_rob_idx <= _GEN_1172;
      end
    end else begin
      rob_payload_19_rob_idx <= _GEN_1172;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h13 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_19_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_19_flits_fired <= _GEN_5783;
      end
    end else begin
      rob_payload_19_flits_fired <= _GEN_5783;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h14 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_20_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_20_tsc <= _GEN_1045;
      end
    end else begin
      rob_payload_20_tsc <= _GEN_1045;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h14 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_20_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_20_rob_idx <= _GEN_1173;
      end
    end else begin
      rob_payload_20_rob_idx <= _GEN_1173;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h14 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_20_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_20_flits_fired <= _GEN_5784;
      end
    end else begin
      rob_payload_20_flits_fired <= _GEN_5784;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h15 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_21_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_21_tsc <= _GEN_1046;
      end
    end else begin
      rob_payload_21_tsc <= _GEN_1046;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h15 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_21_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_21_rob_idx <= _GEN_1174;
      end
    end else begin
      rob_payload_21_rob_idx <= _GEN_1174;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h15 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_21_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_21_flits_fired <= _GEN_5785;
      end
    end else begin
      rob_payload_21_flits_fired <= _GEN_5785;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h16 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_22_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_22_tsc <= _GEN_1047;
      end
    end else begin
      rob_payload_22_tsc <= _GEN_1047;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h16 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_22_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_22_rob_idx <= _GEN_1175;
      end
    end else begin
      rob_payload_22_rob_idx <= _GEN_1175;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h16 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_22_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_22_flits_fired <= _GEN_5786;
      end
    end else begin
      rob_payload_22_flits_fired <= _GEN_5786;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h17 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_23_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_23_tsc <= _GEN_1048;
      end
    end else begin
      rob_payload_23_tsc <= _GEN_1048;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h17 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_23_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_23_rob_idx <= _GEN_1176;
      end
    end else begin
      rob_payload_23_rob_idx <= _GEN_1176;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h17 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_23_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_23_flits_fired <= _GEN_5787;
      end
    end else begin
      rob_payload_23_flits_fired <= _GEN_5787;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h18 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_24_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_24_tsc <= _GEN_1049;
      end
    end else begin
      rob_payload_24_tsc <= _GEN_1049;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h18 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_24_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_24_rob_idx <= _GEN_1177;
      end
    end else begin
      rob_payload_24_rob_idx <= _GEN_1177;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h18 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_24_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_24_flits_fired <= _GEN_5788;
      end
    end else begin
      rob_payload_24_flits_fired <= _GEN_5788;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h19 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_25_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_25_tsc <= _GEN_1050;
      end
    end else begin
      rob_payload_25_tsc <= _GEN_1050;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h19 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_25_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_25_rob_idx <= _GEN_1178;
      end
    end else begin
      rob_payload_25_rob_idx <= _GEN_1178;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h19 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_25_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_25_flits_fired <= _GEN_5789;
      end
    end else begin
      rob_payload_25_flits_fired <= _GEN_5789;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1a == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_26_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_26_tsc <= _GEN_1051;
      end
    end else begin
      rob_payload_26_tsc <= _GEN_1051;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1a == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_26_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_26_rob_idx <= _GEN_1179;
      end
    end else begin
      rob_payload_26_rob_idx <= _GEN_1179;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h1a == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_26_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_26_flits_fired <= _GEN_5790;
      end
    end else begin
      rob_payload_26_flits_fired <= _GEN_5790;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1b == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_27_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_27_tsc <= _GEN_1052;
      end
    end else begin
      rob_payload_27_tsc <= _GEN_1052;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1b == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_27_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_27_rob_idx <= _GEN_1180;
      end
    end else begin
      rob_payload_27_rob_idx <= _GEN_1180;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h1b == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_27_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_27_flits_fired <= _GEN_5791;
      end
    end else begin
      rob_payload_27_flits_fired <= _GEN_5791;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1c == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_28_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_28_tsc <= _GEN_1053;
      end
    end else begin
      rob_payload_28_tsc <= _GEN_1053;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1c == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_28_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_28_rob_idx <= _GEN_1181;
      end
    end else begin
      rob_payload_28_rob_idx <= _GEN_1181;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h1c == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_28_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_28_flits_fired <= _GEN_5792;
      end
    end else begin
      rob_payload_28_flits_fired <= _GEN_5792;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1d == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_29_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_29_tsc <= _GEN_1054;
      end
    end else begin
      rob_payload_29_tsc <= _GEN_1054;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1d == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_29_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_29_rob_idx <= _GEN_1182;
      end
    end else begin
      rob_payload_29_rob_idx <= _GEN_1182;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h1d == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_29_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_29_flits_fired <= _GEN_5793;
      end
    end else begin
      rob_payload_29_flits_fired <= _GEN_5793;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1e == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_30_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_30_tsc <= _GEN_1055;
      end
    end else begin
      rob_payload_30_tsc <= _GEN_1055;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1e == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_30_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_30_rob_idx <= _GEN_1183;
      end
    end else begin
      rob_payload_30_rob_idx <= _GEN_1183;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h1e == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_30_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_30_flits_fired <= _GEN_5794;
      end
    end else begin
      rob_payload_30_flits_fired <= _GEN_5794;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1f == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_31_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_31_tsc <= _GEN_1056;
      end
    end else begin
      rob_payload_31_tsc <= _GEN_1056;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1f == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_31_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_31_rob_idx <= _GEN_1184;
      end
    end else begin
      rob_payload_31_rob_idx <= _GEN_1184;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h1f == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_31_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_31_flits_fired <= _GEN_5795;
      end
    end else begin
      rob_payload_31_flits_fired <= _GEN_5795;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h20 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_32_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_32_tsc <= _GEN_1057;
      end
    end else begin
      rob_payload_32_tsc <= _GEN_1057;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h20 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_32_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_32_rob_idx <= _GEN_1185;
      end
    end else begin
      rob_payload_32_rob_idx <= _GEN_1185;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h20 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_32_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_32_flits_fired <= _GEN_5796;
      end
    end else begin
      rob_payload_32_flits_fired <= _GEN_5796;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h21 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_33_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_33_tsc <= _GEN_1058;
      end
    end else begin
      rob_payload_33_tsc <= _GEN_1058;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h21 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_33_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_33_rob_idx <= _GEN_1186;
      end
    end else begin
      rob_payload_33_rob_idx <= _GEN_1186;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h21 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_33_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_33_flits_fired <= _GEN_5797;
      end
    end else begin
      rob_payload_33_flits_fired <= _GEN_5797;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h22 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_34_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_34_tsc <= _GEN_1059;
      end
    end else begin
      rob_payload_34_tsc <= _GEN_1059;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h22 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_34_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_34_rob_idx <= _GEN_1187;
      end
    end else begin
      rob_payload_34_rob_idx <= _GEN_1187;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h22 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_34_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_34_flits_fired <= _GEN_5798;
      end
    end else begin
      rob_payload_34_flits_fired <= _GEN_5798;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h23 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_35_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_35_tsc <= _GEN_1060;
      end
    end else begin
      rob_payload_35_tsc <= _GEN_1060;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h23 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_35_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_35_rob_idx <= _GEN_1188;
      end
    end else begin
      rob_payload_35_rob_idx <= _GEN_1188;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h23 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_35_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_35_flits_fired <= _GEN_5799;
      end
    end else begin
      rob_payload_35_flits_fired <= _GEN_5799;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h24 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_36_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_36_tsc <= _GEN_1061;
      end
    end else begin
      rob_payload_36_tsc <= _GEN_1061;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h24 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_36_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_36_rob_idx <= _GEN_1189;
      end
    end else begin
      rob_payload_36_rob_idx <= _GEN_1189;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h24 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_36_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_36_flits_fired <= _GEN_5800;
      end
    end else begin
      rob_payload_36_flits_fired <= _GEN_5800;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h25 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_37_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_37_tsc <= _GEN_1062;
      end
    end else begin
      rob_payload_37_tsc <= _GEN_1062;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h25 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_37_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_37_rob_idx <= _GEN_1190;
      end
    end else begin
      rob_payload_37_rob_idx <= _GEN_1190;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h25 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_37_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_37_flits_fired <= _GEN_5801;
      end
    end else begin
      rob_payload_37_flits_fired <= _GEN_5801;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h26 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_38_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_38_tsc <= _GEN_1063;
      end
    end else begin
      rob_payload_38_tsc <= _GEN_1063;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h26 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_38_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_38_rob_idx <= _GEN_1191;
      end
    end else begin
      rob_payload_38_rob_idx <= _GEN_1191;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h26 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_38_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_38_flits_fired <= _GEN_5802;
      end
    end else begin
      rob_payload_38_flits_fired <= _GEN_5802;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h27 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_39_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_39_tsc <= _GEN_1064;
      end
    end else begin
      rob_payload_39_tsc <= _GEN_1064;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h27 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_39_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_39_rob_idx <= _GEN_1192;
      end
    end else begin
      rob_payload_39_rob_idx <= _GEN_1192;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h27 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_39_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_39_flits_fired <= _GEN_5803;
      end
    end else begin
      rob_payload_39_flits_fired <= _GEN_5803;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h28 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_40_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_40_tsc <= _GEN_1065;
      end
    end else begin
      rob_payload_40_tsc <= _GEN_1065;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h28 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_40_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_40_rob_idx <= _GEN_1193;
      end
    end else begin
      rob_payload_40_rob_idx <= _GEN_1193;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h28 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_40_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_40_flits_fired <= _GEN_5804;
      end
    end else begin
      rob_payload_40_flits_fired <= _GEN_5804;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h29 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_41_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_41_tsc <= _GEN_1066;
      end
    end else begin
      rob_payload_41_tsc <= _GEN_1066;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h29 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_41_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_41_rob_idx <= _GEN_1194;
      end
    end else begin
      rob_payload_41_rob_idx <= _GEN_1194;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h29 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_41_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_41_flits_fired <= _GEN_5805;
      end
    end else begin
      rob_payload_41_flits_fired <= _GEN_5805;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2a == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_42_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_42_tsc <= _GEN_1067;
      end
    end else begin
      rob_payload_42_tsc <= _GEN_1067;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2a == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_42_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_42_rob_idx <= _GEN_1195;
      end
    end else begin
      rob_payload_42_rob_idx <= _GEN_1195;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h2a == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_42_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_42_flits_fired <= _GEN_5806;
      end
    end else begin
      rob_payload_42_flits_fired <= _GEN_5806;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2b == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_43_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_43_tsc <= _GEN_1068;
      end
    end else begin
      rob_payload_43_tsc <= _GEN_1068;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2b == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_43_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_43_rob_idx <= _GEN_1196;
      end
    end else begin
      rob_payload_43_rob_idx <= _GEN_1196;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h2b == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_43_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_43_flits_fired <= _GEN_5807;
      end
    end else begin
      rob_payload_43_flits_fired <= _GEN_5807;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2c == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_44_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_44_tsc <= _GEN_1069;
      end
    end else begin
      rob_payload_44_tsc <= _GEN_1069;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2c == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_44_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_44_rob_idx <= _GEN_1197;
      end
    end else begin
      rob_payload_44_rob_idx <= _GEN_1197;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h2c == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_44_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_44_flits_fired <= _GEN_5808;
      end
    end else begin
      rob_payload_44_flits_fired <= _GEN_5808;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2d == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_45_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_45_tsc <= _GEN_1070;
      end
    end else begin
      rob_payload_45_tsc <= _GEN_1070;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2d == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_45_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_45_rob_idx <= _GEN_1198;
      end
    end else begin
      rob_payload_45_rob_idx <= _GEN_1198;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h2d == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_45_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_45_flits_fired <= _GEN_5809;
      end
    end else begin
      rob_payload_45_flits_fired <= _GEN_5809;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2e == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_46_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_46_tsc <= _GEN_1071;
      end
    end else begin
      rob_payload_46_tsc <= _GEN_1071;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2e == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_46_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_46_rob_idx <= _GEN_1199;
      end
    end else begin
      rob_payload_46_rob_idx <= _GEN_1199;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h2e == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_46_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_46_flits_fired <= _GEN_5810;
      end
    end else begin
      rob_payload_46_flits_fired <= _GEN_5810;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2f == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_47_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_47_tsc <= _GEN_1072;
      end
    end else begin
      rob_payload_47_tsc <= _GEN_1072;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2f == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_47_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_47_rob_idx <= _GEN_1200;
      end
    end else begin
      rob_payload_47_rob_idx <= _GEN_1200;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h2f == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_47_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_47_flits_fired <= _GEN_5811;
      end
    end else begin
      rob_payload_47_flits_fired <= _GEN_5811;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h30 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_48_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_48_tsc <= _GEN_1073;
      end
    end else begin
      rob_payload_48_tsc <= _GEN_1073;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h30 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_48_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_48_rob_idx <= _GEN_1201;
      end
    end else begin
      rob_payload_48_rob_idx <= _GEN_1201;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h30 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_48_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_48_flits_fired <= _GEN_5812;
      end
    end else begin
      rob_payload_48_flits_fired <= _GEN_5812;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h31 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_49_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_49_tsc <= _GEN_1074;
      end
    end else begin
      rob_payload_49_tsc <= _GEN_1074;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h31 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_49_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_49_rob_idx <= _GEN_1202;
      end
    end else begin
      rob_payload_49_rob_idx <= _GEN_1202;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h31 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_49_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_49_flits_fired <= _GEN_5813;
      end
    end else begin
      rob_payload_49_flits_fired <= _GEN_5813;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h32 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_50_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_50_tsc <= _GEN_1075;
      end
    end else begin
      rob_payload_50_tsc <= _GEN_1075;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h32 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_50_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_50_rob_idx <= _GEN_1203;
      end
    end else begin
      rob_payload_50_rob_idx <= _GEN_1203;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h32 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_50_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_50_flits_fired <= _GEN_5814;
      end
    end else begin
      rob_payload_50_flits_fired <= _GEN_5814;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h33 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_51_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_51_tsc <= _GEN_1076;
      end
    end else begin
      rob_payload_51_tsc <= _GEN_1076;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h33 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_51_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_51_rob_idx <= _GEN_1204;
      end
    end else begin
      rob_payload_51_rob_idx <= _GEN_1204;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h33 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_51_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_51_flits_fired <= _GEN_5815;
      end
    end else begin
      rob_payload_51_flits_fired <= _GEN_5815;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h34 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_52_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_52_tsc <= _GEN_1077;
      end
    end else begin
      rob_payload_52_tsc <= _GEN_1077;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h34 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_52_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_52_rob_idx <= _GEN_1205;
      end
    end else begin
      rob_payload_52_rob_idx <= _GEN_1205;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h34 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_52_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_52_flits_fired <= _GEN_5816;
      end
    end else begin
      rob_payload_52_flits_fired <= _GEN_5816;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h35 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_53_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_53_tsc <= _GEN_1078;
      end
    end else begin
      rob_payload_53_tsc <= _GEN_1078;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h35 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_53_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_53_rob_idx <= _GEN_1206;
      end
    end else begin
      rob_payload_53_rob_idx <= _GEN_1206;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h35 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_53_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_53_flits_fired <= _GEN_5817;
      end
    end else begin
      rob_payload_53_flits_fired <= _GEN_5817;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h36 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_54_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_54_tsc <= _GEN_1079;
      end
    end else begin
      rob_payload_54_tsc <= _GEN_1079;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h36 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_54_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_54_rob_idx <= _GEN_1207;
      end
    end else begin
      rob_payload_54_rob_idx <= _GEN_1207;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h36 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_54_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_54_flits_fired <= _GEN_5818;
      end
    end else begin
      rob_payload_54_flits_fired <= _GEN_5818;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h37 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_55_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_55_tsc <= _GEN_1080;
      end
    end else begin
      rob_payload_55_tsc <= _GEN_1080;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h37 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_55_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_55_rob_idx <= _GEN_1208;
      end
    end else begin
      rob_payload_55_rob_idx <= _GEN_1208;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h37 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_55_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_55_flits_fired <= _GEN_5819;
      end
    end else begin
      rob_payload_55_flits_fired <= _GEN_5819;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h38 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_56_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_56_tsc <= _GEN_1081;
      end
    end else begin
      rob_payload_56_tsc <= _GEN_1081;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h38 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_56_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_56_rob_idx <= _GEN_1209;
      end
    end else begin
      rob_payload_56_rob_idx <= _GEN_1209;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h38 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_56_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_56_flits_fired <= _GEN_5820;
      end
    end else begin
      rob_payload_56_flits_fired <= _GEN_5820;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h39 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_57_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_57_tsc <= _GEN_1082;
      end
    end else begin
      rob_payload_57_tsc <= _GEN_1082;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h39 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_57_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_57_rob_idx <= _GEN_1210;
      end
    end else begin
      rob_payload_57_rob_idx <= _GEN_1210;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h39 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_57_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_57_flits_fired <= _GEN_5821;
      end
    end else begin
      rob_payload_57_flits_fired <= _GEN_5821;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3a == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_58_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_58_tsc <= _GEN_1083;
      end
    end else begin
      rob_payload_58_tsc <= _GEN_1083;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3a == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_58_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_58_rob_idx <= _GEN_1211;
      end
    end else begin
      rob_payload_58_rob_idx <= _GEN_1211;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h3a == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_58_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_58_flits_fired <= _GEN_5822;
      end
    end else begin
      rob_payload_58_flits_fired <= _GEN_5822;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3b == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_59_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_59_tsc <= _GEN_1084;
      end
    end else begin
      rob_payload_59_tsc <= _GEN_1084;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3b == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_59_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_59_rob_idx <= _GEN_1212;
      end
    end else begin
      rob_payload_59_rob_idx <= _GEN_1212;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h3b == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_59_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_59_flits_fired <= _GEN_5823;
      end
    end else begin
      rob_payload_59_flits_fired <= _GEN_5823;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3c == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_60_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_60_tsc <= _GEN_1085;
      end
    end else begin
      rob_payload_60_tsc <= _GEN_1085;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3c == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_60_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_60_rob_idx <= _GEN_1213;
      end
    end else begin
      rob_payload_60_rob_idx <= _GEN_1213;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h3c == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_60_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_60_flits_fired <= _GEN_5824;
      end
    end else begin
      rob_payload_60_flits_fired <= _GEN_5824;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3d == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_61_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_61_tsc <= _GEN_1086;
      end
    end else begin
      rob_payload_61_tsc <= _GEN_1086;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3d == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_61_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_61_rob_idx <= _GEN_1214;
      end
    end else begin
      rob_payload_61_rob_idx <= _GEN_1214;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h3d == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_61_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_61_flits_fired <= _GEN_5825;
      end
    end else begin
      rob_payload_61_flits_fired <= _GEN_5825;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3e == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_62_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_62_tsc <= _GEN_1087;
      end
    end else begin
      rob_payload_62_tsc <= _GEN_1087;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3e == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_62_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_62_rob_idx <= _GEN_1215;
      end
    end else begin
      rob_payload_62_rob_idx <= _GEN_1215;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h3e == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_62_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_62_flits_fired <= _GEN_5826;
      end
    end else begin
      rob_payload_62_flits_fired <= _GEN_5826;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3f == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_63_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_63_tsc <= _GEN_1088;
      end
    end else begin
      rob_payload_63_tsc <= _GEN_1088;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3f == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_63_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_63_rob_idx <= _GEN_1216;
      end
    end else begin
      rob_payload_63_rob_idx <= _GEN_1216;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h3f == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_63_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_63_flits_fired <= _GEN_5827;
      end
    end else begin
      rob_payload_63_flits_fired <= _GEN_5827;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h40 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_64_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_64_tsc <= _GEN_1089;
      end
    end else begin
      rob_payload_64_tsc <= _GEN_1089;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h40 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_64_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_64_rob_idx <= _GEN_1217;
      end
    end else begin
      rob_payload_64_rob_idx <= _GEN_1217;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h40 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_64_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_64_flits_fired <= _GEN_5828;
      end
    end else begin
      rob_payload_64_flits_fired <= _GEN_5828;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h41 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_65_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_65_tsc <= _GEN_1090;
      end
    end else begin
      rob_payload_65_tsc <= _GEN_1090;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h41 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_65_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_65_rob_idx <= _GEN_1218;
      end
    end else begin
      rob_payload_65_rob_idx <= _GEN_1218;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h41 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_65_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_65_flits_fired <= _GEN_5829;
      end
    end else begin
      rob_payload_65_flits_fired <= _GEN_5829;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h42 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_66_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_66_tsc <= _GEN_1091;
      end
    end else begin
      rob_payload_66_tsc <= _GEN_1091;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h42 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_66_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_66_rob_idx <= _GEN_1219;
      end
    end else begin
      rob_payload_66_rob_idx <= _GEN_1219;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h42 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_66_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_66_flits_fired <= _GEN_5830;
      end
    end else begin
      rob_payload_66_flits_fired <= _GEN_5830;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h43 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_67_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_67_tsc <= _GEN_1092;
      end
    end else begin
      rob_payload_67_tsc <= _GEN_1092;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h43 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_67_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_67_rob_idx <= _GEN_1220;
      end
    end else begin
      rob_payload_67_rob_idx <= _GEN_1220;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h43 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_67_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_67_flits_fired <= _GEN_5831;
      end
    end else begin
      rob_payload_67_flits_fired <= _GEN_5831;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h44 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_68_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_68_tsc <= _GEN_1093;
      end
    end else begin
      rob_payload_68_tsc <= _GEN_1093;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h44 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_68_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_68_rob_idx <= _GEN_1221;
      end
    end else begin
      rob_payload_68_rob_idx <= _GEN_1221;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h44 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_68_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_68_flits_fired <= _GEN_5832;
      end
    end else begin
      rob_payload_68_flits_fired <= _GEN_5832;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h45 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_69_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_69_tsc <= _GEN_1094;
      end
    end else begin
      rob_payload_69_tsc <= _GEN_1094;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h45 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_69_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_69_rob_idx <= _GEN_1222;
      end
    end else begin
      rob_payload_69_rob_idx <= _GEN_1222;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h45 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_69_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_69_flits_fired <= _GEN_5833;
      end
    end else begin
      rob_payload_69_flits_fired <= _GEN_5833;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h46 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_70_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_70_tsc <= _GEN_1095;
      end
    end else begin
      rob_payload_70_tsc <= _GEN_1095;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h46 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_70_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_70_rob_idx <= _GEN_1223;
      end
    end else begin
      rob_payload_70_rob_idx <= _GEN_1223;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h46 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_70_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_70_flits_fired <= _GEN_5834;
      end
    end else begin
      rob_payload_70_flits_fired <= _GEN_5834;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h47 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_71_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_71_tsc <= _GEN_1096;
      end
    end else begin
      rob_payload_71_tsc <= _GEN_1096;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h47 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_71_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_71_rob_idx <= _GEN_1224;
      end
    end else begin
      rob_payload_71_rob_idx <= _GEN_1224;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h47 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_71_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_71_flits_fired <= _GEN_5835;
      end
    end else begin
      rob_payload_71_flits_fired <= _GEN_5835;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h48 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_72_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_72_tsc <= _GEN_1097;
      end
    end else begin
      rob_payload_72_tsc <= _GEN_1097;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h48 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_72_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_72_rob_idx <= _GEN_1225;
      end
    end else begin
      rob_payload_72_rob_idx <= _GEN_1225;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h48 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_72_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_72_flits_fired <= _GEN_5836;
      end
    end else begin
      rob_payload_72_flits_fired <= _GEN_5836;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h49 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_73_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_73_tsc <= _GEN_1098;
      end
    end else begin
      rob_payload_73_tsc <= _GEN_1098;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h49 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_73_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_73_rob_idx <= _GEN_1226;
      end
    end else begin
      rob_payload_73_rob_idx <= _GEN_1226;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h49 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_73_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_73_flits_fired <= _GEN_5837;
      end
    end else begin
      rob_payload_73_flits_fired <= _GEN_5837;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4a == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_74_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_74_tsc <= _GEN_1099;
      end
    end else begin
      rob_payload_74_tsc <= _GEN_1099;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4a == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_74_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_74_rob_idx <= _GEN_1227;
      end
    end else begin
      rob_payload_74_rob_idx <= _GEN_1227;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h4a == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_74_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_74_flits_fired <= _GEN_5838;
      end
    end else begin
      rob_payload_74_flits_fired <= _GEN_5838;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4b == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_75_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_75_tsc <= _GEN_1100;
      end
    end else begin
      rob_payload_75_tsc <= _GEN_1100;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4b == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_75_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_75_rob_idx <= _GEN_1228;
      end
    end else begin
      rob_payload_75_rob_idx <= _GEN_1228;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h4b == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_75_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_75_flits_fired <= _GEN_5839;
      end
    end else begin
      rob_payload_75_flits_fired <= _GEN_5839;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4c == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_76_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_76_tsc <= _GEN_1101;
      end
    end else begin
      rob_payload_76_tsc <= _GEN_1101;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4c == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_76_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_76_rob_idx <= _GEN_1229;
      end
    end else begin
      rob_payload_76_rob_idx <= _GEN_1229;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h4c == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_76_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_76_flits_fired <= _GEN_5840;
      end
    end else begin
      rob_payload_76_flits_fired <= _GEN_5840;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4d == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_77_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_77_tsc <= _GEN_1102;
      end
    end else begin
      rob_payload_77_tsc <= _GEN_1102;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4d == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_77_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_77_rob_idx <= _GEN_1230;
      end
    end else begin
      rob_payload_77_rob_idx <= _GEN_1230;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h4d == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_77_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_77_flits_fired <= _GEN_5841;
      end
    end else begin
      rob_payload_77_flits_fired <= _GEN_5841;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4e == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_78_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_78_tsc <= _GEN_1103;
      end
    end else begin
      rob_payload_78_tsc <= _GEN_1103;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4e == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_78_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_78_rob_idx <= _GEN_1231;
      end
    end else begin
      rob_payload_78_rob_idx <= _GEN_1231;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h4e == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_78_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_78_flits_fired <= _GEN_5842;
      end
    end else begin
      rob_payload_78_flits_fired <= _GEN_5842;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4f == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_79_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_79_tsc <= _GEN_1104;
      end
    end else begin
      rob_payload_79_tsc <= _GEN_1104;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4f == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_79_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_79_rob_idx <= _GEN_1232;
      end
    end else begin
      rob_payload_79_rob_idx <= _GEN_1232;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h4f == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_79_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_79_flits_fired <= _GEN_5843;
      end
    end else begin
      rob_payload_79_flits_fired <= _GEN_5843;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h50 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_80_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_80_tsc <= _GEN_1105;
      end
    end else begin
      rob_payload_80_tsc <= _GEN_1105;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h50 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_80_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_80_rob_idx <= _GEN_1233;
      end
    end else begin
      rob_payload_80_rob_idx <= _GEN_1233;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h50 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_80_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_80_flits_fired <= _GEN_5844;
      end
    end else begin
      rob_payload_80_flits_fired <= _GEN_5844;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h51 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_81_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_81_tsc <= _GEN_1106;
      end
    end else begin
      rob_payload_81_tsc <= _GEN_1106;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h51 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_81_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_81_rob_idx <= _GEN_1234;
      end
    end else begin
      rob_payload_81_rob_idx <= _GEN_1234;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h51 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_81_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_81_flits_fired <= _GEN_5845;
      end
    end else begin
      rob_payload_81_flits_fired <= _GEN_5845;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h52 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_82_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_82_tsc <= _GEN_1107;
      end
    end else begin
      rob_payload_82_tsc <= _GEN_1107;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h52 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_82_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_82_rob_idx <= _GEN_1235;
      end
    end else begin
      rob_payload_82_rob_idx <= _GEN_1235;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h52 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_82_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_82_flits_fired <= _GEN_5846;
      end
    end else begin
      rob_payload_82_flits_fired <= _GEN_5846;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h53 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_83_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_83_tsc <= _GEN_1108;
      end
    end else begin
      rob_payload_83_tsc <= _GEN_1108;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h53 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_83_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_83_rob_idx <= _GEN_1236;
      end
    end else begin
      rob_payload_83_rob_idx <= _GEN_1236;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h53 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_83_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_83_flits_fired <= _GEN_5847;
      end
    end else begin
      rob_payload_83_flits_fired <= _GEN_5847;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h54 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_84_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_84_tsc <= _GEN_1109;
      end
    end else begin
      rob_payload_84_tsc <= _GEN_1109;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h54 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_84_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_84_rob_idx <= _GEN_1237;
      end
    end else begin
      rob_payload_84_rob_idx <= _GEN_1237;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h54 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_84_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_84_flits_fired <= _GEN_5848;
      end
    end else begin
      rob_payload_84_flits_fired <= _GEN_5848;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h55 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_85_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_85_tsc <= _GEN_1110;
      end
    end else begin
      rob_payload_85_tsc <= _GEN_1110;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h55 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_85_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_85_rob_idx <= _GEN_1238;
      end
    end else begin
      rob_payload_85_rob_idx <= _GEN_1238;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h55 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_85_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_85_flits_fired <= _GEN_5849;
      end
    end else begin
      rob_payload_85_flits_fired <= _GEN_5849;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h56 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_86_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_86_tsc <= _GEN_1111;
      end
    end else begin
      rob_payload_86_tsc <= _GEN_1111;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h56 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_86_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_86_rob_idx <= _GEN_1239;
      end
    end else begin
      rob_payload_86_rob_idx <= _GEN_1239;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h56 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_86_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_86_flits_fired <= _GEN_5850;
      end
    end else begin
      rob_payload_86_flits_fired <= _GEN_5850;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h57 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_87_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_87_tsc <= _GEN_1112;
      end
    end else begin
      rob_payload_87_tsc <= _GEN_1112;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h57 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_87_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_87_rob_idx <= _GEN_1240;
      end
    end else begin
      rob_payload_87_rob_idx <= _GEN_1240;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h57 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_87_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_87_flits_fired <= _GEN_5851;
      end
    end else begin
      rob_payload_87_flits_fired <= _GEN_5851;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h58 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_88_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_88_tsc <= _GEN_1113;
      end
    end else begin
      rob_payload_88_tsc <= _GEN_1113;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h58 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_88_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_88_rob_idx <= _GEN_1241;
      end
    end else begin
      rob_payload_88_rob_idx <= _GEN_1241;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h58 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_88_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_88_flits_fired <= _GEN_5852;
      end
    end else begin
      rob_payload_88_flits_fired <= _GEN_5852;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h59 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_89_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_89_tsc <= _GEN_1114;
      end
    end else begin
      rob_payload_89_tsc <= _GEN_1114;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h59 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_89_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_89_rob_idx <= _GEN_1242;
      end
    end else begin
      rob_payload_89_rob_idx <= _GEN_1242;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h59 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_89_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_89_flits_fired <= _GEN_5853;
      end
    end else begin
      rob_payload_89_flits_fired <= _GEN_5853;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5a == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_90_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_90_tsc <= _GEN_1115;
      end
    end else begin
      rob_payload_90_tsc <= _GEN_1115;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5a == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_90_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_90_rob_idx <= _GEN_1243;
      end
    end else begin
      rob_payload_90_rob_idx <= _GEN_1243;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h5a == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_90_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_90_flits_fired <= _GEN_5854;
      end
    end else begin
      rob_payload_90_flits_fired <= _GEN_5854;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5b == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_91_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_91_tsc <= _GEN_1116;
      end
    end else begin
      rob_payload_91_tsc <= _GEN_1116;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5b == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_91_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_91_rob_idx <= _GEN_1244;
      end
    end else begin
      rob_payload_91_rob_idx <= _GEN_1244;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h5b == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_91_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_91_flits_fired <= _GEN_5855;
      end
    end else begin
      rob_payload_91_flits_fired <= _GEN_5855;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5c == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_92_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_92_tsc <= _GEN_1117;
      end
    end else begin
      rob_payload_92_tsc <= _GEN_1117;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5c == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_92_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_92_rob_idx <= _GEN_1245;
      end
    end else begin
      rob_payload_92_rob_idx <= _GEN_1245;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h5c == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_92_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_92_flits_fired <= _GEN_5856;
      end
    end else begin
      rob_payload_92_flits_fired <= _GEN_5856;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5d == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_93_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_93_tsc <= _GEN_1118;
      end
    end else begin
      rob_payload_93_tsc <= _GEN_1118;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5d == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_93_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_93_rob_idx <= _GEN_1246;
      end
    end else begin
      rob_payload_93_rob_idx <= _GEN_1246;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h5d == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_93_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_93_flits_fired <= _GEN_5857;
      end
    end else begin
      rob_payload_93_flits_fired <= _GEN_5857;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5e == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_94_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_94_tsc <= _GEN_1119;
      end
    end else begin
      rob_payload_94_tsc <= _GEN_1119;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5e == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_94_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_94_rob_idx <= _GEN_1247;
      end
    end else begin
      rob_payload_94_rob_idx <= _GEN_1247;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h5e == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_94_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_94_flits_fired <= _GEN_5858;
      end
    end else begin
      rob_payload_94_flits_fired <= _GEN_5858;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5f == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_95_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_95_tsc <= _GEN_1120;
      end
    end else begin
      rob_payload_95_tsc <= _GEN_1120;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5f == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_95_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_95_rob_idx <= _GEN_1248;
      end
    end else begin
      rob_payload_95_rob_idx <= _GEN_1248;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h5f == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_95_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_95_flits_fired <= _GEN_5859;
      end
    end else begin
      rob_payload_95_flits_fired <= _GEN_5859;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h60 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_96_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_96_tsc <= _GEN_1121;
      end
    end else begin
      rob_payload_96_tsc <= _GEN_1121;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h60 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_96_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_96_rob_idx <= _GEN_1249;
      end
    end else begin
      rob_payload_96_rob_idx <= _GEN_1249;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h60 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_96_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_96_flits_fired <= _GEN_5860;
      end
    end else begin
      rob_payload_96_flits_fired <= _GEN_5860;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h61 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_97_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_97_tsc <= _GEN_1122;
      end
    end else begin
      rob_payload_97_tsc <= _GEN_1122;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h61 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_97_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_97_rob_idx <= _GEN_1250;
      end
    end else begin
      rob_payload_97_rob_idx <= _GEN_1250;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h61 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_97_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_97_flits_fired <= _GEN_5861;
      end
    end else begin
      rob_payload_97_flits_fired <= _GEN_5861;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h62 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_98_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_98_tsc <= _GEN_1123;
      end
    end else begin
      rob_payload_98_tsc <= _GEN_1123;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h62 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_98_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_98_rob_idx <= _GEN_1251;
      end
    end else begin
      rob_payload_98_rob_idx <= _GEN_1251;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h62 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_98_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_98_flits_fired <= _GEN_5862;
      end
    end else begin
      rob_payload_98_flits_fired <= _GEN_5862;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h63 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_99_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_99_tsc <= _GEN_1124;
      end
    end else begin
      rob_payload_99_tsc <= _GEN_1124;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h63 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_99_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_99_rob_idx <= _GEN_1252;
      end
    end else begin
      rob_payload_99_rob_idx <= _GEN_1252;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h63 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_99_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_99_flits_fired <= _GEN_5863;
      end
    end else begin
      rob_payload_99_flits_fired <= _GEN_5863;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h64 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_100_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_100_tsc <= _GEN_1125;
      end
    end else begin
      rob_payload_100_tsc <= _GEN_1125;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h64 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_100_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_100_rob_idx <= _GEN_1253;
      end
    end else begin
      rob_payload_100_rob_idx <= _GEN_1253;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h64 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_100_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_100_flits_fired <= _GEN_5864;
      end
    end else begin
      rob_payload_100_flits_fired <= _GEN_5864;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h65 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_101_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_101_tsc <= _GEN_1126;
      end
    end else begin
      rob_payload_101_tsc <= _GEN_1126;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h65 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_101_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_101_rob_idx <= _GEN_1254;
      end
    end else begin
      rob_payload_101_rob_idx <= _GEN_1254;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h65 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_101_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_101_flits_fired <= _GEN_5865;
      end
    end else begin
      rob_payload_101_flits_fired <= _GEN_5865;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h66 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_102_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_102_tsc <= _GEN_1127;
      end
    end else begin
      rob_payload_102_tsc <= _GEN_1127;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h66 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_102_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_102_rob_idx <= _GEN_1255;
      end
    end else begin
      rob_payload_102_rob_idx <= _GEN_1255;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h66 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_102_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_102_flits_fired <= _GEN_5866;
      end
    end else begin
      rob_payload_102_flits_fired <= _GEN_5866;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h67 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_103_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_103_tsc <= _GEN_1128;
      end
    end else begin
      rob_payload_103_tsc <= _GEN_1128;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h67 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_103_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_103_rob_idx <= _GEN_1256;
      end
    end else begin
      rob_payload_103_rob_idx <= _GEN_1256;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h67 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_103_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_103_flits_fired <= _GEN_5867;
      end
    end else begin
      rob_payload_103_flits_fired <= _GEN_5867;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h68 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_104_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_104_tsc <= _GEN_1129;
      end
    end else begin
      rob_payload_104_tsc <= _GEN_1129;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h68 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_104_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_104_rob_idx <= _GEN_1257;
      end
    end else begin
      rob_payload_104_rob_idx <= _GEN_1257;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h68 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_104_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_104_flits_fired <= _GEN_5868;
      end
    end else begin
      rob_payload_104_flits_fired <= _GEN_5868;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h69 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_105_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_105_tsc <= _GEN_1130;
      end
    end else begin
      rob_payload_105_tsc <= _GEN_1130;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h69 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_105_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_105_rob_idx <= _GEN_1258;
      end
    end else begin
      rob_payload_105_rob_idx <= _GEN_1258;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h69 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_105_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_105_flits_fired <= _GEN_5869;
      end
    end else begin
      rob_payload_105_flits_fired <= _GEN_5869;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6a == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_106_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_106_tsc <= _GEN_1131;
      end
    end else begin
      rob_payload_106_tsc <= _GEN_1131;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6a == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_106_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_106_rob_idx <= _GEN_1259;
      end
    end else begin
      rob_payload_106_rob_idx <= _GEN_1259;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h6a == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_106_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_106_flits_fired <= _GEN_5870;
      end
    end else begin
      rob_payload_106_flits_fired <= _GEN_5870;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6b == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_107_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_107_tsc <= _GEN_1132;
      end
    end else begin
      rob_payload_107_tsc <= _GEN_1132;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6b == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_107_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_107_rob_idx <= _GEN_1260;
      end
    end else begin
      rob_payload_107_rob_idx <= _GEN_1260;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h6b == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_107_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_107_flits_fired <= _GEN_5871;
      end
    end else begin
      rob_payload_107_flits_fired <= _GEN_5871;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6c == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_108_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_108_tsc <= _GEN_1133;
      end
    end else begin
      rob_payload_108_tsc <= _GEN_1133;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6c == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_108_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_108_rob_idx <= _GEN_1261;
      end
    end else begin
      rob_payload_108_rob_idx <= _GEN_1261;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h6c == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_108_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_108_flits_fired <= _GEN_5872;
      end
    end else begin
      rob_payload_108_flits_fired <= _GEN_5872;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6d == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_109_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_109_tsc <= _GEN_1134;
      end
    end else begin
      rob_payload_109_tsc <= _GEN_1134;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6d == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_109_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_109_rob_idx <= _GEN_1262;
      end
    end else begin
      rob_payload_109_rob_idx <= _GEN_1262;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h6d == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_109_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_109_flits_fired <= _GEN_5873;
      end
    end else begin
      rob_payload_109_flits_fired <= _GEN_5873;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6e == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_110_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_110_tsc <= _GEN_1135;
      end
    end else begin
      rob_payload_110_tsc <= _GEN_1135;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6e == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_110_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_110_rob_idx <= _GEN_1263;
      end
    end else begin
      rob_payload_110_rob_idx <= _GEN_1263;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h6e == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_110_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_110_flits_fired <= _GEN_5874;
      end
    end else begin
      rob_payload_110_flits_fired <= _GEN_5874;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6f == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_111_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_111_tsc <= _GEN_1136;
      end
    end else begin
      rob_payload_111_tsc <= _GEN_1136;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6f == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_111_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_111_rob_idx <= _GEN_1264;
      end
    end else begin
      rob_payload_111_rob_idx <= _GEN_1264;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h6f == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_111_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_111_flits_fired <= _GEN_5875;
      end
    end else begin
      rob_payload_111_flits_fired <= _GEN_5875;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h70 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_112_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_112_tsc <= _GEN_1137;
      end
    end else begin
      rob_payload_112_tsc <= _GEN_1137;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h70 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_112_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_112_rob_idx <= _GEN_1265;
      end
    end else begin
      rob_payload_112_rob_idx <= _GEN_1265;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h70 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_112_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_112_flits_fired <= _GEN_5876;
      end
    end else begin
      rob_payload_112_flits_fired <= _GEN_5876;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h71 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_113_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_113_tsc <= _GEN_1138;
      end
    end else begin
      rob_payload_113_tsc <= _GEN_1138;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h71 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_113_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_113_rob_idx <= _GEN_1266;
      end
    end else begin
      rob_payload_113_rob_idx <= _GEN_1266;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h71 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_113_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_113_flits_fired <= _GEN_5877;
      end
    end else begin
      rob_payload_113_flits_fired <= _GEN_5877;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h72 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_114_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_114_tsc <= _GEN_1139;
      end
    end else begin
      rob_payload_114_tsc <= _GEN_1139;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h72 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_114_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_114_rob_idx <= _GEN_1267;
      end
    end else begin
      rob_payload_114_rob_idx <= _GEN_1267;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h72 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_114_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_114_flits_fired <= _GEN_5878;
      end
    end else begin
      rob_payload_114_flits_fired <= _GEN_5878;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h73 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_115_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_115_tsc <= _GEN_1140;
      end
    end else begin
      rob_payload_115_tsc <= _GEN_1140;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h73 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_115_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_115_rob_idx <= _GEN_1268;
      end
    end else begin
      rob_payload_115_rob_idx <= _GEN_1268;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h73 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_115_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_115_flits_fired <= _GEN_5879;
      end
    end else begin
      rob_payload_115_flits_fired <= _GEN_5879;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h74 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_116_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_116_tsc <= _GEN_1141;
      end
    end else begin
      rob_payload_116_tsc <= _GEN_1141;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h74 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_116_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_116_rob_idx <= _GEN_1269;
      end
    end else begin
      rob_payload_116_rob_idx <= _GEN_1269;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h74 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_116_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_116_flits_fired <= _GEN_5880;
      end
    end else begin
      rob_payload_116_flits_fired <= _GEN_5880;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h75 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_117_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_117_tsc <= _GEN_1142;
      end
    end else begin
      rob_payload_117_tsc <= _GEN_1142;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h75 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_117_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_117_rob_idx <= _GEN_1270;
      end
    end else begin
      rob_payload_117_rob_idx <= _GEN_1270;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h75 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_117_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_117_flits_fired <= _GEN_5881;
      end
    end else begin
      rob_payload_117_flits_fired <= _GEN_5881;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h76 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_118_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_118_tsc <= _GEN_1143;
      end
    end else begin
      rob_payload_118_tsc <= _GEN_1143;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h76 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_118_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_118_rob_idx <= _GEN_1271;
      end
    end else begin
      rob_payload_118_rob_idx <= _GEN_1271;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h76 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_118_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_118_flits_fired <= _GEN_5882;
      end
    end else begin
      rob_payload_118_flits_fired <= _GEN_5882;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h77 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_119_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_119_tsc <= _GEN_1144;
      end
    end else begin
      rob_payload_119_tsc <= _GEN_1144;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h77 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_119_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_119_rob_idx <= _GEN_1272;
      end
    end else begin
      rob_payload_119_rob_idx <= _GEN_1272;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h77 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_119_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_119_flits_fired <= _GEN_5883;
      end
    end else begin
      rob_payload_119_flits_fired <= _GEN_5883;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h78 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_120_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_120_tsc <= _GEN_1145;
      end
    end else begin
      rob_payload_120_tsc <= _GEN_1145;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h78 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_120_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_120_rob_idx <= _GEN_1273;
      end
    end else begin
      rob_payload_120_rob_idx <= _GEN_1273;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h78 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_120_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_120_flits_fired <= _GEN_5884;
      end
    end else begin
      rob_payload_120_flits_fired <= _GEN_5884;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h79 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_121_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_121_tsc <= _GEN_1146;
      end
    end else begin
      rob_payload_121_tsc <= _GEN_1146;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h79 == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_121_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_121_rob_idx <= _GEN_1274;
      end
    end else begin
      rob_payload_121_rob_idx <= _GEN_1274;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h79 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_121_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_121_flits_fired <= _GEN_5885;
      end
    end else begin
      rob_payload_121_flits_fired <= _GEN_5885;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7a == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_122_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_122_tsc <= _GEN_1147;
      end
    end else begin
      rob_payload_122_tsc <= _GEN_1147;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7a == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_122_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_122_rob_idx <= _GEN_1275;
      end
    end else begin
      rob_payload_122_rob_idx <= _GEN_1275;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h7a == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_122_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_122_flits_fired <= _GEN_5886;
      end
    end else begin
      rob_payload_122_flits_fired <= _GEN_5886;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7b == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_123_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_123_tsc <= _GEN_1148;
      end
    end else begin
      rob_payload_123_tsc <= _GEN_1148;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7b == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_123_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_123_rob_idx <= _GEN_1276;
      end
    end else begin
      rob_payload_123_rob_idx <= _GEN_1276;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h7b == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_123_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_123_flits_fired <= _GEN_5887;
      end
    end else begin
      rob_payload_123_flits_fired <= _GEN_5887;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7c == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_124_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_124_tsc <= _GEN_1149;
      end
    end else begin
      rob_payload_124_tsc <= _GEN_1149;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7c == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_124_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_124_rob_idx <= _GEN_1277;
      end
    end else begin
      rob_payload_124_rob_idx <= _GEN_1277;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h7c == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_124_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_124_flits_fired <= _GEN_5888;
      end
    end else begin
      rob_payload_124_flits_fired <= _GEN_5888;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7d == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_125_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_125_tsc <= _GEN_1150;
      end
    end else begin
      rob_payload_125_tsc <= _GEN_1150;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7d == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_125_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_125_rob_idx <= _GEN_1278;
      end
    end else begin
      rob_payload_125_rob_idx <= _GEN_1278;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h7d == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_125_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_125_flits_fired <= _GEN_5889;
      end
    end else begin
      rob_payload_125_flits_fired <= _GEN_5889;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7e == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_126_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_126_tsc <= _GEN_1151;
      end
    end else begin
      rob_payload_126_tsc <= _GEN_1151;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7e == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_126_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_126_rob_idx <= _GEN_1279;
      end
    end else begin
      rob_payload_126_rob_idx <= _GEN_1279;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h7e == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_126_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_126_flits_fired <= _GEN_5890;
      end
    end else begin
      rob_payload_126_flits_fired <= _GEN_5890;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7f == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_127_tsc <= _rob_payload_WIRE_3[63:32]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_127_tsc <= _GEN_1152;
      end
    end else begin
      rob_payload_127_tsc <= _GEN_1152;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7f == rob_alloc_ids_1) begin // @[TestHarness.scala 179:36]
        rob_payload_127_rob_idx <= _rob_payload_WIRE_3[31:16]; // @[TestHarness.scala 179:36]
      end else begin
        rob_payload_127_rob_idx <= _GEN_1280;
      end
    end else begin
      rob_payload_127_rob_idx <= _GEN_1280;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h7f == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 214:40]
        rob_payload_127_flits_fired <= _rob_payload_flits_fired_T_5; // @[TestHarness.scala 214:40]
      end else begin
        rob_payload_127_flits_fired <= _GEN_5891;
      end
    end else begin
      rob_payload_127_flits_fired <= _GEN_5891;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h0 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_0 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_0 <= _GEN_1409;
      end
    end else begin
      rob_egress_id_0 <= _GEN_1409;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_1 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_1 <= _GEN_1410;
      end
    end else begin
      rob_egress_id_1 <= _GEN_1410;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_2 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_2 <= _GEN_1411;
      end
    end else begin
      rob_egress_id_2 <= _GEN_1411;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_3 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_3 <= _GEN_1412;
      end
    end else begin
      rob_egress_id_3 <= _GEN_1412;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_4 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_4 <= _GEN_1413;
      end
    end else begin
      rob_egress_id_4 <= _GEN_1413;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_5 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_5 <= _GEN_1414;
      end
    end else begin
      rob_egress_id_5 <= _GEN_1414;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_6 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_6 <= _GEN_1415;
      end
    end else begin
      rob_egress_id_6 <= _GEN_1415;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_7 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_7 <= _GEN_1416;
      end
    end else begin
      rob_egress_id_7 <= _GEN_1416;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h8 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_8 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_8 <= _GEN_1417;
      end
    end else begin
      rob_egress_id_8 <= _GEN_1417;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h9 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_9 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_9 <= _GEN_1418;
      end
    end else begin
      rob_egress_id_9 <= _GEN_1418;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'ha == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_10 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_10 <= _GEN_1419;
      end
    end else begin
      rob_egress_id_10 <= _GEN_1419;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hb == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_11 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_11 <= _GEN_1420;
      end
    end else begin
      rob_egress_id_11 <= _GEN_1420;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hc == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_12 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_12 <= _GEN_1421;
      end
    end else begin
      rob_egress_id_12 <= _GEN_1421;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hd == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_13 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_13 <= _GEN_1422;
      end
    end else begin
      rob_egress_id_13 <= _GEN_1422;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'he == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_14 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_14 <= _GEN_1423;
      end
    end else begin
      rob_egress_id_14 <= _GEN_1423;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hf == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_15 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_15 <= _GEN_1424;
      end
    end else begin
      rob_egress_id_15 <= _GEN_1424;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h10 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_16 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_16 <= _GEN_1425;
      end
    end else begin
      rob_egress_id_16 <= _GEN_1425;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h11 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_17 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_17 <= _GEN_1426;
      end
    end else begin
      rob_egress_id_17 <= _GEN_1426;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h12 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_18 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_18 <= _GEN_1427;
      end
    end else begin
      rob_egress_id_18 <= _GEN_1427;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h13 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_19 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_19 <= _GEN_1428;
      end
    end else begin
      rob_egress_id_19 <= _GEN_1428;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h14 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_20 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_20 <= _GEN_1429;
      end
    end else begin
      rob_egress_id_20 <= _GEN_1429;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h15 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_21 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_21 <= _GEN_1430;
      end
    end else begin
      rob_egress_id_21 <= _GEN_1430;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h16 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_22 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_22 <= _GEN_1431;
      end
    end else begin
      rob_egress_id_22 <= _GEN_1431;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h17 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_23 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_23 <= _GEN_1432;
      end
    end else begin
      rob_egress_id_23 <= _GEN_1432;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h18 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_24 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_24 <= _GEN_1433;
      end
    end else begin
      rob_egress_id_24 <= _GEN_1433;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h19 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_25 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_25 <= _GEN_1434;
      end
    end else begin
      rob_egress_id_25 <= _GEN_1434;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1a == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_26 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_26 <= _GEN_1435;
      end
    end else begin
      rob_egress_id_26 <= _GEN_1435;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1b == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_27 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_27 <= _GEN_1436;
      end
    end else begin
      rob_egress_id_27 <= _GEN_1436;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1c == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_28 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_28 <= _GEN_1437;
      end
    end else begin
      rob_egress_id_28 <= _GEN_1437;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1d == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_29 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_29 <= _GEN_1438;
      end
    end else begin
      rob_egress_id_29 <= _GEN_1438;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1e == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_30 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_30 <= _GEN_1439;
      end
    end else begin
      rob_egress_id_30 <= _GEN_1439;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1f == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_31 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_31 <= _GEN_1440;
      end
    end else begin
      rob_egress_id_31 <= _GEN_1440;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h20 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_32 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_32 <= _GEN_1441;
      end
    end else begin
      rob_egress_id_32 <= _GEN_1441;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h21 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_33 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_33 <= _GEN_1442;
      end
    end else begin
      rob_egress_id_33 <= _GEN_1442;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h22 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_34 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_34 <= _GEN_1443;
      end
    end else begin
      rob_egress_id_34 <= _GEN_1443;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h23 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_35 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_35 <= _GEN_1444;
      end
    end else begin
      rob_egress_id_35 <= _GEN_1444;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h24 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_36 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_36 <= _GEN_1445;
      end
    end else begin
      rob_egress_id_36 <= _GEN_1445;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h25 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_37 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_37 <= _GEN_1446;
      end
    end else begin
      rob_egress_id_37 <= _GEN_1446;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h26 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_38 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_38 <= _GEN_1447;
      end
    end else begin
      rob_egress_id_38 <= _GEN_1447;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h27 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_39 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_39 <= _GEN_1448;
      end
    end else begin
      rob_egress_id_39 <= _GEN_1448;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h28 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_40 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_40 <= _GEN_1449;
      end
    end else begin
      rob_egress_id_40 <= _GEN_1449;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h29 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_41 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_41 <= _GEN_1450;
      end
    end else begin
      rob_egress_id_41 <= _GEN_1450;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2a == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_42 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_42 <= _GEN_1451;
      end
    end else begin
      rob_egress_id_42 <= _GEN_1451;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2b == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_43 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_43 <= _GEN_1452;
      end
    end else begin
      rob_egress_id_43 <= _GEN_1452;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2c == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_44 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_44 <= _GEN_1453;
      end
    end else begin
      rob_egress_id_44 <= _GEN_1453;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2d == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_45 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_45 <= _GEN_1454;
      end
    end else begin
      rob_egress_id_45 <= _GEN_1454;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2e == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_46 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_46 <= _GEN_1455;
      end
    end else begin
      rob_egress_id_46 <= _GEN_1455;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2f == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_47 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_47 <= _GEN_1456;
      end
    end else begin
      rob_egress_id_47 <= _GEN_1456;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h30 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_48 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_48 <= _GEN_1457;
      end
    end else begin
      rob_egress_id_48 <= _GEN_1457;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h31 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_49 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_49 <= _GEN_1458;
      end
    end else begin
      rob_egress_id_49 <= _GEN_1458;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h32 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_50 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_50 <= _GEN_1459;
      end
    end else begin
      rob_egress_id_50 <= _GEN_1459;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h33 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_51 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_51 <= _GEN_1460;
      end
    end else begin
      rob_egress_id_51 <= _GEN_1460;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h34 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_52 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_52 <= _GEN_1461;
      end
    end else begin
      rob_egress_id_52 <= _GEN_1461;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h35 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_53 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_53 <= _GEN_1462;
      end
    end else begin
      rob_egress_id_53 <= _GEN_1462;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h36 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_54 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_54 <= _GEN_1463;
      end
    end else begin
      rob_egress_id_54 <= _GEN_1463;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h37 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_55 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_55 <= _GEN_1464;
      end
    end else begin
      rob_egress_id_55 <= _GEN_1464;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h38 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_56 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_56 <= _GEN_1465;
      end
    end else begin
      rob_egress_id_56 <= _GEN_1465;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h39 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_57 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_57 <= _GEN_1466;
      end
    end else begin
      rob_egress_id_57 <= _GEN_1466;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3a == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_58 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_58 <= _GEN_1467;
      end
    end else begin
      rob_egress_id_58 <= _GEN_1467;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3b == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_59 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_59 <= _GEN_1468;
      end
    end else begin
      rob_egress_id_59 <= _GEN_1468;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3c == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_60 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_60 <= _GEN_1469;
      end
    end else begin
      rob_egress_id_60 <= _GEN_1469;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3d == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_61 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_61 <= _GEN_1470;
      end
    end else begin
      rob_egress_id_61 <= _GEN_1470;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3e == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_62 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_62 <= _GEN_1471;
      end
    end else begin
      rob_egress_id_62 <= _GEN_1471;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3f == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_63 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_63 <= _GEN_1472;
      end
    end else begin
      rob_egress_id_63 <= _GEN_1472;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h40 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_64 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_64 <= _GEN_1473;
      end
    end else begin
      rob_egress_id_64 <= _GEN_1473;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h41 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_65 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_65 <= _GEN_1474;
      end
    end else begin
      rob_egress_id_65 <= _GEN_1474;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h42 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_66 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_66 <= _GEN_1475;
      end
    end else begin
      rob_egress_id_66 <= _GEN_1475;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h43 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_67 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_67 <= _GEN_1476;
      end
    end else begin
      rob_egress_id_67 <= _GEN_1476;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h44 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_68 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_68 <= _GEN_1477;
      end
    end else begin
      rob_egress_id_68 <= _GEN_1477;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h45 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_69 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_69 <= _GEN_1478;
      end
    end else begin
      rob_egress_id_69 <= _GEN_1478;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h46 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_70 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_70 <= _GEN_1479;
      end
    end else begin
      rob_egress_id_70 <= _GEN_1479;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h47 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_71 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_71 <= _GEN_1480;
      end
    end else begin
      rob_egress_id_71 <= _GEN_1480;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h48 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_72 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_72 <= _GEN_1481;
      end
    end else begin
      rob_egress_id_72 <= _GEN_1481;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h49 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_73 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_73 <= _GEN_1482;
      end
    end else begin
      rob_egress_id_73 <= _GEN_1482;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4a == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_74 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_74 <= _GEN_1483;
      end
    end else begin
      rob_egress_id_74 <= _GEN_1483;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4b == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_75 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_75 <= _GEN_1484;
      end
    end else begin
      rob_egress_id_75 <= _GEN_1484;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4c == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_76 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_76 <= _GEN_1485;
      end
    end else begin
      rob_egress_id_76 <= _GEN_1485;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4d == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_77 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_77 <= _GEN_1486;
      end
    end else begin
      rob_egress_id_77 <= _GEN_1486;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4e == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_78 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_78 <= _GEN_1487;
      end
    end else begin
      rob_egress_id_78 <= _GEN_1487;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4f == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_79 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_79 <= _GEN_1488;
      end
    end else begin
      rob_egress_id_79 <= _GEN_1488;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h50 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_80 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_80 <= _GEN_1489;
      end
    end else begin
      rob_egress_id_80 <= _GEN_1489;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h51 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_81 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_81 <= _GEN_1490;
      end
    end else begin
      rob_egress_id_81 <= _GEN_1490;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h52 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_82 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_82 <= _GEN_1491;
      end
    end else begin
      rob_egress_id_82 <= _GEN_1491;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h53 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_83 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_83 <= _GEN_1492;
      end
    end else begin
      rob_egress_id_83 <= _GEN_1492;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h54 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_84 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_84 <= _GEN_1493;
      end
    end else begin
      rob_egress_id_84 <= _GEN_1493;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h55 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_85 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_85 <= _GEN_1494;
      end
    end else begin
      rob_egress_id_85 <= _GEN_1494;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h56 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_86 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_86 <= _GEN_1495;
      end
    end else begin
      rob_egress_id_86 <= _GEN_1495;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h57 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_87 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_87 <= _GEN_1496;
      end
    end else begin
      rob_egress_id_87 <= _GEN_1496;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h58 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_88 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_88 <= _GEN_1497;
      end
    end else begin
      rob_egress_id_88 <= _GEN_1497;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h59 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_89 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_89 <= _GEN_1498;
      end
    end else begin
      rob_egress_id_89 <= _GEN_1498;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5a == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_90 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_90 <= _GEN_1499;
      end
    end else begin
      rob_egress_id_90 <= _GEN_1499;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5b == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_91 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_91 <= _GEN_1500;
      end
    end else begin
      rob_egress_id_91 <= _GEN_1500;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5c == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_92 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_92 <= _GEN_1501;
      end
    end else begin
      rob_egress_id_92 <= _GEN_1501;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5d == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_93 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_93 <= _GEN_1502;
      end
    end else begin
      rob_egress_id_93 <= _GEN_1502;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5e == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_94 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_94 <= _GEN_1503;
      end
    end else begin
      rob_egress_id_94 <= _GEN_1503;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5f == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_95 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_95 <= _GEN_1504;
      end
    end else begin
      rob_egress_id_95 <= _GEN_1504;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h60 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_96 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_96 <= _GEN_1505;
      end
    end else begin
      rob_egress_id_96 <= _GEN_1505;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h61 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_97 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_97 <= _GEN_1506;
      end
    end else begin
      rob_egress_id_97 <= _GEN_1506;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h62 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_98 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_98 <= _GEN_1507;
      end
    end else begin
      rob_egress_id_98 <= _GEN_1507;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h63 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_99 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_99 <= _GEN_1508;
      end
    end else begin
      rob_egress_id_99 <= _GEN_1508;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h64 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_100 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_100 <= _GEN_1509;
      end
    end else begin
      rob_egress_id_100 <= _GEN_1509;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h65 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_101 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_101 <= _GEN_1510;
      end
    end else begin
      rob_egress_id_101 <= _GEN_1510;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h66 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_102 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_102 <= _GEN_1511;
      end
    end else begin
      rob_egress_id_102 <= _GEN_1511;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h67 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_103 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_103 <= _GEN_1512;
      end
    end else begin
      rob_egress_id_103 <= _GEN_1512;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h68 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_104 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_104 <= _GEN_1513;
      end
    end else begin
      rob_egress_id_104 <= _GEN_1513;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h69 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_105 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_105 <= _GEN_1514;
      end
    end else begin
      rob_egress_id_105 <= _GEN_1514;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6a == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_106 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_106 <= _GEN_1515;
      end
    end else begin
      rob_egress_id_106 <= _GEN_1515;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6b == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_107 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_107 <= _GEN_1516;
      end
    end else begin
      rob_egress_id_107 <= _GEN_1516;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6c == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_108 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_108 <= _GEN_1517;
      end
    end else begin
      rob_egress_id_108 <= _GEN_1517;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6d == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_109 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_109 <= _GEN_1518;
      end
    end else begin
      rob_egress_id_109 <= _GEN_1518;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6e == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_110 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_110 <= _GEN_1519;
      end
    end else begin
      rob_egress_id_110 <= _GEN_1519;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6f == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_111 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_111 <= _GEN_1520;
      end
    end else begin
      rob_egress_id_111 <= _GEN_1520;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h70 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_112 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_112 <= _GEN_1521;
      end
    end else begin
      rob_egress_id_112 <= _GEN_1521;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h71 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_113 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_113 <= _GEN_1522;
      end
    end else begin
      rob_egress_id_113 <= _GEN_1522;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h72 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_114 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_114 <= _GEN_1523;
      end
    end else begin
      rob_egress_id_114 <= _GEN_1523;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h73 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_115 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_115 <= _GEN_1524;
      end
    end else begin
      rob_egress_id_115 <= _GEN_1524;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h74 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_116 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_116 <= _GEN_1525;
      end
    end else begin
      rob_egress_id_116 <= _GEN_1525;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h75 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_117 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_117 <= _GEN_1526;
      end
    end else begin
      rob_egress_id_117 <= _GEN_1526;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h76 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_118 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_118 <= _GEN_1527;
      end
    end else begin
      rob_egress_id_118 <= _GEN_1527;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h77 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_119 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_119 <= _GEN_1528;
      end
    end else begin
      rob_egress_id_119 <= _GEN_1528;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h78 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_120 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_120 <= _GEN_1529;
      end
    end else begin
      rob_egress_id_120 <= _GEN_1529;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h79 == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_121 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_121 <= _GEN_1530;
      end
    end else begin
      rob_egress_id_121 <= _GEN_1530;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7a == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_122 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_122 <= _GEN_1531;
      end
    end else begin
      rob_egress_id_122 <= _GEN_1531;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7b == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_123 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_123 <= _GEN_1532;
      end
    end else begin
      rob_egress_id_123 <= _GEN_1532;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7c == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_124 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_124 <= _GEN_1533;
      end
    end else begin
      rob_egress_id_124 <= _GEN_1533;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7d == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_125 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_125 <= _GEN_1534;
      end
    end else begin
      rob_egress_id_125 <= _GEN_1534;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7e == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_126 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_126 <= _GEN_1535;
      end
    end else begin
      rob_egress_id_126 <= _GEN_1535;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7f == rob_alloc_ids_1) begin // @[TestHarness.scala 180:36]
        rob_egress_id_127 <= igen_1_io_out_bits_egress_id; // @[TestHarness.scala 180:36]
      end else begin
        rob_egress_id_127 <= _GEN_1536;
      end
    end else begin
      rob_egress_id_127 <= _GEN_1536;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_0 <= _GEN_2561;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h0 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_0 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_1 <= _GEN_2562;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_1 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_2 <= _GEN_2563;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_2 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_3 <= _GEN_2564;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_3 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_4 <= _GEN_2565;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_4 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_5 <= _GEN_2566;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_5 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_6 <= _GEN_2567;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_6 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_7 <= _GEN_2568;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_7 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_8 <= _GEN_2569;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h8 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_8 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_9 <= _GEN_2570;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h9 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_9 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_10 <= _GEN_2571;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'ha == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_10 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_11 <= _GEN_2572;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hb == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_11 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_12 <= _GEN_2573;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hc == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_12 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_13 <= _GEN_2574;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hd == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_13 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_14 <= _GEN_2575;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'he == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_14 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_15 <= _GEN_2576;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hf == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_15 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_16 <= _GEN_2577;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h10 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_16 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_17 <= _GEN_2578;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h11 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_17 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_18 <= _GEN_2579;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h12 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_18 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_19 <= _GEN_2580;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h13 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_19 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_20 <= _GEN_2581;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h14 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_20 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_21 <= _GEN_2582;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h15 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_21 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_22 <= _GEN_2583;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h16 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_22 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_23 <= _GEN_2584;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h17 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_23 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_24 <= _GEN_2585;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h18 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_24 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_25 <= _GEN_2586;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h19 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_25 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_26 <= _GEN_2587;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1a == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_26 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_27 <= _GEN_2588;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1b == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_27 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_28 <= _GEN_2589;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1c == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_28 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_29 <= _GEN_2590;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1d == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_29 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_30 <= _GEN_2591;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1e == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_30 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_31 <= _GEN_2592;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1f == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_31 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_32 <= _GEN_2593;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h20 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_32 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_33 <= _GEN_2594;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h21 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_33 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_34 <= _GEN_2595;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h22 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_34 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_35 <= _GEN_2596;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h23 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_35 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_36 <= _GEN_2597;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h24 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_36 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_37 <= _GEN_2598;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h25 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_37 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_38 <= _GEN_2599;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h26 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_38 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_39 <= _GEN_2600;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h27 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_39 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_40 <= _GEN_2601;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h28 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_40 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_41 <= _GEN_2602;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h29 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_41 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_42 <= _GEN_2603;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2a == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_42 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_43 <= _GEN_2604;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2b == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_43 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_44 <= _GEN_2605;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2c == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_44 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_45 <= _GEN_2606;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2d == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_45 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_46 <= _GEN_2607;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2e == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_46 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_47 <= _GEN_2608;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2f == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_47 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_48 <= _GEN_2609;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h30 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_48 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_49 <= _GEN_2610;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h31 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_49 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_50 <= _GEN_2611;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h32 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_50 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_51 <= _GEN_2612;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h33 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_51 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_52 <= _GEN_2613;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h34 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_52 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_53 <= _GEN_2614;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h35 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_53 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_54 <= _GEN_2615;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h36 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_54 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_55 <= _GEN_2616;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h37 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_55 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_56 <= _GEN_2617;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h38 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_56 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_57 <= _GEN_2618;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h39 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_57 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_58 <= _GEN_2619;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3a == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_58 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_59 <= _GEN_2620;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3b == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_59 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_60 <= _GEN_2621;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3c == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_60 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_61 <= _GEN_2622;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3d == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_61 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_62 <= _GEN_2623;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3e == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_62 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_63 <= _GEN_2624;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3f == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_63 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_64 <= _GEN_2625;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h40 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_64 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_65 <= _GEN_2626;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h41 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_65 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_66 <= _GEN_2627;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h42 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_66 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_67 <= _GEN_2628;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h43 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_67 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_68 <= _GEN_2629;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h44 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_68 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_69 <= _GEN_2630;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h45 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_69 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_70 <= _GEN_2631;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h46 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_70 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_71 <= _GEN_2632;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h47 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_71 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_72 <= _GEN_2633;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h48 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_72 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_73 <= _GEN_2634;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h49 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_73 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_74 <= _GEN_2635;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4a == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_74 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_75 <= _GEN_2636;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4b == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_75 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_76 <= _GEN_2637;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4c == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_76 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_77 <= _GEN_2638;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4d == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_77 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_78 <= _GEN_2639;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4e == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_78 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_79 <= _GEN_2640;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4f == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_79 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_80 <= _GEN_2641;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h50 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_80 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_81 <= _GEN_2642;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h51 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_81 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_82 <= _GEN_2643;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h52 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_82 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_83 <= _GEN_2644;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h53 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_83 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_84 <= _GEN_2645;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h54 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_84 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_85 <= _GEN_2646;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h55 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_85 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_86 <= _GEN_2647;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h56 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_86 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_87 <= _GEN_2648;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h57 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_87 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_88 <= _GEN_2649;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h58 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_88 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_89 <= _GEN_2650;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h59 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_89 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_90 <= _GEN_2651;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5a == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_90 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_91 <= _GEN_2652;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5b == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_91 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_92 <= _GEN_2653;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5c == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_92 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_93 <= _GEN_2654;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5d == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_93 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_94 <= _GEN_2655;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5e == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_94 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_95 <= _GEN_2656;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5f == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_95 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_96 <= _GEN_2657;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h60 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_96 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_97 <= _GEN_2658;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h61 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_97 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_98 <= _GEN_2659;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h62 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_98 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_99 <= _GEN_2660;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h63 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_99 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_100 <= _GEN_2661;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h64 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_100 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_101 <= _GEN_2662;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h65 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_101 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_102 <= _GEN_2663;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h66 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_102 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_103 <= _GEN_2664;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h67 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_103 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_104 <= _GEN_2665;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h68 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_104 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_105 <= _GEN_2666;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h69 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_105 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_106 <= _GEN_2667;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6a == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_106 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_107 <= _GEN_2668;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6b == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_107 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_108 <= _GEN_2669;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6c == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_108 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_109 <= _GEN_2670;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6d == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_109 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_110 <= _GEN_2671;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6e == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_110 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_111 <= _GEN_2672;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6f == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_111 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_112 <= _GEN_2673;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h70 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_112 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_113 <= _GEN_2674;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h71 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_113 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_114 <= _GEN_2675;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h72 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_114 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_115 <= _GEN_2676;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h73 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_115 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_116 <= _GEN_2677;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h74 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_116 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_117 <= _GEN_2678;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h75 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_117 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_118 <= _GEN_2679;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h76 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_118 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_119 <= _GEN_2680;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h77 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_119 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_120 <= _GEN_2681;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h78 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_120 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_121 <= _GEN_2682;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h79 == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_121 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_122 <= _GEN_2683;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7a == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_122 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_123 <= _GEN_2684;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7b == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_123 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_124 <= _GEN_2685;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7c == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_124 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_125 <= _GEN_2686;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7d == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_125 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_126 <= _GEN_2687;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7e == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_126 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      rob_ingress_id_127 <= _GEN_2688;
    end else if (igen_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7f == rob_alloc_ids_0) begin // @[TestHarness.scala 181:36]
        rob_ingress_id_127 <= 1'h0; // @[TestHarness.scala 181:36]
      end
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h0 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_0 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_0 <= _GEN_1665;
      end
    end else begin
      rob_n_flits_0 <= _GEN_1665;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_1 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_1 <= _GEN_1666;
      end
    end else begin
      rob_n_flits_1 <= _GEN_1666;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_2 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_2 <= _GEN_1667;
      end
    end else begin
      rob_n_flits_2 <= _GEN_1667;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_3 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_3 <= _GEN_1668;
      end
    end else begin
      rob_n_flits_3 <= _GEN_1668;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_4 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_4 <= _GEN_1669;
      end
    end else begin
      rob_n_flits_4 <= _GEN_1669;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_5 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_5 <= _GEN_1670;
      end
    end else begin
      rob_n_flits_5 <= _GEN_1670;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_6 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_6 <= _GEN_1671;
      end
    end else begin
      rob_n_flits_6 <= _GEN_1671;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_7 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_7 <= _GEN_1672;
      end
    end else begin
      rob_n_flits_7 <= _GEN_1672;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h8 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_8 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_8 <= _GEN_1673;
      end
    end else begin
      rob_n_flits_8 <= _GEN_1673;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h9 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_9 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_9 <= _GEN_1674;
      end
    end else begin
      rob_n_flits_9 <= _GEN_1674;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'ha == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_10 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_10 <= _GEN_1675;
      end
    end else begin
      rob_n_flits_10 <= _GEN_1675;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hb == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_11 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_11 <= _GEN_1676;
      end
    end else begin
      rob_n_flits_11 <= _GEN_1676;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hc == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_12 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_12 <= _GEN_1677;
      end
    end else begin
      rob_n_flits_12 <= _GEN_1677;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hd == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_13 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_13 <= _GEN_1678;
      end
    end else begin
      rob_n_flits_13 <= _GEN_1678;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'he == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_14 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_14 <= _GEN_1679;
      end
    end else begin
      rob_n_flits_14 <= _GEN_1679;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hf == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_15 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_15 <= _GEN_1680;
      end
    end else begin
      rob_n_flits_15 <= _GEN_1680;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h10 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_16 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_16 <= _GEN_1681;
      end
    end else begin
      rob_n_flits_16 <= _GEN_1681;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h11 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_17 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_17 <= _GEN_1682;
      end
    end else begin
      rob_n_flits_17 <= _GEN_1682;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h12 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_18 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_18 <= _GEN_1683;
      end
    end else begin
      rob_n_flits_18 <= _GEN_1683;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h13 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_19 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_19 <= _GEN_1684;
      end
    end else begin
      rob_n_flits_19 <= _GEN_1684;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h14 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_20 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_20 <= _GEN_1685;
      end
    end else begin
      rob_n_flits_20 <= _GEN_1685;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h15 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_21 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_21 <= _GEN_1686;
      end
    end else begin
      rob_n_flits_21 <= _GEN_1686;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h16 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_22 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_22 <= _GEN_1687;
      end
    end else begin
      rob_n_flits_22 <= _GEN_1687;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h17 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_23 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_23 <= _GEN_1688;
      end
    end else begin
      rob_n_flits_23 <= _GEN_1688;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h18 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_24 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_24 <= _GEN_1689;
      end
    end else begin
      rob_n_flits_24 <= _GEN_1689;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h19 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_25 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_25 <= _GEN_1690;
      end
    end else begin
      rob_n_flits_25 <= _GEN_1690;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1a == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_26 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_26 <= _GEN_1691;
      end
    end else begin
      rob_n_flits_26 <= _GEN_1691;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1b == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_27 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_27 <= _GEN_1692;
      end
    end else begin
      rob_n_flits_27 <= _GEN_1692;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1c == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_28 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_28 <= _GEN_1693;
      end
    end else begin
      rob_n_flits_28 <= _GEN_1693;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1d == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_29 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_29 <= _GEN_1694;
      end
    end else begin
      rob_n_flits_29 <= _GEN_1694;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1e == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_30 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_30 <= _GEN_1695;
      end
    end else begin
      rob_n_flits_30 <= _GEN_1695;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1f == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_31 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_31 <= _GEN_1696;
      end
    end else begin
      rob_n_flits_31 <= _GEN_1696;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h20 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_32 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_32 <= _GEN_1697;
      end
    end else begin
      rob_n_flits_32 <= _GEN_1697;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h21 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_33 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_33 <= _GEN_1698;
      end
    end else begin
      rob_n_flits_33 <= _GEN_1698;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h22 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_34 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_34 <= _GEN_1699;
      end
    end else begin
      rob_n_flits_34 <= _GEN_1699;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h23 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_35 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_35 <= _GEN_1700;
      end
    end else begin
      rob_n_flits_35 <= _GEN_1700;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h24 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_36 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_36 <= _GEN_1701;
      end
    end else begin
      rob_n_flits_36 <= _GEN_1701;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h25 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_37 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_37 <= _GEN_1702;
      end
    end else begin
      rob_n_flits_37 <= _GEN_1702;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h26 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_38 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_38 <= _GEN_1703;
      end
    end else begin
      rob_n_flits_38 <= _GEN_1703;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h27 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_39 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_39 <= _GEN_1704;
      end
    end else begin
      rob_n_flits_39 <= _GEN_1704;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h28 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_40 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_40 <= _GEN_1705;
      end
    end else begin
      rob_n_flits_40 <= _GEN_1705;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h29 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_41 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_41 <= _GEN_1706;
      end
    end else begin
      rob_n_flits_41 <= _GEN_1706;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2a == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_42 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_42 <= _GEN_1707;
      end
    end else begin
      rob_n_flits_42 <= _GEN_1707;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2b == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_43 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_43 <= _GEN_1708;
      end
    end else begin
      rob_n_flits_43 <= _GEN_1708;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2c == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_44 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_44 <= _GEN_1709;
      end
    end else begin
      rob_n_flits_44 <= _GEN_1709;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2d == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_45 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_45 <= _GEN_1710;
      end
    end else begin
      rob_n_flits_45 <= _GEN_1710;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2e == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_46 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_46 <= _GEN_1711;
      end
    end else begin
      rob_n_flits_46 <= _GEN_1711;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2f == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_47 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_47 <= _GEN_1712;
      end
    end else begin
      rob_n_flits_47 <= _GEN_1712;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h30 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_48 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_48 <= _GEN_1713;
      end
    end else begin
      rob_n_flits_48 <= _GEN_1713;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h31 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_49 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_49 <= _GEN_1714;
      end
    end else begin
      rob_n_flits_49 <= _GEN_1714;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h32 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_50 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_50 <= _GEN_1715;
      end
    end else begin
      rob_n_flits_50 <= _GEN_1715;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h33 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_51 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_51 <= _GEN_1716;
      end
    end else begin
      rob_n_flits_51 <= _GEN_1716;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h34 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_52 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_52 <= _GEN_1717;
      end
    end else begin
      rob_n_flits_52 <= _GEN_1717;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h35 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_53 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_53 <= _GEN_1718;
      end
    end else begin
      rob_n_flits_53 <= _GEN_1718;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h36 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_54 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_54 <= _GEN_1719;
      end
    end else begin
      rob_n_flits_54 <= _GEN_1719;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h37 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_55 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_55 <= _GEN_1720;
      end
    end else begin
      rob_n_flits_55 <= _GEN_1720;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h38 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_56 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_56 <= _GEN_1721;
      end
    end else begin
      rob_n_flits_56 <= _GEN_1721;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h39 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_57 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_57 <= _GEN_1722;
      end
    end else begin
      rob_n_flits_57 <= _GEN_1722;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3a == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_58 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_58 <= _GEN_1723;
      end
    end else begin
      rob_n_flits_58 <= _GEN_1723;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3b == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_59 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_59 <= _GEN_1724;
      end
    end else begin
      rob_n_flits_59 <= _GEN_1724;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3c == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_60 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_60 <= _GEN_1725;
      end
    end else begin
      rob_n_flits_60 <= _GEN_1725;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3d == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_61 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_61 <= _GEN_1726;
      end
    end else begin
      rob_n_flits_61 <= _GEN_1726;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3e == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_62 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_62 <= _GEN_1727;
      end
    end else begin
      rob_n_flits_62 <= _GEN_1727;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3f == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_63 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_63 <= _GEN_1728;
      end
    end else begin
      rob_n_flits_63 <= _GEN_1728;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h40 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_64 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_64 <= _GEN_1729;
      end
    end else begin
      rob_n_flits_64 <= _GEN_1729;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h41 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_65 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_65 <= _GEN_1730;
      end
    end else begin
      rob_n_flits_65 <= _GEN_1730;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h42 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_66 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_66 <= _GEN_1731;
      end
    end else begin
      rob_n_flits_66 <= _GEN_1731;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h43 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_67 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_67 <= _GEN_1732;
      end
    end else begin
      rob_n_flits_67 <= _GEN_1732;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h44 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_68 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_68 <= _GEN_1733;
      end
    end else begin
      rob_n_flits_68 <= _GEN_1733;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h45 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_69 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_69 <= _GEN_1734;
      end
    end else begin
      rob_n_flits_69 <= _GEN_1734;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h46 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_70 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_70 <= _GEN_1735;
      end
    end else begin
      rob_n_flits_70 <= _GEN_1735;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h47 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_71 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_71 <= _GEN_1736;
      end
    end else begin
      rob_n_flits_71 <= _GEN_1736;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h48 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_72 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_72 <= _GEN_1737;
      end
    end else begin
      rob_n_flits_72 <= _GEN_1737;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h49 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_73 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_73 <= _GEN_1738;
      end
    end else begin
      rob_n_flits_73 <= _GEN_1738;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4a == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_74 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_74 <= _GEN_1739;
      end
    end else begin
      rob_n_flits_74 <= _GEN_1739;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4b == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_75 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_75 <= _GEN_1740;
      end
    end else begin
      rob_n_flits_75 <= _GEN_1740;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4c == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_76 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_76 <= _GEN_1741;
      end
    end else begin
      rob_n_flits_76 <= _GEN_1741;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4d == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_77 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_77 <= _GEN_1742;
      end
    end else begin
      rob_n_flits_77 <= _GEN_1742;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4e == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_78 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_78 <= _GEN_1743;
      end
    end else begin
      rob_n_flits_78 <= _GEN_1743;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4f == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_79 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_79 <= _GEN_1744;
      end
    end else begin
      rob_n_flits_79 <= _GEN_1744;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h50 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_80 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_80 <= _GEN_1745;
      end
    end else begin
      rob_n_flits_80 <= _GEN_1745;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h51 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_81 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_81 <= _GEN_1746;
      end
    end else begin
      rob_n_flits_81 <= _GEN_1746;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h52 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_82 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_82 <= _GEN_1747;
      end
    end else begin
      rob_n_flits_82 <= _GEN_1747;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h53 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_83 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_83 <= _GEN_1748;
      end
    end else begin
      rob_n_flits_83 <= _GEN_1748;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h54 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_84 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_84 <= _GEN_1749;
      end
    end else begin
      rob_n_flits_84 <= _GEN_1749;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h55 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_85 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_85 <= _GEN_1750;
      end
    end else begin
      rob_n_flits_85 <= _GEN_1750;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h56 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_86 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_86 <= _GEN_1751;
      end
    end else begin
      rob_n_flits_86 <= _GEN_1751;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h57 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_87 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_87 <= _GEN_1752;
      end
    end else begin
      rob_n_flits_87 <= _GEN_1752;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h58 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_88 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_88 <= _GEN_1753;
      end
    end else begin
      rob_n_flits_88 <= _GEN_1753;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h59 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_89 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_89 <= _GEN_1754;
      end
    end else begin
      rob_n_flits_89 <= _GEN_1754;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5a == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_90 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_90 <= _GEN_1755;
      end
    end else begin
      rob_n_flits_90 <= _GEN_1755;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5b == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_91 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_91 <= _GEN_1756;
      end
    end else begin
      rob_n_flits_91 <= _GEN_1756;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5c == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_92 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_92 <= _GEN_1757;
      end
    end else begin
      rob_n_flits_92 <= _GEN_1757;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5d == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_93 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_93 <= _GEN_1758;
      end
    end else begin
      rob_n_flits_93 <= _GEN_1758;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5e == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_94 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_94 <= _GEN_1759;
      end
    end else begin
      rob_n_flits_94 <= _GEN_1759;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5f == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_95 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_95 <= _GEN_1760;
      end
    end else begin
      rob_n_flits_95 <= _GEN_1760;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h60 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_96 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_96 <= _GEN_1761;
      end
    end else begin
      rob_n_flits_96 <= _GEN_1761;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h61 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_97 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_97 <= _GEN_1762;
      end
    end else begin
      rob_n_flits_97 <= _GEN_1762;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h62 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_98 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_98 <= _GEN_1763;
      end
    end else begin
      rob_n_flits_98 <= _GEN_1763;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h63 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_99 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_99 <= _GEN_1764;
      end
    end else begin
      rob_n_flits_99 <= _GEN_1764;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h64 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_100 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_100 <= _GEN_1765;
      end
    end else begin
      rob_n_flits_100 <= _GEN_1765;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h65 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_101 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_101 <= _GEN_1766;
      end
    end else begin
      rob_n_flits_101 <= _GEN_1766;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h66 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_102 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_102 <= _GEN_1767;
      end
    end else begin
      rob_n_flits_102 <= _GEN_1767;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h67 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_103 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_103 <= _GEN_1768;
      end
    end else begin
      rob_n_flits_103 <= _GEN_1768;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h68 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_104 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_104 <= _GEN_1769;
      end
    end else begin
      rob_n_flits_104 <= _GEN_1769;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h69 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_105 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_105 <= _GEN_1770;
      end
    end else begin
      rob_n_flits_105 <= _GEN_1770;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6a == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_106 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_106 <= _GEN_1771;
      end
    end else begin
      rob_n_flits_106 <= _GEN_1771;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6b == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_107 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_107 <= _GEN_1772;
      end
    end else begin
      rob_n_flits_107 <= _GEN_1772;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6c == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_108 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_108 <= _GEN_1773;
      end
    end else begin
      rob_n_flits_108 <= _GEN_1773;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6d == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_109 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_109 <= _GEN_1774;
      end
    end else begin
      rob_n_flits_109 <= _GEN_1774;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6e == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_110 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_110 <= _GEN_1775;
      end
    end else begin
      rob_n_flits_110 <= _GEN_1775;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6f == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_111 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_111 <= _GEN_1776;
      end
    end else begin
      rob_n_flits_111 <= _GEN_1776;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h70 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_112 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_112 <= _GEN_1777;
      end
    end else begin
      rob_n_flits_112 <= _GEN_1777;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h71 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_113 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_113 <= _GEN_1778;
      end
    end else begin
      rob_n_flits_113 <= _GEN_1778;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h72 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_114 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_114 <= _GEN_1779;
      end
    end else begin
      rob_n_flits_114 <= _GEN_1779;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h73 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_115 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_115 <= _GEN_1780;
      end
    end else begin
      rob_n_flits_115 <= _GEN_1780;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h74 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_116 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_116 <= _GEN_1781;
      end
    end else begin
      rob_n_flits_116 <= _GEN_1781;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h75 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_117 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_117 <= _GEN_1782;
      end
    end else begin
      rob_n_flits_117 <= _GEN_1782;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h76 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_118 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_118 <= _GEN_1783;
      end
    end else begin
      rob_n_flits_118 <= _GEN_1783;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h77 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_119 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_119 <= _GEN_1784;
      end
    end else begin
      rob_n_flits_119 <= _GEN_1784;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h78 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_120 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_120 <= _GEN_1785;
      end
    end else begin
      rob_n_flits_120 <= _GEN_1785;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h79 == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_121 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_121 <= _GEN_1786;
      end
    end else begin
      rob_n_flits_121 <= _GEN_1786;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7a == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_122 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_122 <= _GEN_1787;
      end
    end else begin
      rob_n_flits_122 <= _GEN_1787;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7b == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_123 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_123 <= _GEN_1788;
      end
    end else begin
      rob_n_flits_123 <= _GEN_1788;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7c == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_124 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_124 <= _GEN_1789;
      end
    end else begin
      rob_n_flits_124 <= _GEN_1789;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7d == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_125 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_125 <= _GEN_1790;
      end
    end else begin
      rob_n_flits_125 <= _GEN_1790;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7e == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_126 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_126 <= _GEN_1791;
      end
    end else begin
      rob_n_flits_126 <= _GEN_1791;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7f == rob_alloc_ids_1) begin // @[TestHarness.scala 182:36]
        rob_n_flits_127 <= _rob_n_flits_T_35; // @[TestHarness.scala 182:36]
      end else begin
        rob_n_flits_127 <= _GEN_1792;
      end
    end else begin
      rob_n_flits_127 <= _GEN_1792;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h0 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_0 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_0 <= _GEN_5636;
      end
    end else begin
      rob_flits_returned_0 <= _GEN_5636;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h1 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_1 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_1 <= _GEN_5637;
      end
    end else begin
      rob_flits_returned_1 <= _GEN_5637;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h2 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_2 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_2 <= _GEN_5638;
      end
    end else begin
      rob_flits_returned_2 <= _GEN_5638;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h3 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_3 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_3 <= _GEN_5639;
      end
    end else begin
      rob_flits_returned_3 <= _GEN_5639;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h4 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_4 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_4 <= _GEN_5640;
      end
    end else begin
      rob_flits_returned_4 <= _GEN_5640;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h5 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_5 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_5 <= _GEN_5641;
      end
    end else begin
      rob_flits_returned_5 <= _GEN_5641;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h6 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_6 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_6 <= _GEN_5642;
      end
    end else begin
      rob_flits_returned_6 <= _GEN_5642;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h7 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_7 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_7 <= _GEN_5643;
      end
    end else begin
      rob_flits_returned_7 <= _GEN_5643;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h8 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_8 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_8 <= _GEN_5644;
      end
    end else begin
      rob_flits_returned_8 <= _GEN_5644;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h9 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_9 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_9 <= _GEN_5645;
      end
    end else begin
      rob_flits_returned_9 <= _GEN_5645;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'ha == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_10 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_10 <= _GEN_5646;
      end
    end else begin
      rob_flits_returned_10 <= _GEN_5646;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'hb == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_11 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_11 <= _GEN_5647;
      end
    end else begin
      rob_flits_returned_11 <= _GEN_5647;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'hc == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_12 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_12 <= _GEN_5648;
      end
    end else begin
      rob_flits_returned_12 <= _GEN_5648;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'hd == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_13 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_13 <= _GEN_5649;
      end
    end else begin
      rob_flits_returned_13 <= _GEN_5649;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'he == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_14 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_14 <= _GEN_5650;
      end
    end else begin
      rob_flits_returned_14 <= _GEN_5650;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'hf == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_15 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_15 <= _GEN_5651;
      end
    end else begin
      rob_flits_returned_15 <= _GEN_5651;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h10 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_16 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_16 <= _GEN_5652;
      end
    end else begin
      rob_flits_returned_16 <= _GEN_5652;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h11 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_17 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_17 <= _GEN_5653;
      end
    end else begin
      rob_flits_returned_17 <= _GEN_5653;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h12 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_18 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_18 <= _GEN_5654;
      end
    end else begin
      rob_flits_returned_18 <= _GEN_5654;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h13 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_19 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_19 <= _GEN_5655;
      end
    end else begin
      rob_flits_returned_19 <= _GEN_5655;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h14 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_20 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_20 <= _GEN_5656;
      end
    end else begin
      rob_flits_returned_20 <= _GEN_5656;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h15 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_21 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_21 <= _GEN_5657;
      end
    end else begin
      rob_flits_returned_21 <= _GEN_5657;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h16 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_22 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_22 <= _GEN_5658;
      end
    end else begin
      rob_flits_returned_22 <= _GEN_5658;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h17 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_23 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_23 <= _GEN_5659;
      end
    end else begin
      rob_flits_returned_23 <= _GEN_5659;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h18 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_24 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_24 <= _GEN_5660;
      end
    end else begin
      rob_flits_returned_24 <= _GEN_5660;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h19 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_25 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_25 <= _GEN_5661;
      end
    end else begin
      rob_flits_returned_25 <= _GEN_5661;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h1a == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_26 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_26 <= _GEN_5662;
      end
    end else begin
      rob_flits_returned_26 <= _GEN_5662;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h1b == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_27 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_27 <= _GEN_5663;
      end
    end else begin
      rob_flits_returned_27 <= _GEN_5663;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h1c == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_28 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_28 <= _GEN_5664;
      end
    end else begin
      rob_flits_returned_28 <= _GEN_5664;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h1d == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_29 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_29 <= _GEN_5665;
      end
    end else begin
      rob_flits_returned_29 <= _GEN_5665;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h1e == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_30 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_30 <= _GEN_5666;
      end
    end else begin
      rob_flits_returned_30 <= _GEN_5666;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h1f == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_31 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_31 <= _GEN_5667;
      end
    end else begin
      rob_flits_returned_31 <= _GEN_5667;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h20 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_32 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_32 <= _GEN_5668;
      end
    end else begin
      rob_flits_returned_32 <= _GEN_5668;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h21 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_33 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_33 <= _GEN_5669;
      end
    end else begin
      rob_flits_returned_33 <= _GEN_5669;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h22 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_34 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_34 <= _GEN_5670;
      end
    end else begin
      rob_flits_returned_34 <= _GEN_5670;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h23 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_35 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_35 <= _GEN_5671;
      end
    end else begin
      rob_flits_returned_35 <= _GEN_5671;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h24 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_36 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_36 <= _GEN_5672;
      end
    end else begin
      rob_flits_returned_36 <= _GEN_5672;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h25 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_37 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_37 <= _GEN_5673;
      end
    end else begin
      rob_flits_returned_37 <= _GEN_5673;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h26 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_38 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_38 <= _GEN_5674;
      end
    end else begin
      rob_flits_returned_38 <= _GEN_5674;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h27 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_39 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_39 <= _GEN_5675;
      end
    end else begin
      rob_flits_returned_39 <= _GEN_5675;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h28 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_40 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_40 <= _GEN_5676;
      end
    end else begin
      rob_flits_returned_40 <= _GEN_5676;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h29 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_41 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_41 <= _GEN_5677;
      end
    end else begin
      rob_flits_returned_41 <= _GEN_5677;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h2a == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_42 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_42 <= _GEN_5678;
      end
    end else begin
      rob_flits_returned_42 <= _GEN_5678;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h2b == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_43 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_43 <= _GEN_5679;
      end
    end else begin
      rob_flits_returned_43 <= _GEN_5679;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h2c == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_44 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_44 <= _GEN_5680;
      end
    end else begin
      rob_flits_returned_44 <= _GEN_5680;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h2d == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_45 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_45 <= _GEN_5681;
      end
    end else begin
      rob_flits_returned_45 <= _GEN_5681;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h2e == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_46 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_46 <= _GEN_5682;
      end
    end else begin
      rob_flits_returned_46 <= _GEN_5682;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h2f == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_47 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_47 <= _GEN_5683;
      end
    end else begin
      rob_flits_returned_47 <= _GEN_5683;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h30 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_48 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_48 <= _GEN_5684;
      end
    end else begin
      rob_flits_returned_48 <= _GEN_5684;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h31 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_49 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_49 <= _GEN_5685;
      end
    end else begin
      rob_flits_returned_49 <= _GEN_5685;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h32 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_50 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_50 <= _GEN_5686;
      end
    end else begin
      rob_flits_returned_50 <= _GEN_5686;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h33 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_51 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_51 <= _GEN_5687;
      end
    end else begin
      rob_flits_returned_51 <= _GEN_5687;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h34 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_52 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_52 <= _GEN_5688;
      end
    end else begin
      rob_flits_returned_52 <= _GEN_5688;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h35 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_53 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_53 <= _GEN_5689;
      end
    end else begin
      rob_flits_returned_53 <= _GEN_5689;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h36 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_54 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_54 <= _GEN_5690;
      end
    end else begin
      rob_flits_returned_54 <= _GEN_5690;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h37 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_55 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_55 <= _GEN_5691;
      end
    end else begin
      rob_flits_returned_55 <= _GEN_5691;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h38 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_56 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_56 <= _GEN_5692;
      end
    end else begin
      rob_flits_returned_56 <= _GEN_5692;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h39 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_57 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_57 <= _GEN_5693;
      end
    end else begin
      rob_flits_returned_57 <= _GEN_5693;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h3a == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_58 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_58 <= _GEN_5694;
      end
    end else begin
      rob_flits_returned_58 <= _GEN_5694;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h3b == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_59 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_59 <= _GEN_5695;
      end
    end else begin
      rob_flits_returned_59 <= _GEN_5695;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h3c == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_60 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_60 <= _GEN_5696;
      end
    end else begin
      rob_flits_returned_60 <= _GEN_5696;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h3d == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_61 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_61 <= _GEN_5697;
      end
    end else begin
      rob_flits_returned_61 <= _GEN_5697;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h3e == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_62 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_62 <= _GEN_5698;
      end
    end else begin
      rob_flits_returned_62 <= _GEN_5698;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h3f == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_63 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_63 <= _GEN_5699;
      end
    end else begin
      rob_flits_returned_63 <= _GEN_5699;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h40 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_64 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_64 <= _GEN_5700;
      end
    end else begin
      rob_flits_returned_64 <= _GEN_5700;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h41 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_65 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_65 <= _GEN_5701;
      end
    end else begin
      rob_flits_returned_65 <= _GEN_5701;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h42 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_66 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_66 <= _GEN_5702;
      end
    end else begin
      rob_flits_returned_66 <= _GEN_5702;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h43 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_67 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_67 <= _GEN_5703;
      end
    end else begin
      rob_flits_returned_67 <= _GEN_5703;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h44 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_68 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_68 <= _GEN_5704;
      end
    end else begin
      rob_flits_returned_68 <= _GEN_5704;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h45 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_69 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_69 <= _GEN_5705;
      end
    end else begin
      rob_flits_returned_69 <= _GEN_5705;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h46 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_70 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_70 <= _GEN_5706;
      end
    end else begin
      rob_flits_returned_70 <= _GEN_5706;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h47 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_71 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_71 <= _GEN_5707;
      end
    end else begin
      rob_flits_returned_71 <= _GEN_5707;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h48 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_72 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_72 <= _GEN_5708;
      end
    end else begin
      rob_flits_returned_72 <= _GEN_5708;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h49 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_73 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_73 <= _GEN_5709;
      end
    end else begin
      rob_flits_returned_73 <= _GEN_5709;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h4a == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_74 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_74 <= _GEN_5710;
      end
    end else begin
      rob_flits_returned_74 <= _GEN_5710;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h4b == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_75 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_75 <= _GEN_5711;
      end
    end else begin
      rob_flits_returned_75 <= _GEN_5711;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h4c == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_76 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_76 <= _GEN_5712;
      end
    end else begin
      rob_flits_returned_76 <= _GEN_5712;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h4d == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_77 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_77 <= _GEN_5713;
      end
    end else begin
      rob_flits_returned_77 <= _GEN_5713;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h4e == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_78 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_78 <= _GEN_5714;
      end
    end else begin
      rob_flits_returned_78 <= _GEN_5714;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h4f == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_79 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_79 <= _GEN_5715;
      end
    end else begin
      rob_flits_returned_79 <= _GEN_5715;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h50 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_80 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_80 <= _GEN_5716;
      end
    end else begin
      rob_flits_returned_80 <= _GEN_5716;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h51 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_81 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_81 <= _GEN_5717;
      end
    end else begin
      rob_flits_returned_81 <= _GEN_5717;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h52 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_82 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_82 <= _GEN_5718;
      end
    end else begin
      rob_flits_returned_82 <= _GEN_5718;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h53 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_83 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_83 <= _GEN_5719;
      end
    end else begin
      rob_flits_returned_83 <= _GEN_5719;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h54 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_84 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_84 <= _GEN_5720;
      end
    end else begin
      rob_flits_returned_84 <= _GEN_5720;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h55 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_85 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_85 <= _GEN_5721;
      end
    end else begin
      rob_flits_returned_85 <= _GEN_5721;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h56 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_86 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_86 <= _GEN_5722;
      end
    end else begin
      rob_flits_returned_86 <= _GEN_5722;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h57 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_87 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_87 <= _GEN_5723;
      end
    end else begin
      rob_flits_returned_87 <= _GEN_5723;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h58 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_88 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_88 <= _GEN_5724;
      end
    end else begin
      rob_flits_returned_88 <= _GEN_5724;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h59 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_89 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_89 <= _GEN_5725;
      end
    end else begin
      rob_flits_returned_89 <= _GEN_5725;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h5a == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_90 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_90 <= _GEN_5726;
      end
    end else begin
      rob_flits_returned_90 <= _GEN_5726;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h5b == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_91 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_91 <= _GEN_5727;
      end
    end else begin
      rob_flits_returned_91 <= _GEN_5727;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h5c == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_92 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_92 <= _GEN_5728;
      end
    end else begin
      rob_flits_returned_92 <= _GEN_5728;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h5d == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_93 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_93 <= _GEN_5729;
      end
    end else begin
      rob_flits_returned_93 <= _GEN_5729;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h5e == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_94 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_94 <= _GEN_5730;
      end
    end else begin
      rob_flits_returned_94 <= _GEN_5730;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h5f == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_95 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_95 <= _GEN_5731;
      end
    end else begin
      rob_flits_returned_95 <= _GEN_5731;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h60 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_96 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_96 <= _GEN_5732;
      end
    end else begin
      rob_flits_returned_96 <= _GEN_5732;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h61 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_97 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_97 <= _GEN_5733;
      end
    end else begin
      rob_flits_returned_97 <= _GEN_5733;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h62 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_98 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_98 <= _GEN_5734;
      end
    end else begin
      rob_flits_returned_98 <= _GEN_5734;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h63 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_99 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_99 <= _GEN_5735;
      end
    end else begin
      rob_flits_returned_99 <= _GEN_5735;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h64 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_100 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_100 <= _GEN_5736;
      end
    end else begin
      rob_flits_returned_100 <= _GEN_5736;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h65 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_101 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_101 <= _GEN_5737;
      end
    end else begin
      rob_flits_returned_101 <= _GEN_5737;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h66 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_102 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_102 <= _GEN_5738;
      end
    end else begin
      rob_flits_returned_102 <= _GEN_5738;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h67 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_103 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_103 <= _GEN_5739;
      end
    end else begin
      rob_flits_returned_103 <= _GEN_5739;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h68 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_104 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_104 <= _GEN_5740;
      end
    end else begin
      rob_flits_returned_104 <= _GEN_5740;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h69 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_105 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_105 <= _GEN_5741;
      end
    end else begin
      rob_flits_returned_105 <= _GEN_5741;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h6a == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_106 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_106 <= _GEN_5742;
      end
    end else begin
      rob_flits_returned_106 <= _GEN_5742;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h6b == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_107 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_107 <= _GEN_5743;
      end
    end else begin
      rob_flits_returned_107 <= _GEN_5743;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h6c == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_108 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_108 <= _GEN_5744;
      end
    end else begin
      rob_flits_returned_108 <= _GEN_5744;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h6d == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_109 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_109 <= _GEN_5745;
      end
    end else begin
      rob_flits_returned_109 <= _GEN_5745;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h6e == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_110 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_110 <= _GEN_5746;
      end
    end else begin
      rob_flits_returned_110 <= _GEN_5746;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h6f == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_111 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_111 <= _GEN_5747;
      end
    end else begin
      rob_flits_returned_111 <= _GEN_5747;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h70 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_112 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_112 <= _GEN_5748;
      end
    end else begin
      rob_flits_returned_112 <= _GEN_5748;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h71 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_113 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_113 <= _GEN_5749;
      end
    end else begin
      rob_flits_returned_113 <= _GEN_5749;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h72 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_114 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_114 <= _GEN_5750;
      end
    end else begin
      rob_flits_returned_114 <= _GEN_5750;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h73 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_115 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_115 <= _GEN_5751;
      end
    end else begin
      rob_flits_returned_115 <= _GEN_5751;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h74 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_116 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_116 <= _GEN_5752;
      end
    end else begin
      rob_flits_returned_116 <= _GEN_5752;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h75 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_117 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_117 <= _GEN_5753;
      end
    end else begin
      rob_flits_returned_117 <= _GEN_5753;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h76 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_118 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_118 <= _GEN_5754;
      end
    end else begin
      rob_flits_returned_118 <= _GEN_5754;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h77 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_119 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_119 <= _GEN_5755;
      end
    end else begin
      rob_flits_returned_119 <= _GEN_5755;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h78 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_120 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_120 <= _GEN_5756;
      end
    end else begin
      rob_flits_returned_120 <= _GEN_5756;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h79 == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_121 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_121 <= _GEN_5757;
      end
    end else begin
      rob_flits_returned_121 <= _GEN_5757;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h7a == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_122 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_122 <= _GEN_5758;
      end
    end else begin
      rob_flits_returned_122 <= _GEN_5758;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h7b == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_123 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_123 <= _GEN_5759;
      end
    end else begin
      rob_flits_returned_123 <= _GEN_5759;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h7c == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_124 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_124 <= _GEN_5760;
      end
    end else begin
      rob_flits_returned_124 <= _GEN_5760;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h7d == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_125 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_125 <= _GEN_5761;
      end
    end else begin
      rob_flits_returned_125 <= _GEN_5761;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h7e == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_126 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_126 <= _GEN_5762;
      end
    end else begin
      rob_flits_returned_126 <= _GEN_5762;
    end
    if (_T_131) begin // @[TestHarness.scala 199:26]
      if (7'h7f == out_payload_1_rob_idx[6:0]) begin // @[TestHarness.scala 213:35]
        rob_flits_returned_127 <= _rob_flits_returned_T_5; // @[TestHarness.scala 213:35]
      end else begin
        rob_flits_returned_127 <= _GEN_5763;
      end
    end else begin
      rob_flits_returned_127 <= _GEN_5763;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h0 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_0 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_0 <= _GEN_1921;
      end
    end else begin
      rob_tscs_0 <= _GEN_1921;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_1 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_1 <= _GEN_1922;
      end
    end else begin
      rob_tscs_1 <= _GEN_1922;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_2 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_2 <= _GEN_1923;
      end
    end else begin
      rob_tscs_2 <= _GEN_1923;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_3 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_3 <= _GEN_1924;
      end
    end else begin
      rob_tscs_3 <= _GEN_1924;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_4 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_4 <= _GEN_1925;
      end
    end else begin
      rob_tscs_4 <= _GEN_1925;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_5 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_5 <= _GEN_1926;
      end
    end else begin
      rob_tscs_5 <= _GEN_1926;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_6 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_6 <= _GEN_1927;
      end
    end else begin
      rob_tscs_6 <= _GEN_1927;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_7 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_7 <= _GEN_1928;
      end
    end else begin
      rob_tscs_7 <= _GEN_1928;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h8 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_8 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_8 <= _GEN_1929;
      end
    end else begin
      rob_tscs_8 <= _GEN_1929;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h9 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_9 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_9 <= _GEN_1930;
      end
    end else begin
      rob_tscs_9 <= _GEN_1930;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'ha == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_10 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_10 <= _GEN_1931;
      end
    end else begin
      rob_tscs_10 <= _GEN_1931;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hb == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_11 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_11 <= _GEN_1932;
      end
    end else begin
      rob_tscs_11 <= _GEN_1932;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hc == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_12 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_12 <= _GEN_1933;
      end
    end else begin
      rob_tscs_12 <= _GEN_1933;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hd == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_13 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_13 <= _GEN_1934;
      end
    end else begin
      rob_tscs_13 <= _GEN_1934;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'he == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_14 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_14 <= _GEN_1935;
      end
    end else begin
      rob_tscs_14 <= _GEN_1935;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'hf == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_15 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_15 <= _GEN_1936;
      end
    end else begin
      rob_tscs_15 <= _GEN_1936;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h10 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_16 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_16 <= _GEN_1937;
      end
    end else begin
      rob_tscs_16 <= _GEN_1937;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h11 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_17 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_17 <= _GEN_1938;
      end
    end else begin
      rob_tscs_17 <= _GEN_1938;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h12 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_18 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_18 <= _GEN_1939;
      end
    end else begin
      rob_tscs_18 <= _GEN_1939;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h13 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_19 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_19 <= _GEN_1940;
      end
    end else begin
      rob_tscs_19 <= _GEN_1940;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h14 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_20 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_20 <= _GEN_1941;
      end
    end else begin
      rob_tscs_20 <= _GEN_1941;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h15 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_21 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_21 <= _GEN_1942;
      end
    end else begin
      rob_tscs_21 <= _GEN_1942;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h16 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_22 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_22 <= _GEN_1943;
      end
    end else begin
      rob_tscs_22 <= _GEN_1943;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h17 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_23 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_23 <= _GEN_1944;
      end
    end else begin
      rob_tscs_23 <= _GEN_1944;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h18 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_24 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_24 <= _GEN_1945;
      end
    end else begin
      rob_tscs_24 <= _GEN_1945;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h19 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_25 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_25 <= _GEN_1946;
      end
    end else begin
      rob_tscs_25 <= _GEN_1946;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1a == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_26 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_26 <= _GEN_1947;
      end
    end else begin
      rob_tscs_26 <= _GEN_1947;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1b == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_27 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_27 <= _GEN_1948;
      end
    end else begin
      rob_tscs_27 <= _GEN_1948;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1c == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_28 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_28 <= _GEN_1949;
      end
    end else begin
      rob_tscs_28 <= _GEN_1949;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1d == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_29 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_29 <= _GEN_1950;
      end
    end else begin
      rob_tscs_29 <= _GEN_1950;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1e == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_30 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_30 <= _GEN_1951;
      end
    end else begin
      rob_tscs_30 <= _GEN_1951;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h1f == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_31 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_31 <= _GEN_1952;
      end
    end else begin
      rob_tscs_31 <= _GEN_1952;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h20 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_32 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_32 <= _GEN_1953;
      end
    end else begin
      rob_tscs_32 <= _GEN_1953;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h21 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_33 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_33 <= _GEN_1954;
      end
    end else begin
      rob_tscs_33 <= _GEN_1954;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h22 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_34 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_34 <= _GEN_1955;
      end
    end else begin
      rob_tscs_34 <= _GEN_1955;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h23 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_35 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_35 <= _GEN_1956;
      end
    end else begin
      rob_tscs_35 <= _GEN_1956;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h24 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_36 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_36 <= _GEN_1957;
      end
    end else begin
      rob_tscs_36 <= _GEN_1957;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h25 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_37 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_37 <= _GEN_1958;
      end
    end else begin
      rob_tscs_37 <= _GEN_1958;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h26 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_38 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_38 <= _GEN_1959;
      end
    end else begin
      rob_tscs_38 <= _GEN_1959;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h27 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_39 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_39 <= _GEN_1960;
      end
    end else begin
      rob_tscs_39 <= _GEN_1960;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h28 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_40 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_40 <= _GEN_1961;
      end
    end else begin
      rob_tscs_40 <= _GEN_1961;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h29 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_41 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_41 <= _GEN_1962;
      end
    end else begin
      rob_tscs_41 <= _GEN_1962;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2a == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_42 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_42 <= _GEN_1963;
      end
    end else begin
      rob_tscs_42 <= _GEN_1963;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2b == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_43 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_43 <= _GEN_1964;
      end
    end else begin
      rob_tscs_43 <= _GEN_1964;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2c == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_44 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_44 <= _GEN_1965;
      end
    end else begin
      rob_tscs_44 <= _GEN_1965;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2d == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_45 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_45 <= _GEN_1966;
      end
    end else begin
      rob_tscs_45 <= _GEN_1966;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2e == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_46 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_46 <= _GEN_1967;
      end
    end else begin
      rob_tscs_46 <= _GEN_1967;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h2f == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_47 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_47 <= _GEN_1968;
      end
    end else begin
      rob_tscs_47 <= _GEN_1968;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h30 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_48 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_48 <= _GEN_1969;
      end
    end else begin
      rob_tscs_48 <= _GEN_1969;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h31 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_49 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_49 <= _GEN_1970;
      end
    end else begin
      rob_tscs_49 <= _GEN_1970;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h32 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_50 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_50 <= _GEN_1971;
      end
    end else begin
      rob_tscs_50 <= _GEN_1971;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h33 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_51 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_51 <= _GEN_1972;
      end
    end else begin
      rob_tscs_51 <= _GEN_1972;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h34 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_52 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_52 <= _GEN_1973;
      end
    end else begin
      rob_tscs_52 <= _GEN_1973;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h35 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_53 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_53 <= _GEN_1974;
      end
    end else begin
      rob_tscs_53 <= _GEN_1974;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h36 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_54 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_54 <= _GEN_1975;
      end
    end else begin
      rob_tscs_54 <= _GEN_1975;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h37 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_55 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_55 <= _GEN_1976;
      end
    end else begin
      rob_tscs_55 <= _GEN_1976;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h38 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_56 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_56 <= _GEN_1977;
      end
    end else begin
      rob_tscs_56 <= _GEN_1977;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h39 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_57 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_57 <= _GEN_1978;
      end
    end else begin
      rob_tscs_57 <= _GEN_1978;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3a == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_58 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_58 <= _GEN_1979;
      end
    end else begin
      rob_tscs_58 <= _GEN_1979;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3b == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_59 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_59 <= _GEN_1980;
      end
    end else begin
      rob_tscs_59 <= _GEN_1980;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3c == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_60 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_60 <= _GEN_1981;
      end
    end else begin
      rob_tscs_60 <= _GEN_1981;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3d == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_61 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_61 <= _GEN_1982;
      end
    end else begin
      rob_tscs_61 <= _GEN_1982;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3e == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_62 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_62 <= _GEN_1983;
      end
    end else begin
      rob_tscs_62 <= _GEN_1983;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h3f == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_63 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_63 <= _GEN_1984;
      end
    end else begin
      rob_tscs_63 <= _GEN_1984;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h40 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_64 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_64 <= _GEN_1985;
      end
    end else begin
      rob_tscs_64 <= _GEN_1985;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h41 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_65 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_65 <= _GEN_1986;
      end
    end else begin
      rob_tscs_65 <= _GEN_1986;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h42 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_66 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_66 <= _GEN_1987;
      end
    end else begin
      rob_tscs_66 <= _GEN_1987;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h43 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_67 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_67 <= _GEN_1988;
      end
    end else begin
      rob_tscs_67 <= _GEN_1988;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h44 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_68 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_68 <= _GEN_1989;
      end
    end else begin
      rob_tscs_68 <= _GEN_1989;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h45 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_69 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_69 <= _GEN_1990;
      end
    end else begin
      rob_tscs_69 <= _GEN_1990;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h46 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_70 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_70 <= _GEN_1991;
      end
    end else begin
      rob_tscs_70 <= _GEN_1991;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h47 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_71 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_71 <= _GEN_1992;
      end
    end else begin
      rob_tscs_71 <= _GEN_1992;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h48 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_72 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_72 <= _GEN_1993;
      end
    end else begin
      rob_tscs_72 <= _GEN_1993;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h49 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_73 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_73 <= _GEN_1994;
      end
    end else begin
      rob_tscs_73 <= _GEN_1994;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4a == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_74 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_74 <= _GEN_1995;
      end
    end else begin
      rob_tscs_74 <= _GEN_1995;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4b == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_75 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_75 <= _GEN_1996;
      end
    end else begin
      rob_tscs_75 <= _GEN_1996;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4c == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_76 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_76 <= _GEN_1997;
      end
    end else begin
      rob_tscs_76 <= _GEN_1997;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4d == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_77 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_77 <= _GEN_1998;
      end
    end else begin
      rob_tscs_77 <= _GEN_1998;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4e == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_78 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_78 <= _GEN_1999;
      end
    end else begin
      rob_tscs_78 <= _GEN_1999;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h4f == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_79 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_79 <= _GEN_2000;
      end
    end else begin
      rob_tscs_79 <= _GEN_2000;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h50 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_80 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_80 <= _GEN_2001;
      end
    end else begin
      rob_tscs_80 <= _GEN_2001;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h51 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_81 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_81 <= _GEN_2002;
      end
    end else begin
      rob_tscs_81 <= _GEN_2002;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h52 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_82 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_82 <= _GEN_2003;
      end
    end else begin
      rob_tscs_82 <= _GEN_2003;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h53 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_83 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_83 <= _GEN_2004;
      end
    end else begin
      rob_tscs_83 <= _GEN_2004;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h54 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_84 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_84 <= _GEN_2005;
      end
    end else begin
      rob_tscs_84 <= _GEN_2005;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h55 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_85 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_85 <= _GEN_2006;
      end
    end else begin
      rob_tscs_85 <= _GEN_2006;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h56 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_86 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_86 <= _GEN_2007;
      end
    end else begin
      rob_tscs_86 <= _GEN_2007;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h57 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_87 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_87 <= _GEN_2008;
      end
    end else begin
      rob_tscs_87 <= _GEN_2008;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h58 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_88 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_88 <= _GEN_2009;
      end
    end else begin
      rob_tscs_88 <= _GEN_2009;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h59 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_89 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_89 <= _GEN_2010;
      end
    end else begin
      rob_tscs_89 <= _GEN_2010;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5a == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_90 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_90 <= _GEN_2011;
      end
    end else begin
      rob_tscs_90 <= _GEN_2011;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5b == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_91 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_91 <= _GEN_2012;
      end
    end else begin
      rob_tscs_91 <= _GEN_2012;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5c == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_92 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_92 <= _GEN_2013;
      end
    end else begin
      rob_tscs_92 <= _GEN_2013;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5d == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_93 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_93 <= _GEN_2014;
      end
    end else begin
      rob_tscs_93 <= _GEN_2014;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5e == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_94 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_94 <= _GEN_2015;
      end
    end else begin
      rob_tscs_94 <= _GEN_2015;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h5f == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_95 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_95 <= _GEN_2016;
      end
    end else begin
      rob_tscs_95 <= _GEN_2016;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h60 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_96 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_96 <= _GEN_2017;
      end
    end else begin
      rob_tscs_96 <= _GEN_2017;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h61 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_97 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_97 <= _GEN_2018;
      end
    end else begin
      rob_tscs_97 <= _GEN_2018;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h62 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_98 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_98 <= _GEN_2019;
      end
    end else begin
      rob_tscs_98 <= _GEN_2019;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h63 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_99 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_99 <= _GEN_2020;
      end
    end else begin
      rob_tscs_99 <= _GEN_2020;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h64 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_100 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_100 <= _GEN_2021;
      end
    end else begin
      rob_tscs_100 <= _GEN_2021;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h65 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_101 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_101 <= _GEN_2022;
      end
    end else begin
      rob_tscs_101 <= _GEN_2022;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h66 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_102 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_102 <= _GEN_2023;
      end
    end else begin
      rob_tscs_102 <= _GEN_2023;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h67 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_103 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_103 <= _GEN_2024;
      end
    end else begin
      rob_tscs_103 <= _GEN_2024;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h68 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_104 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_104 <= _GEN_2025;
      end
    end else begin
      rob_tscs_104 <= _GEN_2025;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h69 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_105 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_105 <= _GEN_2026;
      end
    end else begin
      rob_tscs_105 <= _GEN_2026;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6a == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_106 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_106 <= _GEN_2027;
      end
    end else begin
      rob_tscs_106 <= _GEN_2027;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6b == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_107 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_107 <= _GEN_2028;
      end
    end else begin
      rob_tscs_107 <= _GEN_2028;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6c == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_108 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_108 <= _GEN_2029;
      end
    end else begin
      rob_tscs_108 <= _GEN_2029;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6d == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_109 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_109 <= _GEN_2030;
      end
    end else begin
      rob_tscs_109 <= _GEN_2030;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6e == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_110 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_110 <= _GEN_2031;
      end
    end else begin
      rob_tscs_110 <= _GEN_2031;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h6f == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_111 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_111 <= _GEN_2032;
      end
    end else begin
      rob_tscs_111 <= _GEN_2032;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h70 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_112 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_112 <= _GEN_2033;
      end
    end else begin
      rob_tscs_112 <= _GEN_2033;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h71 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_113 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_113 <= _GEN_2034;
      end
    end else begin
      rob_tscs_113 <= _GEN_2034;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h72 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_114 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_114 <= _GEN_2035;
      end
    end else begin
      rob_tscs_114 <= _GEN_2035;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h73 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_115 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_115 <= _GEN_2036;
      end
    end else begin
      rob_tscs_115 <= _GEN_2036;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h74 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_116 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_116 <= _GEN_2037;
      end
    end else begin
      rob_tscs_116 <= _GEN_2037;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h75 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_117 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_117 <= _GEN_2038;
      end
    end else begin
      rob_tscs_117 <= _GEN_2038;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h76 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_118 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_118 <= _GEN_2039;
      end
    end else begin
      rob_tscs_118 <= _GEN_2039;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h77 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_119 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_119 <= _GEN_2040;
      end
    end else begin
      rob_tscs_119 <= _GEN_2040;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h78 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_120 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_120 <= _GEN_2041;
      end
    end else begin
      rob_tscs_120 <= _GEN_2041;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h79 == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_121 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_121 <= _GEN_2042;
      end
    end else begin
      rob_tscs_121 <= _GEN_2042;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7a == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_122 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_122 <= _GEN_2043;
      end
    end else begin
      rob_tscs_122 <= _GEN_2043;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7b == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_123 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_123 <= _GEN_2044;
      end
    end else begin
      rob_tscs_123 <= _GEN_2044;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7c == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_124 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_124 <= _GEN_2045;
      end
    end else begin
      rob_tscs_124 <= _GEN_2045;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7d == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_125 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_125 <= _GEN_2046;
      end
    end else begin
      rob_tscs_125 <= _GEN_2046;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7e == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_126 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_126 <= _GEN_2047;
      end
    end else begin
      rob_tscs_126 <= _GEN_2047;
    end
    if (igen_1_io_fire) begin // @[TestHarness.scala 178:25]
      if (7'h7f == rob_alloc_ids_1) begin // @[TestHarness.scala 184:36]
        rob_tscs_127 <= _rob_tscs_T_25; // @[TestHarness.scala 184:36]
      end else begin
        rob_tscs_127 <= _GEN_2048;
      end
    end else begin
      rob_tscs_127 <= _GEN_2048;
    end
    if (reset) begin // @[TestHarness.scala 164:24]
      io_success_REG <= 1'h0; // @[TestHarness.scala 164:24]
    end else begin
      io_success_REG <= success; // @[TestHarness.scala 164:24]
    end
    if (reset) begin // @[TestHarness.scala 196:31]
      packet_valid <= 1'h0; // @[TestHarness.scala 196:31]
    end else if (_T_84) begin // @[TestHarness.scala 199:26]
      if (io_from_noc_0_flit_bits_tail) begin // @[TestHarness.scala 216:31]
        packet_valid <= 1'h0; // @[TestHarness.scala 216:46]
      end else begin
        packet_valid <= _GEN_5633;
      end
    end
    packet_rob_idx <= _GEN_5893[6:0];
    if (reset) begin // @[TestHarness.scala 196:31]
      packet_valid_1 <= 1'h0; // @[TestHarness.scala 196:31]
    end else if (_T_131) begin // @[TestHarness.scala 199:26]
      if (io_from_noc_1_flit_bits_tail) begin // @[TestHarness.scala 216:31]
        packet_valid_1 <= 1'h0; // @[TestHarness.scala 216:46]
      end else begin
        packet_valid_1 <= _GEN_7430;
      end
    end
    packet_rob_idx_1 <= _GEN_7690[6:0];
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~idle_counter[10])) begin
          $fwrite(32'h80000002,"Assertion failed\n    at TestHarness.scala:148 assert(!idle_counter(10))\n"); // @[TestHarness.scala 148:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (success & _T_3) begin
          $fwrite(32'h80000002,"%d flits, %d cycles\n",flits,tsc); // @[TestHarness.scala 166:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_84 & _T_3 & ~_T_42[0]) begin
          $fwrite(32'h80000002,
            "Assertion failed: out[0] unexpected response\n    at TestHarness.scala:201 assert(rob_valids(rob_idx), cf\"out[${i.toString}] unexpected response\")\n"
            ); // @[TestHarness.scala 201:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_7953 & ~(_T_48 == io_from_noc_0_flit_bits_payload)) begin
          $fwrite(32'h80000002,
            "Assertion failed: out[0] incorrect payload\n    at TestHarness.scala:202 assert(rob_payload(rob_idx).asUInt === o.flit.bits.payload.asUInt, cf\"out[${i.toString}] incorrect payload\");\n"
            ); // @[TestHarness.scala 202:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_7953 & ~(io_from_noc_0_flit_bits_ingress_id == _GEN_4608)) begin
          $fwrite(32'h80000002,
            "Assertion failed: out[0] incorrect source\n    at TestHarness.scala:203 assert(o.flit.bits.ingress_id === rob_ingress_id(rob_idx), cf\"out[${i.toString}] incorrect source\")\n"
            ); // @[TestHarness.scala 203:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_7953 & ~(~_GEN_4736)) begin
          $fwrite(32'h80000002,
            "Assertion failed: out[0] incorrect destination\n    at TestHarness.scala:204 assert(i.U === rob_egress_id(rob_idx), cf\"out[${i.toString}] incorrect destination\")\n"
            ); // @[TestHarness.scala 204:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_7953 & ~(_GEN_4864 < _GEN_4992)) begin
          $fwrite(32'h80000002,
            "Assertion failed: out[0] too many flits returned\n    at TestHarness.scala:205 assert(rob_flits_returned(rob_idx) < rob_n_flits(rob_idx), cf\"out[${i.toString}] too many flits returned\")\n"
            ); // @[TestHarness.scala 205:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_7953 & ~(~packet_valid & io_from_noc_0_flit_bits_head | out_payload_rob_idx == _GEN_7819)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at TestHarness.scala:206 assert((!packet_valid && o.flit.bits.head) || rob_idx === packet_rob_idx)\n"
            ); // @[TestHarness.scala 206:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_84 & _T_76 & _T_3) begin
          $fwrite(32'h80000002,"%d, 0, %d\n",_GEN_4608,tsc - out_payload_tsc); // @[TestHarness.scala 210:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_131 & _T_3 & ~_T_89[0]) begin
          $fwrite(32'h80000002,
            "Assertion failed: out[1] unexpected response\n    at TestHarness.scala:201 assert(rob_valids(rob_idx), cf\"out[${i.toString}] unexpected response\")\n"
            ); // @[TestHarness.scala 201:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_7960 & ~(_T_95 == io_from_noc_1_flit_bits_payload)) begin
          $fwrite(32'h80000002,
            "Assertion failed: out[1] incorrect payload\n    at TestHarness.scala:202 assert(rob_payload(rob_idx).asUInt === o.flit.bits.payload.asUInt, cf\"out[${i.toString}] incorrect payload\");\n"
            ); // @[TestHarness.scala 202:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_7960 & ~(io_from_noc_1_flit_bits_ingress_id == _GEN_6405)) begin
          $fwrite(32'h80000002,
            "Assertion failed: out[1] incorrect source\n    at TestHarness.scala:203 assert(o.flit.bits.ingress_id === rob_ingress_id(rob_idx), cf\"out[${i.toString}] incorrect source\")\n"
            ); // @[TestHarness.scala 203:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_7960 & ~_GEN_6533) begin
          $fwrite(32'h80000002,
            "Assertion failed: out[1] incorrect destination\n    at TestHarness.scala:204 assert(i.U === rob_egress_id(rob_idx), cf\"out[${i.toString}] incorrect destination\")\n"
            ); // @[TestHarness.scala 204:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_7960 & ~(_GEN_6661 < _GEN_6789)) begin
          $fwrite(32'h80000002,
            "Assertion failed: out[1] too many flits returned\n    at TestHarness.scala:205 assert(rob_flits_returned(rob_idx) < rob_n_flits(rob_idx), cf\"out[${i.toString}] too many flits returned\")\n"
            ); // @[TestHarness.scala 205:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_7960 & ~(~packet_valid_1 & io_from_noc_1_flit_bits_head | out_payload_1_rob_idx == _GEN_7820)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at TestHarness.scala:206 assert((!packet_valid && o.flit.bits.head) || rob_idx === packet_rob_idx)\n"
            ); // @[TestHarness.scala 206:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_131 & _T_123 & _T_3) begin
          $fwrite(32'h80000002,"%d, 1, %d\n",_GEN_6405,tsc - out_payload_1_tsc); // @[TestHarness.scala 210:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[0] & _T_3 & ~(_T_136 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 0 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[1] & _T_3 & ~(_T_143 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 1 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[2] & _T_3 & ~(_T_150 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 2 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[3] & _T_3 & ~(_T_157 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 3 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[4] & _T_3 & ~(_T_164 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 4 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[5] & _T_3 & ~(_T_171 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 5 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[6] & _T_3 & ~(_T_178 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 6 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[7] & _T_3 & ~(_T_185 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 7 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[8] & _T_3 & ~(_T_192 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 8 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[9] & _T_3 & ~(_T_199 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 9 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[10] & _T_3 & ~(_T_206 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 10 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[11] & _T_3 & ~(_T_213 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 11 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[12] & _T_3 & ~(_T_220 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 12 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[13] & _T_3 & ~(_T_227 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 13 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[14] & _T_3 & ~(_T_234 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 14 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[15] & _T_3 & ~(_T_241 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 15 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[16] & _T_3 & ~(_T_248 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 16 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[17] & _T_3 & ~(_T_255 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 17 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[18] & _T_3 & ~(_T_262 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 18 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[19] & _T_3 & ~(_T_269 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 19 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[20] & _T_3 & ~(_T_276 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 20 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[21] & _T_3 & ~(_T_283 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 21 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[22] & _T_3 & ~(_T_290 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 22 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[23] & _T_3 & ~(_T_297 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 23 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[24] & _T_3 & ~(_T_304 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 24 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[25] & _T_3 & ~(_T_311 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 25 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[26] & _T_3 & ~(_T_318 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 26 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[27] & _T_3 & ~(_T_325 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 27 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[28] & _T_3 & ~(_T_332 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 28 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[29] & _T_3 & ~(_T_339 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 29 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[30] & _T_3 & ~(_T_346 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 30 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[31] & _T_3 & ~(_T_353 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 31 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[32] & _T_3 & ~(_T_360 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 32 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[33] & _T_3 & ~(_T_367 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 33 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[34] & _T_3 & ~(_T_374 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 34 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[35] & _T_3 & ~(_T_381 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 35 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[36] & _T_3 & ~(_T_388 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 36 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[37] & _T_3 & ~(_T_395 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 37 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[38] & _T_3 & ~(_T_402 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 38 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[39] & _T_3 & ~(_T_409 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 39 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[40] & _T_3 & ~(_T_416 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 40 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[41] & _T_3 & ~(_T_423 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 41 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[42] & _T_3 & ~(_T_430 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 42 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[43] & _T_3 & ~(_T_437 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 43 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[44] & _T_3 & ~(_T_444 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 44 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[45] & _T_3 & ~(_T_451 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 45 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[46] & _T_3 & ~(_T_458 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 46 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[47] & _T_3 & ~(_T_465 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 47 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[48] & _T_3 & ~(_T_472 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 48 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[49] & _T_3 & ~(_T_479 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 49 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[50] & _T_3 & ~(_T_486 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 50 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[51] & _T_3 & ~(_T_493 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 51 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[52] & _T_3 & ~(_T_500 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 52 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[53] & _T_3 & ~(_T_507 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 53 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[54] & _T_3 & ~(_T_514 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 54 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[55] & _T_3 & ~(_T_521 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 55 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[56] & _T_3 & ~(_T_528 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 56 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[57] & _T_3 & ~(_T_535 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 57 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[58] & _T_3 & ~(_T_542 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 58 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[59] & _T_3 & ~(_T_549 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 59 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[60] & _T_3 & ~(_T_556 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 60 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[61] & _T_3 & ~(_T_563 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 61 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[62] & _T_3 & ~(_T_570 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 62 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[63] & _T_3 & ~(_T_577 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 63 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[64] & _T_3 & ~(_T_584 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 64 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[65] & _T_3 & ~(_T_591 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 65 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[66] & _T_3 & ~(_T_598 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 66 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[67] & _T_3 & ~(_T_605 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 67 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[68] & _T_3 & ~(_T_612 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 68 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[69] & _T_3 & ~(_T_619 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 69 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[70] & _T_3 & ~(_T_626 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 70 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[71] & _T_3 & ~(_T_633 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 71 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[72] & _T_3 & ~(_T_640 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 72 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[73] & _T_3 & ~(_T_647 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 73 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[74] & _T_3 & ~(_T_654 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 74 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[75] & _T_3 & ~(_T_661 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 75 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[76] & _T_3 & ~(_T_668 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 76 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[77] & _T_3 & ~(_T_675 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 77 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[78] & _T_3 & ~(_T_682 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 78 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[79] & _T_3 & ~(_T_689 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 79 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[80] & _T_3 & ~(_T_696 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 80 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[81] & _T_3 & ~(_T_703 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 81 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[82] & _T_3 & ~(_T_710 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 82 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[83] & _T_3 & ~(_T_717 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 83 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[84] & _T_3 & ~(_T_724 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 84 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[85] & _T_3 & ~(_T_731 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 85 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[86] & _T_3 & ~(_T_738 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 86 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[87] & _T_3 & ~(_T_745 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 87 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[88] & _T_3 & ~(_T_752 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 88 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[89] & _T_3 & ~(_T_759 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 89 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[90] & _T_3 & ~(_T_766 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 90 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[91] & _T_3 & ~(_T_773 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 91 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[92] & _T_3 & ~(_T_780 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 92 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[93] & _T_3 & ~(_T_787 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 93 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[94] & _T_3 & ~(_T_794 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 94 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[95] & _T_3 & ~(_T_801 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 95 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[96] & _T_3 & ~(_T_808 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 96 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[97] & _T_3 & ~(_T_815 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 97 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[98] & _T_3 & ~(_T_822 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 98 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[99] & _T_3 & ~(_T_829 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 99 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[100] & _T_3 & ~(_T_836 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 100 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[101] & _T_3 & ~(_T_843 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 101 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[102] & _T_3 & ~(_T_850 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 102 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[103] & _T_3 & ~(_T_857 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 103 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[104] & _T_3 & ~(_T_864 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 104 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[105] & _T_3 & ~(_T_871 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 105 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[106] & _T_3 & ~(_T_878 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 106 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[107] & _T_3 & ~(_T_885 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 107 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[108] & _T_3 & ~(_T_892 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 108 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[109] & _T_3 & ~(_T_899 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 109 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[110] & _T_3 & ~(_T_906 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 110 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[111] & _T_3 & ~(_T_913 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 111 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[112] & _T_3 & ~(_T_920 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 112 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[113] & _T_3 & ~(_T_927 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 113 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[114] & _T_3 & ~(_T_934 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 114 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[115] & _T_3 & ~(_T_941 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 115 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[116] & _T_3 & ~(_T_948 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 116 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[117] & _T_3 & ~(_T_955 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 117 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[118] & _T_3 & ~(_T_962 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 118 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[119] & _T_3 & ~(_T_969 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 119 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[120] & _T_3 & ~(_T_976 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 120 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[121] & _T_3 & ~(_T_983 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 121 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[122] & _T_3 & ~(_T_990 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 122 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[123] & _T_3 & ~(_T_997 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 123 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[124] & _T_3 & ~(_T_1004 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 124 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[125] & _T_3 & ~(_T_1011 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 125 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[126] & _T_3 & ~(_T_1018 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 126 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rob_valids[127] & _T_3 & ~(_T_1025 < 64'h4000)) begin
          $fwrite(32'h80000002,
            "Assertion failed: ROB Entry 127 took too long\n    at TestHarness.scala:229 assert(tsc - rob_tscs(i) < (16 << 10).U, cf\"ROB Entry ${i.toString} took too long\")\n"
            ); // @[TestHarness.scala 229:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  txs = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  flits = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  tsc = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  idle_counter = _RAND_3[10:0];
  _RAND_4 = {4{`RANDOM}};
  rob_valids = _RAND_4[127:0];
  _RAND_5 = {1{`RANDOM}};
  rob_payload_0_tsc = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  rob_payload_0_rob_idx = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  rob_payload_0_flits_fired = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  rob_payload_1_tsc = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  rob_payload_1_rob_idx = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  rob_payload_1_flits_fired = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  rob_payload_2_tsc = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  rob_payload_2_rob_idx = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  rob_payload_2_flits_fired = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  rob_payload_3_tsc = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  rob_payload_3_rob_idx = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  rob_payload_3_flits_fired = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  rob_payload_4_tsc = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  rob_payload_4_rob_idx = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  rob_payload_4_flits_fired = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  rob_payload_5_tsc = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  rob_payload_5_rob_idx = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  rob_payload_5_flits_fired = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  rob_payload_6_tsc = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  rob_payload_6_rob_idx = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  rob_payload_6_flits_fired = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  rob_payload_7_tsc = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  rob_payload_7_rob_idx = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  rob_payload_7_flits_fired = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  rob_payload_8_tsc = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  rob_payload_8_rob_idx = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  rob_payload_8_flits_fired = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  rob_payload_9_tsc = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  rob_payload_9_rob_idx = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  rob_payload_9_flits_fired = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  rob_payload_10_tsc = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  rob_payload_10_rob_idx = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  rob_payload_10_flits_fired = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  rob_payload_11_tsc = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  rob_payload_11_rob_idx = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  rob_payload_11_flits_fired = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  rob_payload_12_tsc = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  rob_payload_12_rob_idx = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  rob_payload_12_flits_fired = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  rob_payload_13_tsc = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  rob_payload_13_rob_idx = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  rob_payload_13_flits_fired = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  rob_payload_14_tsc = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  rob_payload_14_rob_idx = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  rob_payload_14_flits_fired = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  rob_payload_15_tsc = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  rob_payload_15_rob_idx = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  rob_payload_15_flits_fired = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  rob_payload_16_tsc = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  rob_payload_16_rob_idx = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  rob_payload_16_flits_fired = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  rob_payload_17_tsc = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  rob_payload_17_rob_idx = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  rob_payload_17_flits_fired = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  rob_payload_18_tsc = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  rob_payload_18_rob_idx = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  rob_payload_18_flits_fired = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  rob_payload_19_tsc = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  rob_payload_19_rob_idx = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  rob_payload_19_flits_fired = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  rob_payload_20_tsc = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  rob_payload_20_rob_idx = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  rob_payload_20_flits_fired = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  rob_payload_21_tsc = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  rob_payload_21_rob_idx = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  rob_payload_21_flits_fired = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  rob_payload_22_tsc = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  rob_payload_22_rob_idx = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  rob_payload_22_flits_fired = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  rob_payload_23_tsc = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  rob_payload_23_rob_idx = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  rob_payload_23_flits_fired = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  rob_payload_24_tsc = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  rob_payload_24_rob_idx = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  rob_payload_24_flits_fired = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  rob_payload_25_tsc = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  rob_payload_25_rob_idx = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  rob_payload_25_flits_fired = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  rob_payload_26_tsc = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  rob_payload_26_rob_idx = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  rob_payload_26_flits_fired = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  rob_payload_27_tsc = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  rob_payload_27_rob_idx = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  rob_payload_27_flits_fired = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  rob_payload_28_tsc = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  rob_payload_28_rob_idx = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  rob_payload_28_flits_fired = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  rob_payload_29_tsc = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  rob_payload_29_rob_idx = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  rob_payload_29_flits_fired = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  rob_payload_30_tsc = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  rob_payload_30_rob_idx = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  rob_payload_30_flits_fired = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  rob_payload_31_tsc = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  rob_payload_31_rob_idx = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  rob_payload_31_flits_fired = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  rob_payload_32_tsc = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  rob_payload_32_rob_idx = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  rob_payload_32_flits_fired = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  rob_payload_33_tsc = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  rob_payload_33_rob_idx = _RAND_105[15:0];
  _RAND_106 = {1{`RANDOM}};
  rob_payload_33_flits_fired = _RAND_106[15:0];
  _RAND_107 = {1{`RANDOM}};
  rob_payload_34_tsc = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  rob_payload_34_rob_idx = _RAND_108[15:0];
  _RAND_109 = {1{`RANDOM}};
  rob_payload_34_flits_fired = _RAND_109[15:0];
  _RAND_110 = {1{`RANDOM}};
  rob_payload_35_tsc = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  rob_payload_35_rob_idx = _RAND_111[15:0];
  _RAND_112 = {1{`RANDOM}};
  rob_payload_35_flits_fired = _RAND_112[15:0];
  _RAND_113 = {1{`RANDOM}};
  rob_payload_36_tsc = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  rob_payload_36_rob_idx = _RAND_114[15:0];
  _RAND_115 = {1{`RANDOM}};
  rob_payload_36_flits_fired = _RAND_115[15:0];
  _RAND_116 = {1{`RANDOM}};
  rob_payload_37_tsc = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  rob_payload_37_rob_idx = _RAND_117[15:0];
  _RAND_118 = {1{`RANDOM}};
  rob_payload_37_flits_fired = _RAND_118[15:0];
  _RAND_119 = {1{`RANDOM}};
  rob_payload_38_tsc = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  rob_payload_38_rob_idx = _RAND_120[15:0];
  _RAND_121 = {1{`RANDOM}};
  rob_payload_38_flits_fired = _RAND_121[15:0];
  _RAND_122 = {1{`RANDOM}};
  rob_payload_39_tsc = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  rob_payload_39_rob_idx = _RAND_123[15:0];
  _RAND_124 = {1{`RANDOM}};
  rob_payload_39_flits_fired = _RAND_124[15:0];
  _RAND_125 = {1{`RANDOM}};
  rob_payload_40_tsc = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  rob_payload_40_rob_idx = _RAND_126[15:0];
  _RAND_127 = {1{`RANDOM}};
  rob_payload_40_flits_fired = _RAND_127[15:0];
  _RAND_128 = {1{`RANDOM}};
  rob_payload_41_tsc = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  rob_payload_41_rob_idx = _RAND_129[15:0];
  _RAND_130 = {1{`RANDOM}};
  rob_payload_41_flits_fired = _RAND_130[15:0];
  _RAND_131 = {1{`RANDOM}};
  rob_payload_42_tsc = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  rob_payload_42_rob_idx = _RAND_132[15:0];
  _RAND_133 = {1{`RANDOM}};
  rob_payload_42_flits_fired = _RAND_133[15:0];
  _RAND_134 = {1{`RANDOM}};
  rob_payload_43_tsc = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  rob_payload_43_rob_idx = _RAND_135[15:0];
  _RAND_136 = {1{`RANDOM}};
  rob_payload_43_flits_fired = _RAND_136[15:0];
  _RAND_137 = {1{`RANDOM}};
  rob_payload_44_tsc = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  rob_payload_44_rob_idx = _RAND_138[15:0];
  _RAND_139 = {1{`RANDOM}};
  rob_payload_44_flits_fired = _RAND_139[15:0];
  _RAND_140 = {1{`RANDOM}};
  rob_payload_45_tsc = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  rob_payload_45_rob_idx = _RAND_141[15:0];
  _RAND_142 = {1{`RANDOM}};
  rob_payload_45_flits_fired = _RAND_142[15:0];
  _RAND_143 = {1{`RANDOM}};
  rob_payload_46_tsc = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  rob_payload_46_rob_idx = _RAND_144[15:0];
  _RAND_145 = {1{`RANDOM}};
  rob_payload_46_flits_fired = _RAND_145[15:0];
  _RAND_146 = {1{`RANDOM}};
  rob_payload_47_tsc = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  rob_payload_47_rob_idx = _RAND_147[15:0];
  _RAND_148 = {1{`RANDOM}};
  rob_payload_47_flits_fired = _RAND_148[15:0];
  _RAND_149 = {1{`RANDOM}};
  rob_payload_48_tsc = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  rob_payload_48_rob_idx = _RAND_150[15:0];
  _RAND_151 = {1{`RANDOM}};
  rob_payload_48_flits_fired = _RAND_151[15:0];
  _RAND_152 = {1{`RANDOM}};
  rob_payload_49_tsc = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  rob_payload_49_rob_idx = _RAND_153[15:0];
  _RAND_154 = {1{`RANDOM}};
  rob_payload_49_flits_fired = _RAND_154[15:0];
  _RAND_155 = {1{`RANDOM}};
  rob_payload_50_tsc = _RAND_155[31:0];
  _RAND_156 = {1{`RANDOM}};
  rob_payload_50_rob_idx = _RAND_156[15:0];
  _RAND_157 = {1{`RANDOM}};
  rob_payload_50_flits_fired = _RAND_157[15:0];
  _RAND_158 = {1{`RANDOM}};
  rob_payload_51_tsc = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  rob_payload_51_rob_idx = _RAND_159[15:0];
  _RAND_160 = {1{`RANDOM}};
  rob_payload_51_flits_fired = _RAND_160[15:0];
  _RAND_161 = {1{`RANDOM}};
  rob_payload_52_tsc = _RAND_161[31:0];
  _RAND_162 = {1{`RANDOM}};
  rob_payload_52_rob_idx = _RAND_162[15:0];
  _RAND_163 = {1{`RANDOM}};
  rob_payload_52_flits_fired = _RAND_163[15:0];
  _RAND_164 = {1{`RANDOM}};
  rob_payload_53_tsc = _RAND_164[31:0];
  _RAND_165 = {1{`RANDOM}};
  rob_payload_53_rob_idx = _RAND_165[15:0];
  _RAND_166 = {1{`RANDOM}};
  rob_payload_53_flits_fired = _RAND_166[15:0];
  _RAND_167 = {1{`RANDOM}};
  rob_payload_54_tsc = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  rob_payload_54_rob_idx = _RAND_168[15:0];
  _RAND_169 = {1{`RANDOM}};
  rob_payload_54_flits_fired = _RAND_169[15:0];
  _RAND_170 = {1{`RANDOM}};
  rob_payload_55_tsc = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  rob_payload_55_rob_idx = _RAND_171[15:0];
  _RAND_172 = {1{`RANDOM}};
  rob_payload_55_flits_fired = _RAND_172[15:0];
  _RAND_173 = {1{`RANDOM}};
  rob_payload_56_tsc = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  rob_payload_56_rob_idx = _RAND_174[15:0];
  _RAND_175 = {1{`RANDOM}};
  rob_payload_56_flits_fired = _RAND_175[15:0];
  _RAND_176 = {1{`RANDOM}};
  rob_payload_57_tsc = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  rob_payload_57_rob_idx = _RAND_177[15:0];
  _RAND_178 = {1{`RANDOM}};
  rob_payload_57_flits_fired = _RAND_178[15:0];
  _RAND_179 = {1{`RANDOM}};
  rob_payload_58_tsc = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  rob_payload_58_rob_idx = _RAND_180[15:0];
  _RAND_181 = {1{`RANDOM}};
  rob_payload_58_flits_fired = _RAND_181[15:0];
  _RAND_182 = {1{`RANDOM}};
  rob_payload_59_tsc = _RAND_182[31:0];
  _RAND_183 = {1{`RANDOM}};
  rob_payload_59_rob_idx = _RAND_183[15:0];
  _RAND_184 = {1{`RANDOM}};
  rob_payload_59_flits_fired = _RAND_184[15:0];
  _RAND_185 = {1{`RANDOM}};
  rob_payload_60_tsc = _RAND_185[31:0];
  _RAND_186 = {1{`RANDOM}};
  rob_payload_60_rob_idx = _RAND_186[15:0];
  _RAND_187 = {1{`RANDOM}};
  rob_payload_60_flits_fired = _RAND_187[15:0];
  _RAND_188 = {1{`RANDOM}};
  rob_payload_61_tsc = _RAND_188[31:0];
  _RAND_189 = {1{`RANDOM}};
  rob_payload_61_rob_idx = _RAND_189[15:0];
  _RAND_190 = {1{`RANDOM}};
  rob_payload_61_flits_fired = _RAND_190[15:0];
  _RAND_191 = {1{`RANDOM}};
  rob_payload_62_tsc = _RAND_191[31:0];
  _RAND_192 = {1{`RANDOM}};
  rob_payload_62_rob_idx = _RAND_192[15:0];
  _RAND_193 = {1{`RANDOM}};
  rob_payload_62_flits_fired = _RAND_193[15:0];
  _RAND_194 = {1{`RANDOM}};
  rob_payload_63_tsc = _RAND_194[31:0];
  _RAND_195 = {1{`RANDOM}};
  rob_payload_63_rob_idx = _RAND_195[15:0];
  _RAND_196 = {1{`RANDOM}};
  rob_payload_63_flits_fired = _RAND_196[15:0];
  _RAND_197 = {1{`RANDOM}};
  rob_payload_64_tsc = _RAND_197[31:0];
  _RAND_198 = {1{`RANDOM}};
  rob_payload_64_rob_idx = _RAND_198[15:0];
  _RAND_199 = {1{`RANDOM}};
  rob_payload_64_flits_fired = _RAND_199[15:0];
  _RAND_200 = {1{`RANDOM}};
  rob_payload_65_tsc = _RAND_200[31:0];
  _RAND_201 = {1{`RANDOM}};
  rob_payload_65_rob_idx = _RAND_201[15:0];
  _RAND_202 = {1{`RANDOM}};
  rob_payload_65_flits_fired = _RAND_202[15:0];
  _RAND_203 = {1{`RANDOM}};
  rob_payload_66_tsc = _RAND_203[31:0];
  _RAND_204 = {1{`RANDOM}};
  rob_payload_66_rob_idx = _RAND_204[15:0];
  _RAND_205 = {1{`RANDOM}};
  rob_payload_66_flits_fired = _RAND_205[15:0];
  _RAND_206 = {1{`RANDOM}};
  rob_payload_67_tsc = _RAND_206[31:0];
  _RAND_207 = {1{`RANDOM}};
  rob_payload_67_rob_idx = _RAND_207[15:0];
  _RAND_208 = {1{`RANDOM}};
  rob_payload_67_flits_fired = _RAND_208[15:0];
  _RAND_209 = {1{`RANDOM}};
  rob_payload_68_tsc = _RAND_209[31:0];
  _RAND_210 = {1{`RANDOM}};
  rob_payload_68_rob_idx = _RAND_210[15:0];
  _RAND_211 = {1{`RANDOM}};
  rob_payload_68_flits_fired = _RAND_211[15:0];
  _RAND_212 = {1{`RANDOM}};
  rob_payload_69_tsc = _RAND_212[31:0];
  _RAND_213 = {1{`RANDOM}};
  rob_payload_69_rob_idx = _RAND_213[15:0];
  _RAND_214 = {1{`RANDOM}};
  rob_payload_69_flits_fired = _RAND_214[15:0];
  _RAND_215 = {1{`RANDOM}};
  rob_payload_70_tsc = _RAND_215[31:0];
  _RAND_216 = {1{`RANDOM}};
  rob_payload_70_rob_idx = _RAND_216[15:0];
  _RAND_217 = {1{`RANDOM}};
  rob_payload_70_flits_fired = _RAND_217[15:0];
  _RAND_218 = {1{`RANDOM}};
  rob_payload_71_tsc = _RAND_218[31:0];
  _RAND_219 = {1{`RANDOM}};
  rob_payload_71_rob_idx = _RAND_219[15:0];
  _RAND_220 = {1{`RANDOM}};
  rob_payload_71_flits_fired = _RAND_220[15:0];
  _RAND_221 = {1{`RANDOM}};
  rob_payload_72_tsc = _RAND_221[31:0];
  _RAND_222 = {1{`RANDOM}};
  rob_payload_72_rob_idx = _RAND_222[15:0];
  _RAND_223 = {1{`RANDOM}};
  rob_payload_72_flits_fired = _RAND_223[15:0];
  _RAND_224 = {1{`RANDOM}};
  rob_payload_73_tsc = _RAND_224[31:0];
  _RAND_225 = {1{`RANDOM}};
  rob_payload_73_rob_idx = _RAND_225[15:0];
  _RAND_226 = {1{`RANDOM}};
  rob_payload_73_flits_fired = _RAND_226[15:0];
  _RAND_227 = {1{`RANDOM}};
  rob_payload_74_tsc = _RAND_227[31:0];
  _RAND_228 = {1{`RANDOM}};
  rob_payload_74_rob_idx = _RAND_228[15:0];
  _RAND_229 = {1{`RANDOM}};
  rob_payload_74_flits_fired = _RAND_229[15:0];
  _RAND_230 = {1{`RANDOM}};
  rob_payload_75_tsc = _RAND_230[31:0];
  _RAND_231 = {1{`RANDOM}};
  rob_payload_75_rob_idx = _RAND_231[15:0];
  _RAND_232 = {1{`RANDOM}};
  rob_payload_75_flits_fired = _RAND_232[15:0];
  _RAND_233 = {1{`RANDOM}};
  rob_payload_76_tsc = _RAND_233[31:0];
  _RAND_234 = {1{`RANDOM}};
  rob_payload_76_rob_idx = _RAND_234[15:0];
  _RAND_235 = {1{`RANDOM}};
  rob_payload_76_flits_fired = _RAND_235[15:0];
  _RAND_236 = {1{`RANDOM}};
  rob_payload_77_tsc = _RAND_236[31:0];
  _RAND_237 = {1{`RANDOM}};
  rob_payload_77_rob_idx = _RAND_237[15:0];
  _RAND_238 = {1{`RANDOM}};
  rob_payload_77_flits_fired = _RAND_238[15:0];
  _RAND_239 = {1{`RANDOM}};
  rob_payload_78_tsc = _RAND_239[31:0];
  _RAND_240 = {1{`RANDOM}};
  rob_payload_78_rob_idx = _RAND_240[15:0];
  _RAND_241 = {1{`RANDOM}};
  rob_payload_78_flits_fired = _RAND_241[15:0];
  _RAND_242 = {1{`RANDOM}};
  rob_payload_79_tsc = _RAND_242[31:0];
  _RAND_243 = {1{`RANDOM}};
  rob_payload_79_rob_idx = _RAND_243[15:0];
  _RAND_244 = {1{`RANDOM}};
  rob_payload_79_flits_fired = _RAND_244[15:0];
  _RAND_245 = {1{`RANDOM}};
  rob_payload_80_tsc = _RAND_245[31:0];
  _RAND_246 = {1{`RANDOM}};
  rob_payload_80_rob_idx = _RAND_246[15:0];
  _RAND_247 = {1{`RANDOM}};
  rob_payload_80_flits_fired = _RAND_247[15:0];
  _RAND_248 = {1{`RANDOM}};
  rob_payload_81_tsc = _RAND_248[31:0];
  _RAND_249 = {1{`RANDOM}};
  rob_payload_81_rob_idx = _RAND_249[15:0];
  _RAND_250 = {1{`RANDOM}};
  rob_payload_81_flits_fired = _RAND_250[15:0];
  _RAND_251 = {1{`RANDOM}};
  rob_payload_82_tsc = _RAND_251[31:0];
  _RAND_252 = {1{`RANDOM}};
  rob_payload_82_rob_idx = _RAND_252[15:0];
  _RAND_253 = {1{`RANDOM}};
  rob_payload_82_flits_fired = _RAND_253[15:0];
  _RAND_254 = {1{`RANDOM}};
  rob_payload_83_tsc = _RAND_254[31:0];
  _RAND_255 = {1{`RANDOM}};
  rob_payload_83_rob_idx = _RAND_255[15:0];
  _RAND_256 = {1{`RANDOM}};
  rob_payload_83_flits_fired = _RAND_256[15:0];
  _RAND_257 = {1{`RANDOM}};
  rob_payload_84_tsc = _RAND_257[31:0];
  _RAND_258 = {1{`RANDOM}};
  rob_payload_84_rob_idx = _RAND_258[15:0];
  _RAND_259 = {1{`RANDOM}};
  rob_payload_84_flits_fired = _RAND_259[15:0];
  _RAND_260 = {1{`RANDOM}};
  rob_payload_85_tsc = _RAND_260[31:0];
  _RAND_261 = {1{`RANDOM}};
  rob_payload_85_rob_idx = _RAND_261[15:0];
  _RAND_262 = {1{`RANDOM}};
  rob_payload_85_flits_fired = _RAND_262[15:0];
  _RAND_263 = {1{`RANDOM}};
  rob_payload_86_tsc = _RAND_263[31:0];
  _RAND_264 = {1{`RANDOM}};
  rob_payload_86_rob_idx = _RAND_264[15:0];
  _RAND_265 = {1{`RANDOM}};
  rob_payload_86_flits_fired = _RAND_265[15:0];
  _RAND_266 = {1{`RANDOM}};
  rob_payload_87_tsc = _RAND_266[31:0];
  _RAND_267 = {1{`RANDOM}};
  rob_payload_87_rob_idx = _RAND_267[15:0];
  _RAND_268 = {1{`RANDOM}};
  rob_payload_87_flits_fired = _RAND_268[15:0];
  _RAND_269 = {1{`RANDOM}};
  rob_payload_88_tsc = _RAND_269[31:0];
  _RAND_270 = {1{`RANDOM}};
  rob_payload_88_rob_idx = _RAND_270[15:0];
  _RAND_271 = {1{`RANDOM}};
  rob_payload_88_flits_fired = _RAND_271[15:0];
  _RAND_272 = {1{`RANDOM}};
  rob_payload_89_tsc = _RAND_272[31:0];
  _RAND_273 = {1{`RANDOM}};
  rob_payload_89_rob_idx = _RAND_273[15:0];
  _RAND_274 = {1{`RANDOM}};
  rob_payload_89_flits_fired = _RAND_274[15:0];
  _RAND_275 = {1{`RANDOM}};
  rob_payload_90_tsc = _RAND_275[31:0];
  _RAND_276 = {1{`RANDOM}};
  rob_payload_90_rob_idx = _RAND_276[15:0];
  _RAND_277 = {1{`RANDOM}};
  rob_payload_90_flits_fired = _RAND_277[15:0];
  _RAND_278 = {1{`RANDOM}};
  rob_payload_91_tsc = _RAND_278[31:0];
  _RAND_279 = {1{`RANDOM}};
  rob_payload_91_rob_idx = _RAND_279[15:0];
  _RAND_280 = {1{`RANDOM}};
  rob_payload_91_flits_fired = _RAND_280[15:0];
  _RAND_281 = {1{`RANDOM}};
  rob_payload_92_tsc = _RAND_281[31:0];
  _RAND_282 = {1{`RANDOM}};
  rob_payload_92_rob_idx = _RAND_282[15:0];
  _RAND_283 = {1{`RANDOM}};
  rob_payload_92_flits_fired = _RAND_283[15:0];
  _RAND_284 = {1{`RANDOM}};
  rob_payload_93_tsc = _RAND_284[31:0];
  _RAND_285 = {1{`RANDOM}};
  rob_payload_93_rob_idx = _RAND_285[15:0];
  _RAND_286 = {1{`RANDOM}};
  rob_payload_93_flits_fired = _RAND_286[15:0];
  _RAND_287 = {1{`RANDOM}};
  rob_payload_94_tsc = _RAND_287[31:0];
  _RAND_288 = {1{`RANDOM}};
  rob_payload_94_rob_idx = _RAND_288[15:0];
  _RAND_289 = {1{`RANDOM}};
  rob_payload_94_flits_fired = _RAND_289[15:0];
  _RAND_290 = {1{`RANDOM}};
  rob_payload_95_tsc = _RAND_290[31:0];
  _RAND_291 = {1{`RANDOM}};
  rob_payload_95_rob_idx = _RAND_291[15:0];
  _RAND_292 = {1{`RANDOM}};
  rob_payload_95_flits_fired = _RAND_292[15:0];
  _RAND_293 = {1{`RANDOM}};
  rob_payload_96_tsc = _RAND_293[31:0];
  _RAND_294 = {1{`RANDOM}};
  rob_payload_96_rob_idx = _RAND_294[15:0];
  _RAND_295 = {1{`RANDOM}};
  rob_payload_96_flits_fired = _RAND_295[15:0];
  _RAND_296 = {1{`RANDOM}};
  rob_payload_97_tsc = _RAND_296[31:0];
  _RAND_297 = {1{`RANDOM}};
  rob_payload_97_rob_idx = _RAND_297[15:0];
  _RAND_298 = {1{`RANDOM}};
  rob_payload_97_flits_fired = _RAND_298[15:0];
  _RAND_299 = {1{`RANDOM}};
  rob_payload_98_tsc = _RAND_299[31:0];
  _RAND_300 = {1{`RANDOM}};
  rob_payload_98_rob_idx = _RAND_300[15:0];
  _RAND_301 = {1{`RANDOM}};
  rob_payload_98_flits_fired = _RAND_301[15:0];
  _RAND_302 = {1{`RANDOM}};
  rob_payload_99_tsc = _RAND_302[31:0];
  _RAND_303 = {1{`RANDOM}};
  rob_payload_99_rob_idx = _RAND_303[15:0];
  _RAND_304 = {1{`RANDOM}};
  rob_payload_99_flits_fired = _RAND_304[15:0];
  _RAND_305 = {1{`RANDOM}};
  rob_payload_100_tsc = _RAND_305[31:0];
  _RAND_306 = {1{`RANDOM}};
  rob_payload_100_rob_idx = _RAND_306[15:0];
  _RAND_307 = {1{`RANDOM}};
  rob_payload_100_flits_fired = _RAND_307[15:0];
  _RAND_308 = {1{`RANDOM}};
  rob_payload_101_tsc = _RAND_308[31:0];
  _RAND_309 = {1{`RANDOM}};
  rob_payload_101_rob_idx = _RAND_309[15:0];
  _RAND_310 = {1{`RANDOM}};
  rob_payload_101_flits_fired = _RAND_310[15:0];
  _RAND_311 = {1{`RANDOM}};
  rob_payload_102_tsc = _RAND_311[31:0];
  _RAND_312 = {1{`RANDOM}};
  rob_payload_102_rob_idx = _RAND_312[15:0];
  _RAND_313 = {1{`RANDOM}};
  rob_payload_102_flits_fired = _RAND_313[15:0];
  _RAND_314 = {1{`RANDOM}};
  rob_payload_103_tsc = _RAND_314[31:0];
  _RAND_315 = {1{`RANDOM}};
  rob_payload_103_rob_idx = _RAND_315[15:0];
  _RAND_316 = {1{`RANDOM}};
  rob_payload_103_flits_fired = _RAND_316[15:0];
  _RAND_317 = {1{`RANDOM}};
  rob_payload_104_tsc = _RAND_317[31:0];
  _RAND_318 = {1{`RANDOM}};
  rob_payload_104_rob_idx = _RAND_318[15:0];
  _RAND_319 = {1{`RANDOM}};
  rob_payload_104_flits_fired = _RAND_319[15:0];
  _RAND_320 = {1{`RANDOM}};
  rob_payload_105_tsc = _RAND_320[31:0];
  _RAND_321 = {1{`RANDOM}};
  rob_payload_105_rob_idx = _RAND_321[15:0];
  _RAND_322 = {1{`RANDOM}};
  rob_payload_105_flits_fired = _RAND_322[15:0];
  _RAND_323 = {1{`RANDOM}};
  rob_payload_106_tsc = _RAND_323[31:0];
  _RAND_324 = {1{`RANDOM}};
  rob_payload_106_rob_idx = _RAND_324[15:0];
  _RAND_325 = {1{`RANDOM}};
  rob_payload_106_flits_fired = _RAND_325[15:0];
  _RAND_326 = {1{`RANDOM}};
  rob_payload_107_tsc = _RAND_326[31:0];
  _RAND_327 = {1{`RANDOM}};
  rob_payload_107_rob_idx = _RAND_327[15:0];
  _RAND_328 = {1{`RANDOM}};
  rob_payload_107_flits_fired = _RAND_328[15:0];
  _RAND_329 = {1{`RANDOM}};
  rob_payload_108_tsc = _RAND_329[31:0];
  _RAND_330 = {1{`RANDOM}};
  rob_payload_108_rob_idx = _RAND_330[15:0];
  _RAND_331 = {1{`RANDOM}};
  rob_payload_108_flits_fired = _RAND_331[15:0];
  _RAND_332 = {1{`RANDOM}};
  rob_payload_109_tsc = _RAND_332[31:0];
  _RAND_333 = {1{`RANDOM}};
  rob_payload_109_rob_idx = _RAND_333[15:0];
  _RAND_334 = {1{`RANDOM}};
  rob_payload_109_flits_fired = _RAND_334[15:0];
  _RAND_335 = {1{`RANDOM}};
  rob_payload_110_tsc = _RAND_335[31:0];
  _RAND_336 = {1{`RANDOM}};
  rob_payload_110_rob_idx = _RAND_336[15:0];
  _RAND_337 = {1{`RANDOM}};
  rob_payload_110_flits_fired = _RAND_337[15:0];
  _RAND_338 = {1{`RANDOM}};
  rob_payload_111_tsc = _RAND_338[31:0];
  _RAND_339 = {1{`RANDOM}};
  rob_payload_111_rob_idx = _RAND_339[15:0];
  _RAND_340 = {1{`RANDOM}};
  rob_payload_111_flits_fired = _RAND_340[15:0];
  _RAND_341 = {1{`RANDOM}};
  rob_payload_112_tsc = _RAND_341[31:0];
  _RAND_342 = {1{`RANDOM}};
  rob_payload_112_rob_idx = _RAND_342[15:0];
  _RAND_343 = {1{`RANDOM}};
  rob_payload_112_flits_fired = _RAND_343[15:0];
  _RAND_344 = {1{`RANDOM}};
  rob_payload_113_tsc = _RAND_344[31:0];
  _RAND_345 = {1{`RANDOM}};
  rob_payload_113_rob_idx = _RAND_345[15:0];
  _RAND_346 = {1{`RANDOM}};
  rob_payload_113_flits_fired = _RAND_346[15:0];
  _RAND_347 = {1{`RANDOM}};
  rob_payload_114_tsc = _RAND_347[31:0];
  _RAND_348 = {1{`RANDOM}};
  rob_payload_114_rob_idx = _RAND_348[15:0];
  _RAND_349 = {1{`RANDOM}};
  rob_payload_114_flits_fired = _RAND_349[15:0];
  _RAND_350 = {1{`RANDOM}};
  rob_payload_115_tsc = _RAND_350[31:0];
  _RAND_351 = {1{`RANDOM}};
  rob_payload_115_rob_idx = _RAND_351[15:0];
  _RAND_352 = {1{`RANDOM}};
  rob_payload_115_flits_fired = _RAND_352[15:0];
  _RAND_353 = {1{`RANDOM}};
  rob_payload_116_tsc = _RAND_353[31:0];
  _RAND_354 = {1{`RANDOM}};
  rob_payload_116_rob_idx = _RAND_354[15:0];
  _RAND_355 = {1{`RANDOM}};
  rob_payload_116_flits_fired = _RAND_355[15:0];
  _RAND_356 = {1{`RANDOM}};
  rob_payload_117_tsc = _RAND_356[31:0];
  _RAND_357 = {1{`RANDOM}};
  rob_payload_117_rob_idx = _RAND_357[15:0];
  _RAND_358 = {1{`RANDOM}};
  rob_payload_117_flits_fired = _RAND_358[15:0];
  _RAND_359 = {1{`RANDOM}};
  rob_payload_118_tsc = _RAND_359[31:0];
  _RAND_360 = {1{`RANDOM}};
  rob_payload_118_rob_idx = _RAND_360[15:0];
  _RAND_361 = {1{`RANDOM}};
  rob_payload_118_flits_fired = _RAND_361[15:0];
  _RAND_362 = {1{`RANDOM}};
  rob_payload_119_tsc = _RAND_362[31:0];
  _RAND_363 = {1{`RANDOM}};
  rob_payload_119_rob_idx = _RAND_363[15:0];
  _RAND_364 = {1{`RANDOM}};
  rob_payload_119_flits_fired = _RAND_364[15:0];
  _RAND_365 = {1{`RANDOM}};
  rob_payload_120_tsc = _RAND_365[31:0];
  _RAND_366 = {1{`RANDOM}};
  rob_payload_120_rob_idx = _RAND_366[15:0];
  _RAND_367 = {1{`RANDOM}};
  rob_payload_120_flits_fired = _RAND_367[15:0];
  _RAND_368 = {1{`RANDOM}};
  rob_payload_121_tsc = _RAND_368[31:0];
  _RAND_369 = {1{`RANDOM}};
  rob_payload_121_rob_idx = _RAND_369[15:0];
  _RAND_370 = {1{`RANDOM}};
  rob_payload_121_flits_fired = _RAND_370[15:0];
  _RAND_371 = {1{`RANDOM}};
  rob_payload_122_tsc = _RAND_371[31:0];
  _RAND_372 = {1{`RANDOM}};
  rob_payload_122_rob_idx = _RAND_372[15:0];
  _RAND_373 = {1{`RANDOM}};
  rob_payload_122_flits_fired = _RAND_373[15:0];
  _RAND_374 = {1{`RANDOM}};
  rob_payload_123_tsc = _RAND_374[31:0];
  _RAND_375 = {1{`RANDOM}};
  rob_payload_123_rob_idx = _RAND_375[15:0];
  _RAND_376 = {1{`RANDOM}};
  rob_payload_123_flits_fired = _RAND_376[15:0];
  _RAND_377 = {1{`RANDOM}};
  rob_payload_124_tsc = _RAND_377[31:0];
  _RAND_378 = {1{`RANDOM}};
  rob_payload_124_rob_idx = _RAND_378[15:0];
  _RAND_379 = {1{`RANDOM}};
  rob_payload_124_flits_fired = _RAND_379[15:0];
  _RAND_380 = {1{`RANDOM}};
  rob_payload_125_tsc = _RAND_380[31:0];
  _RAND_381 = {1{`RANDOM}};
  rob_payload_125_rob_idx = _RAND_381[15:0];
  _RAND_382 = {1{`RANDOM}};
  rob_payload_125_flits_fired = _RAND_382[15:0];
  _RAND_383 = {1{`RANDOM}};
  rob_payload_126_tsc = _RAND_383[31:0];
  _RAND_384 = {1{`RANDOM}};
  rob_payload_126_rob_idx = _RAND_384[15:0];
  _RAND_385 = {1{`RANDOM}};
  rob_payload_126_flits_fired = _RAND_385[15:0];
  _RAND_386 = {1{`RANDOM}};
  rob_payload_127_tsc = _RAND_386[31:0];
  _RAND_387 = {1{`RANDOM}};
  rob_payload_127_rob_idx = _RAND_387[15:0];
  _RAND_388 = {1{`RANDOM}};
  rob_payload_127_flits_fired = _RAND_388[15:0];
  _RAND_389 = {1{`RANDOM}};
  rob_egress_id_0 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  rob_egress_id_1 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  rob_egress_id_2 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  rob_egress_id_3 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  rob_egress_id_4 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  rob_egress_id_5 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  rob_egress_id_6 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  rob_egress_id_7 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  rob_egress_id_8 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  rob_egress_id_9 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  rob_egress_id_10 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  rob_egress_id_11 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  rob_egress_id_12 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  rob_egress_id_13 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  rob_egress_id_14 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  rob_egress_id_15 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  rob_egress_id_16 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  rob_egress_id_17 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  rob_egress_id_18 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  rob_egress_id_19 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  rob_egress_id_20 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  rob_egress_id_21 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  rob_egress_id_22 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  rob_egress_id_23 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  rob_egress_id_24 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  rob_egress_id_25 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  rob_egress_id_26 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  rob_egress_id_27 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  rob_egress_id_28 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  rob_egress_id_29 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  rob_egress_id_30 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  rob_egress_id_31 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  rob_egress_id_32 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  rob_egress_id_33 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  rob_egress_id_34 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  rob_egress_id_35 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  rob_egress_id_36 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  rob_egress_id_37 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  rob_egress_id_38 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  rob_egress_id_39 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  rob_egress_id_40 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  rob_egress_id_41 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  rob_egress_id_42 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  rob_egress_id_43 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  rob_egress_id_44 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  rob_egress_id_45 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  rob_egress_id_46 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  rob_egress_id_47 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  rob_egress_id_48 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  rob_egress_id_49 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  rob_egress_id_50 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  rob_egress_id_51 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  rob_egress_id_52 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  rob_egress_id_53 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  rob_egress_id_54 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  rob_egress_id_55 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  rob_egress_id_56 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  rob_egress_id_57 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  rob_egress_id_58 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  rob_egress_id_59 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  rob_egress_id_60 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  rob_egress_id_61 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  rob_egress_id_62 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  rob_egress_id_63 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  rob_egress_id_64 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  rob_egress_id_65 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  rob_egress_id_66 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  rob_egress_id_67 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  rob_egress_id_68 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  rob_egress_id_69 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  rob_egress_id_70 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  rob_egress_id_71 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  rob_egress_id_72 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  rob_egress_id_73 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  rob_egress_id_74 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  rob_egress_id_75 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  rob_egress_id_76 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  rob_egress_id_77 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  rob_egress_id_78 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  rob_egress_id_79 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  rob_egress_id_80 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  rob_egress_id_81 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  rob_egress_id_82 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  rob_egress_id_83 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  rob_egress_id_84 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  rob_egress_id_85 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  rob_egress_id_86 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  rob_egress_id_87 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  rob_egress_id_88 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  rob_egress_id_89 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  rob_egress_id_90 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  rob_egress_id_91 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  rob_egress_id_92 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  rob_egress_id_93 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  rob_egress_id_94 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  rob_egress_id_95 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  rob_egress_id_96 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  rob_egress_id_97 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  rob_egress_id_98 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  rob_egress_id_99 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  rob_egress_id_100 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  rob_egress_id_101 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  rob_egress_id_102 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  rob_egress_id_103 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  rob_egress_id_104 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  rob_egress_id_105 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  rob_egress_id_106 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  rob_egress_id_107 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  rob_egress_id_108 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  rob_egress_id_109 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  rob_egress_id_110 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  rob_egress_id_111 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  rob_egress_id_112 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  rob_egress_id_113 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  rob_egress_id_114 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  rob_egress_id_115 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  rob_egress_id_116 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  rob_egress_id_117 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  rob_egress_id_118 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  rob_egress_id_119 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  rob_egress_id_120 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  rob_egress_id_121 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  rob_egress_id_122 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  rob_egress_id_123 = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  rob_egress_id_124 = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  rob_egress_id_125 = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  rob_egress_id_126 = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  rob_egress_id_127 = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  rob_ingress_id_0 = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  rob_ingress_id_1 = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  rob_ingress_id_2 = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  rob_ingress_id_3 = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  rob_ingress_id_4 = _RAND_521[0:0];
  _RAND_522 = {1{`RANDOM}};
  rob_ingress_id_5 = _RAND_522[0:0];
  _RAND_523 = {1{`RANDOM}};
  rob_ingress_id_6 = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  rob_ingress_id_7 = _RAND_524[0:0];
  _RAND_525 = {1{`RANDOM}};
  rob_ingress_id_8 = _RAND_525[0:0];
  _RAND_526 = {1{`RANDOM}};
  rob_ingress_id_9 = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  rob_ingress_id_10 = _RAND_527[0:0];
  _RAND_528 = {1{`RANDOM}};
  rob_ingress_id_11 = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  rob_ingress_id_12 = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  rob_ingress_id_13 = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  rob_ingress_id_14 = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  rob_ingress_id_15 = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  rob_ingress_id_16 = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  rob_ingress_id_17 = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  rob_ingress_id_18 = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  rob_ingress_id_19 = _RAND_536[0:0];
  _RAND_537 = {1{`RANDOM}};
  rob_ingress_id_20 = _RAND_537[0:0];
  _RAND_538 = {1{`RANDOM}};
  rob_ingress_id_21 = _RAND_538[0:0];
  _RAND_539 = {1{`RANDOM}};
  rob_ingress_id_22 = _RAND_539[0:0];
  _RAND_540 = {1{`RANDOM}};
  rob_ingress_id_23 = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  rob_ingress_id_24 = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  rob_ingress_id_25 = _RAND_542[0:0];
  _RAND_543 = {1{`RANDOM}};
  rob_ingress_id_26 = _RAND_543[0:0];
  _RAND_544 = {1{`RANDOM}};
  rob_ingress_id_27 = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  rob_ingress_id_28 = _RAND_545[0:0];
  _RAND_546 = {1{`RANDOM}};
  rob_ingress_id_29 = _RAND_546[0:0];
  _RAND_547 = {1{`RANDOM}};
  rob_ingress_id_30 = _RAND_547[0:0];
  _RAND_548 = {1{`RANDOM}};
  rob_ingress_id_31 = _RAND_548[0:0];
  _RAND_549 = {1{`RANDOM}};
  rob_ingress_id_32 = _RAND_549[0:0];
  _RAND_550 = {1{`RANDOM}};
  rob_ingress_id_33 = _RAND_550[0:0];
  _RAND_551 = {1{`RANDOM}};
  rob_ingress_id_34 = _RAND_551[0:0];
  _RAND_552 = {1{`RANDOM}};
  rob_ingress_id_35 = _RAND_552[0:0];
  _RAND_553 = {1{`RANDOM}};
  rob_ingress_id_36 = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  rob_ingress_id_37 = _RAND_554[0:0];
  _RAND_555 = {1{`RANDOM}};
  rob_ingress_id_38 = _RAND_555[0:0];
  _RAND_556 = {1{`RANDOM}};
  rob_ingress_id_39 = _RAND_556[0:0];
  _RAND_557 = {1{`RANDOM}};
  rob_ingress_id_40 = _RAND_557[0:0];
  _RAND_558 = {1{`RANDOM}};
  rob_ingress_id_41 = _RAND_558[0:0];
  _RAND_559 = {1{`RANDOM}};
  rob_ingress_id_42 = _RAND_559[0:0];
  _RAND_560 = {1{`RANDOM}};
  rob_ingress_id_43 = _RAND_560[0:0];
  _RAND_561 = {1{`RANDOM}};
  rob_ingress_id_44 = _RAND_561[0:0];
  _RAND_562 = {1{`RANDOM}};
  rob_ingress_id_45 = _RAND_562[0:0];
  _RAND_563 = {1{`RANDOM}};
  rob_ingress_id_46 = _RAND_563[0:0];
  _RAND_564 = {1{`RANDOM}};
  rob_ingress_id_47 = _RAND_564[0:0];
  _RAND_565 = {1{`RANDOM}};
  rob_ingress_id_48 = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  rob_ingress_id_49 = _RAND_566[0:0];
  _RAND_567 = {1{`RANDOM}};
  rob_ingress_id_50 = _RAND_567[0:0];
  _RAND_568 = {1{`RANDOM}};
  rob_ingress_id_51 = _RAND_568[0:0];
  _RAND_569 = {1{`RANDOM}};
  rob_ingress_id_52 = _RAND_569[0:0];
  _RAND_570 = {1{`RANDOM}};
  rob_ingress_id_53 = _RAND_570[0:0];
  _RAND_571 = {1{`RANDOM}};
  rob_ingress_id_54 = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  rob_ingress_id_55 = _RAND_572[0:0];
  _RAND_573 = {1{`RANDOM}};
  rob_ingress_id_56 = _RAND_573[0:0];
  _RAND_574 = {1{`RANDOM}};
  rob_ingress_id_57 = _RAND_574[0:0];
  _RAND_575 = {1{`RANDOM}};
  rob_ingress_id_58 = _RAND_575[0:0];
  _RAND_576 = {1{`RANDOM}};
  rob_ingress_id_59 = _RAND_576[0:0];
  _RAND_577 = {1{`RANDOM}};
  rob_ingress_id_60 = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  rob_ingress_id_61 = _RAND_578[0:0];
  _RAND_579 = {1{`RANDOM}};
  rob_ingress_id_62 = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  rob_ingress_id_63 = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  rob_ingress_id_64 = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  rob_ingress_id_65 = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  rob_ingress_id_66 = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  rob_ingress_id_67 = _RAND_584[0:0];
  _RAND_585 = {1{`RANDOM}};
  rob_ingress_id_68 = _RAND_585[0:0];
  _RAND_586 = {1{`RANDOM}};
  rob_ingress_id_69 = _RAND_586[0:0];
  _RAND_587 = {1{`RANDOM}};
  rob_ingress_id_70 = _RAND_587[0:0];
  _RAND_588 = {1{`RANDOM}};
  rob_ingress_id_71 = _RAND_588[0:0];
  _RAND_589 = {1{`RANDOM}};
  rob_ingress_id_72 = _RAND_589[0:0];
  _RAND_590 = {1{`RANDOM}};
  rob_ingress_id_73 = _RAND_590[0:0];
  _RAND_591 = {1{`RANDOM}};
  rob_ingress_id_74 = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  rob_ingress_id_75 = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  rob_ingress_id_76 = _RAND_593[0:0];
  _RAND_594 = {1{`RANDOM}};
  rob_ingress_id_77 = _RAND_594[0:0];
  _RAND_595 = {1{`RANDOM}};
  rob_ingress_id_78 = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  rob_ingress_id_79 = _RAND_596[0:0];
  _RAND_597 = {1{`RANDOM}};
  rob_ingress_id_80 = _RAND_597[0:0];
  _RAND_598 = {1{`RANDOM}};
  rob_ingress_id_81 = _RAND_598[0:0];
  _RAND_599 = {1{`RANDOM}};
  rob_ingress_id_82 = _RAND_599[0:0];
  _RAND_600 = {1{`RANDOM}};
  rob_ingress_id_83 = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  rob_ingress_id_84 = _RAND_601[0:0];
  _RAND_602 = {1{`RANDOM}};
  rob_ingress_id_85 = _RAND_602[0:0];
  _RAND_603 = {1{`RANDOM}};
  rob_ingress_id_86 = _RAND_603[0:0];
  _RAND_604 = {1{`RANDOM}};
  rob_ingress_id_87 = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  rob_ingress_id_88 = _RAND_605[0:0];
  _RAND_606 = {1{`RANDOM}};
  rob_ingress_id_89 = _RAND_606[0:0];
  _RAND_607 = {1{`RANDOM}};
  rob_ingress_id_90 = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  rob_ingress_id_91 = _RAND_608[0:0];
  _RAND_609 = {1{`RANDOM}};
  rob_ingress_id_92 = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  rob_ingress_id_93 = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  rob_ingress_id_94 = _RAND_611[0:0];
  _RAND_612 = {1{`RANDOM}};
  rob_ingress_id_95 = _RAND_612[0:0];
  _RAND_613 = {1{`RANDOM}};
  rob_ingress_id_96 = _RAND_613[0:0];
  _RAND_614 = {1{`RANDOM}};
  rob_ingress_id_97 = _RAND_614[0:0];
  _RAND_615 = {1{`RANDOM}};
  rob_ingress_id_98 = _RAND_615[0:0];
  _RAND_616 = {1{`RANDOM}};
  rob_ingress_id_99 = _RAND_616[0:0];
  _RAND_617 = {1{`RANDOM}};
  rob_ingress_id_100 = _RAND_617[0:0];
  _RAND_618 = {1{`RANDOM}};
  rob_ingress_id_101 = _RAND_618[0:0];
  _RAND_619 = {1{`RANDOM}};
  rob_ingress_id_102 = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  rob_ingress_id_103 = _RAND_620[0:0];
  _RAND_621 = {1{`RANDOM}};
  rob_ingress_id_104 = _RAND_621[0:0];
  _RAND_622 = {1{`RANDOM}};
  rob_ingress_id_105 = _RAND_622[0:0];
  _RAND_623 = {1{`RANDOM}};
  rob_ingress_id_106 = _RAND_623[0:0];
  _RAND_624 = {1{`RANDOM}};
  rob_ingress_id_107 = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  rob_ingress_id_108 = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  rob_ingress_id_109 = _RAND_626[0:0];
  _RAND_627 = {1{`RANDOM}};
  rob_ingress_id_110 = _RAND_627[0:0];
  _RAND_628 = {1{`RANDOM}};
  rob_ingress_id_111 = _RAND_628[0:0];
  _RAND_629 = {1{`RANDOM}};
  rob_ingress_id_112 = _RAND_629[0:0];
  _RAND_630 = {1{`RANDOM}};
  rob_ingress_id_113 = _RAND_630[0:0];
  _RAND_631 = {1{`RANDOM}};
  rob_ingress_id_114 = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  rob_ingress_id_115 = _RAND_632[0:0];
  _RAND_633 = {1{`RANDOM}};
  rob_ingress_id_116 = _RAND_633[0:0];
  _RAND_634 = {1{`RANDOM}};
  rob_ingress_id_117 = _RAND_634[0:0];
  _RAND_635 = {1{`RANDOM}};
  rob_ingress_id_118 = _RAND_635[0:0];
  _RAND_636 = {1{`RANDOM}};
  rob_ingress_id_119 = _RAND_636[0:0];
  _RAND_637 = {1{`RANDOM}};
  rob_ingress_id_120 = _RAND_637[0:0];
  _RAND_638 = {1{`RANDOM}};
  rob_ingress_id_121 = _RAND_638[0:0];
  _RAND_639 = {1{`RANDOM}};
  rob_ingress_id_122 = _RAND_639[0:0];
  _RAND_640 = {1{`RANDOM}};
  rob_ingress_id_123 = _RAND_640[0:0];
  _RAND_641 = {1{`RANDOM}};
  rob_ingress_id_124 = _RAND_641[0:0];
  _RAND_642 = {1{`RANDOM}};
  rob_ingress_id_125 = _RAND_642[0:0];
  _RAND_643 = {1{`RANDOM}};
  rob_ingress_id_126 = _RAND_643[0:0];
  _RAND_644 = {1{`RANDOM}};
  rob_ingress_id_127 = _RAND_644[0:0];
  _RAND_645 = {1{`RANDOM}};
  rob_n_flits_0 = _RAND_645[3:0];
  _RAND_646 = {1{`RANDOM}};
  rob_n_flits_1 = _RAND_646[3:0];
  _RAND_647 = {1{`RANDOM}};
  rob_n_flits_2 = _RAND_647[3:0];
  _RAND_648 = {1{`RANDOM}};
  rob_n_flits_3 = _RAND_648[3:0];
  _RAND_649 = {1{`RANDOM}};
  rob_n_flits_4 = _RAND_649[3:0];
  _RAND_650 = {1{`RANDOM}};
  rob_n_flits_5 = _RAND_650[3:0];
  _RAND_651 = {1{`RANDOM}};
  rob_n_flits_6 = _RAND_651[3:0];
  _RAND_652 = {1{`RANDOM}};
  rob_n_flits_7 = _RAND_652[3:0];
  _RAND_653 = {1{`RANDOM}};
  rob_n_flits_8 = _RAND_653[3:0];
  _RAND_654 = {1{`RANDOM}};
  rob_n_flits_9 = _RAND_654[3:0];
  _RAND_655 = {1{`RANDOM}};
  rob_n_flits_10 = _RAND_655[3:0];
  _RAND_656 = {1{`RANDOM}};
  rob_n_flits_11 = _RAND_656[3:0];
  _RAND_657 = {1{`RANDOM}};
  rob_n_flits_12 = _RAND_657[3:0];
  _RAND_658 = {1{`RANDOM}};
  rob_n_flits_13 = _RAND_658[3:0];
  _RAND_659 = {1{`RANDOM}};
  rob_n_flits_14 = _RAND_659[3:0];
  _RAND_660 = {1{`RANDOM}};
  rob_n_flits_15 = _RAND_660[3:0];
  _RAND_661 = {1{`RANDOM}};
  rob_n_flits_16 = _RAND_661[3:0];
  _RAND_662 = {1{`RANDOM}};
  rob_n_flits_17 = _RAND_662[3:0];
  _RAND_663 = {1{`RANDOM}};
  rob_n_flits_18 = _RAND_663[3:0];
  _RAND_664 = {1{`RANDOM}};
  rob_n_flits_19 = _RAND_664[3:0];
  _RAND_665 = {1{`RANDOM}};
  rob_n_flits_20 = _RAND_665[3:0];
  _RAND_666 = {1{`RANDOM}};
  rob_n_flits_21 = _RAND_666[3:0];
  _RAND_667 = {1{`RANDOM}};
  rob_n_flits_22 = _RAND_667[3:0];
  _RAND_668 = {1{`RANDOM}};
  rob_n_flits_23 = _RAND_668[3:0];
  _RAND_669 = {1{`RANDOM}};
  rob_n_flits_24 = _RAND_669[3:0];
  _RAND_670 = {1{`RANDOM}};
  rob_n_flits_25 = _RAND_670[3:0];
  _RAND_671 = {1{`RANDOM}};
  rob_n_flits_26 = _RAND_671[3:0];
  _RAND_672 = {1{`RANDOM}};
  rob_n_flits_27 = _RAND_672[3:0];
  _RAND_673 = {1{`RANDOM}};
  rob_n_flits_28 = _RAND_673[3:0];
  _RAND_674 = {1{`RANDOM}};
  rob_n_flits_29 = _RAND_674[3:0];
  _RAND_675 = {1{`RANDOM}};
  rob_n_flits_30 = _RAND_675[3:0];
  _RAND_676 = {1{`RANDOM}};
  rob_n_flits_31 = _RAND_676[3:0];
  _RAND_677 = {1{`RANDOM}};
  rob_n_flits_32 = _RAND_677[3:0];
  _RAND_678 = {1{`RANDOM}};
  rob_n_flits_33 = _RAND_678[3:0];
  _RAND_679 = {1{`RANDOM}};
  rob_n_flits_34 = _RAND_679[3:0];
  _RAND_680 = {1{`RANDOM}};
  rob_n_flits_35 = _RAND_680[3:0];
  _RAND_681 = {1{`RANDOM}};
  rob_n_flits_36 = _RAND_681[3:0];
  _RAND_682 = {1{`RANDOM}};
  rob_n_flits_37 = _RAND_682[3:0];
  _RAND_683 = {1{`RANDOM}};
  rob_n_flits_38 = _RAND_683[3:0];
  _RAND_684 = {1{`RANDOM}};
  rob_n_flits_39 = _RAND_684[3:0];
  _RAND_685 = {1{`RANDOM}};
  rob_n_flits_40 = _RAND_685[3:0];
  _RAND_686 = {1{`RANDOM}};
  rob_n_flits_41 = _RAND_686[3:0];
  _RAND_687 = {1{`RANDOM}};
  rob_n_flits_42 = _RAND_687[3:0];
  _RAND_688 = {1{`RANDOM}};
  rob_n_flits_43 = _RAND_688[3:0];
  _RAND_689 = {1{`RANDOM}};
  rob_n_flits_44 = _RAND_689[3:0];
  _RAND_690 = {1{`RANDOM}};
  rob_n_flits_45 = _RAND_690[3:0];
  _RAND_691 = {1{`RANDOM}};
  rob_n_flits_46 = _RAND_691[3:0];
  _RAND_692 = {1{`RANDOM}};
  rob_n_flits_47 = _RAND_692[3:0];
  _RAND_693 = {1{`RANDOM}};
  rob_n_flits_48 = _RAND_693[3:0];
  _RAND_694 = {1{`RANDOM}};
  rob_n_flits_49 = _RAND_694[3:0];
  _RAND_695 = {1{`RANDOM}};
  rob_n_flits_50 = _RAND_695[3:0];
  _RAND_696 = {1{`RANDOM}};
  rob_n_flits_51 = _RAND_696[3:0];
  _RAND_697 = {1{`RANDOM}};
  rob_n_flits_52 = _RAND_697[3:0];
  _RAND_698 = {1{`RANDOM}};
  rob_n_flits_53 = _RAND_698[3:0];
  _RAND_699 = {1{`RANDOM}};
  rob_n_flits_54 = _RAND_699[3:0];
  _RAND_700 = {1{`RANDOM}};
  rob_n_flits_55 = _RAND_700[3:0];
  _RAND_701 = {1{`RANDOM}};
  rob_n_flits_56 = _RAND_701[3:0];
  _RAND_702 = {1{`RANDOM}};
  rob_n_flits_57 = _RAND_702[3:0];
  _RAND_703 = {1{`RANDOM}};
  rob_n_flits_58 = _RAND_703[3:0];
  _RAND_704 = {1{`RANDOM}};
  rob_n_flits_59 = _RAND_704[3:0];
  _RAND_705 = {1{`RANDOM}};
  rob_n_flits_60 = _RAND_705[3:0];
  _RAND_706 = {1{`RANDOM}};
  rob_n_flits_61 = _RAND_706[3:0];
  _RAND_707 = {1{`RANDOM}};
  rob_n_flits_62 = _RAND_707[3:0];
  _RAND_708 = {1{`RANDOM}};
  rob_n_flits_63 = _RAND_708[3:0];
  _RAND_709 = {1{`RANDOM}};
  rob_n_flits_64 = _RAND_709[3:0];
  _RAND_710 = {1{`RANDOM}};
  rob_n_flits_65 = _RAND_710[3:0];
  _RAND_711 = {1{`RANDOM}};
  rob_n_flits_66 = _RAND_711[3:0];
  _RAND_712 = {1{`RANDOM}};
  rob_n_flits_67 = _RAND_712[3:0];
  _RAND_713 = {1{`RANDOM}};
  rob_n_flits_68 = _RAND_713[3:0];
  _RAND_714 = {1{`RANDOM}};
  rob_n_flits_69 = _RAND_714[3:0];
  _RAND_715 = {1{`RANDOM}};
  rob_n_flits_70 = _RAND_715[3:0];
  _RAND_716 = {1{`RANDOM}};
  rob_n_flits_71 = _RAND_716[3:0];
  _RAND_717 = {1{`RANDOM}};
  rob_n_flits_72 = _RAND_717[3:0];
  _RAND_718 = {1{`RANDOM}};
  rob_n_flits_73 = _RAND_718[3:0];
  _RAND_719 = {1{`RANDOM}};
  rob_n_flits_74 = _RAND_719[3:0];
  _RAND_720 = {1{`RANDOM}};
  rob_n_flits_75 = _RAND_720[3:0];
  _RAND_721 = {1{`RANDOM}};
  rob_n_flits_76 = _RAND_721[3:0];
  _RAND_722 = {1{`RANDOM}};
  rob_n_flits_77 = _RAND_722[3:0];
  _RAND_723 = {1{`RANDOM}};
  rob_n_flits_78 = _RAND_723[3:0];
  _RAND_724 = {1{`RANDOM}};
  rob_n_flits_79 = _RAND_724[3:0];
  _RAND_725 = {1{`RANDOM}};
  rob_n_flits_80 = _RAND_725[3:0];
  _RAND_726 = {1{`RANDOM}};
  rob_n_flits_81 = _RAND_726[3:0];
  _RAND_727 = {1{`RANDOM}};
  rob_n_flits_82 = _RAND_727[3:0];
  _RAND_728 = {1{`RANDOM}};
  rob_n_flits_83 = _RAND_728[3:0];
  _RAND_729 = {1{`RANDOM}};
  rob_n_flits_84 = _RAND_729[3:0];
  _RAND_730 = {1{`RANDOM}};
  rob_n_flits_85 = _RAND_730[3:0];
  _RAND_731 = {1{`RANDOM}};
  rob_n_flits_86 = _RAND_731[3:0];
  _RAND_732 = {1{`RANDOM}};
  rob_n_flits_87 = _RAND_732[3:0];
  _RAND_733 = {1{`RANDOM}};
  rob_n_flits_88 = _RAND_733[3:0];
  _RAND_734 = {1{`RANDOM}};
  rob_n_flits_89 = _RAND_734[3:0];
  _RAND_735 = {1{`RANDOM}};
  rob_n_flits_90 = _RAND_735[3:0];
  _RAND_736 = {1{`RANDOM}};
  rob_n_flits_91 = _RAND_736[3:0];
  _RAND_737 = {1{`RANDOM}};
  rob_n_flits_92 = _RAND_737[3:0];
  _RAND_738 = {1{`RANDOM}};
  rob_n_flits_93 = _RAND_738[3:0];
  _RAND_739 = {1{`RANDOM}};
  rob_n_flits_94 = _RAND_739[3:0];
  _RAND_740 = {1{`RANDOM}};
  rob_n_flits_95 = _RAND_740[3:0];
  _RAND_741 = {1{`RANDOM}};
  rob_n_flits_96 = _RAND_741[3:0];
  _RAND_742 = {1{`RANDOM}};
  rob_n_flits_97 = _RAND_742[3:0];
  _RAND_743 = {1{`RANDOM}};
  rob_n_flits_98 = _RAND_743[3:0];
  _RAND_744 = {1{`RANDOM}};
  rob_n_flits_99 = _RAND_744[3:0];
  _RAND_745 = {1{`RANDOM}};
  rob_n_flits_100 = _RAND_745[3:0];
  _RAND_746 = {1{`RANDOM}};
  rob_n_flits_101 = _RAND_746[3:0];
  _RAND_747 = {1{`RANDOM}};
  rob_n_flits_102 = _RAND_747[3:0];
  _RAND_748 = {1{`RANDOM}};
  rob_n_flits_103 = _RAND_748[3:0];
  _RAND_749 = {1{`RANDOM}};
  rob_n_flits_104 = _RAND_749[3:0];
  _RAND_750 = {1{`RANDOM}};
  rob_n_flits_105 = _RAND_750[3:0];
  _RAND_751 = {1{`RANDOM}};
  rob_n_flits_106 = _RAND_751[3:0];
  _RAND_752 = {1{`RANDOM}};
  rob_n_flits_107 = _RAND_752[3:0];
  _RAND_753 = {1{`RANDOM}};
  rob_n_flits_108 = _RAND_753[3:0];
  _RAND_754 = {1{`RANDOM}};
  rob_n_flits_109 = _RAND_754[3:0];
  _RAND_755 = {1{`RANDOM}};
  rob_n_flits_110 = _RAND_755[3:0];
  _RAND_756 = {1{`RANDOM}};
  rob_n_flits_111 = _RAND_756[3:0];
  _RAND_757 = {1{`RANDOM}};
  rob_n_flits_112 = _RAND_757[3:0];
  _RAND_758 = {1{`RANDOM}};
  rob_n_flits_113 = _RAND_758[3:0];
  _RAND_759 = {1{`RANDOM}};
  rob_n_flits_114 = _RAND_759[3:0];
  _RAND_760 = {1{`RANDOM}};
  rob_n_flits_115 = _RAND_760[3:0];
  _RAND_761 = {1{`RANDOM}};
  rob_n_flits_116 = _RAND_761[3:0];
  _RAND_762 = {1{`RANDOM}};
  rob_n_flits_117 = _RAND_762[3:0];
  _RAND_763 = {1{`RANDOM}};
  rob_n_flits_118 = _RAND_763[3:0];
  _RAND_764 = {1{`RANDOM}};
  rob_n_flits_119 = _RAND_764[3:0];
  _RAND_765 = {1{`RANDOM}};
  rob_n_flits_120 = _RAND_765[3:0];
  _RAND_766 = {1{`RANDOM}};
  rob_n_flits_121 = _RAND_766[3:0];
  _RAND_767 = {1{`RANDOM}};
  rob_n_flits_122 = _RAND_767[3:0];
  _RAND_768 = {1{`RANDOM}};
  rob_n_flits_123 = _RAND_768[3:0];
  _RAND_769 = {1{`RANDOM}};
  rob_n_flits_124 = _RAND_769[3:0];
  _RAND_770 = {1{`RANDOM}};
  rob_n_flits_125 = _RAND_770[3:0];
  _RAND_771 = {1{`RANDOM}};
  rob_n_flits_126 = _RAND_771[3:0];
  _RAND_772 = {1{`RANDOM}};
  rob_n_flits_127 = _RAND_772[3:0];
  _RAND_773 = {1{`RANDOM}};
  rob_flits_returned_0 = _RAND_773[3:0];
  _RAND_774 = {1{`RANDOM}};
  rob_flits_returned_1 = _RAND_774[3:0];
  _RAND_775 = {1{`RANDOM}};
  rob_flits_returned_2 = _RAND_775[3:0];
  _RAND_776 = {1{`RANDOM}};
  rob_flits_returned_3 = _RAND_776[3:0];
  _RAND_777 = {1{`RANDOM}};
  rob_flits_returned_4 = _RAND_777[3:0];
  _RAND_778 = {1{`RANDOM}};
  rob_flits_returned_5 = _RAND_778[3:0];
  _RAND_779 = {1{`RANDOM}};
  rob_flits_returned_6 = _RAND_779[3:0];
  _RAND_780 = {1{`RANDOM}};
  rob_flits_returned_7 = _RAND_780[3:0];
  _RAND_781 = {1{`RANDOM}};
  rob_flits_returned_8 = _RAND_781[3:0];
  _RAND_782 = {1{`RANDOM}};
  rob_flits_returned_9 = _RAND_782[3:0];
  _RAND_783 = {1{`RANDOM}};
  rob_flits_returned_10 = _RAND_783[3:0];
  _RAND_784 = {1{`RANDOM}};
  rob_flits_returned_11 = _RAND_784[3:0];
  _RAND_785 = {1{`RANDOM}};
  rob_flits_returned_12 = _RAND_785[3:0];
  _RAND_786 = {1{`RANDOM}};
  rob_flits_returned_13 = _RAND_786[3:0];
  _RAND_787 = {1{`RANDOM}};
  rob_flits_returned_14 = _RAND_787[3:0];
  _RAND_788 = {1{`RANDOM}};
  rob_flits_returned_15 = _RAND_788[3:0];
  _RAND_789 = {1{`RANDOM}};
  rob_flits_returned_16 = _RAND_789[3:0];
  _RAND_790 = {1{`RANDOM}};
  rob_flits_returned_17 = _RAND_790[3:0];
  _RAND_791 = {1{`RANDOM}};
  rob_flits_returned_18 = _RAND_791[3:0];
  _RAND_792 = {1{`RANDOM}};
  rob_flits_returned_19 = _RAND_792[3:0];
  _RAND_793 = {1{`RANDOM}};
  rob_flits_returned_20 = _RAND_793[3:0];
  _RAND_794 = {1{`RANDOM}};
  rob_flits_returned_21 = _RAND_794[3:0];
  _RAND_795 = {1{`RANDOM}};
  rob_flits_returned_22 = _RAND_795[3:0];
  _RAND_796 = {1{`RANDOM}};
  rob_flits_returned_23 = _RAND_796[3:0];
  _RAND_797 = {1{`RANDOM}};
  rob_flits_returned_24 = _RAND_797[3:0];
  _RAND_798 = {1{`RANDOM}};
  rob_flits_returned_25 = _RAND_798[3:0];
  _RAND_799 = {1{`RANDOM}};
  rob_flits_returned_26 = _RAND_799[3:0];
  _RAND_800 = {1{`RANDOM}};
  rob_flits_returned_27 = _RAND_800[3:0];
  _RAND_801 = {1{`RANDOM}};
  rob_flits_returned_28 = _RAND_801[3:0];
  _RAND_802 = {1{`RANDOM}};
  rob_flits_returned_29 = _RAND_802[3:0];
  _RAND_803 = {1{`RANDOM}};
  rob_flits_returned_30 = _RAND_803[3:0];
  _RAND_804 = {1{`RANDOM}};
  rob_flits_returned_31 = _RAND_804[3:0];
  _RAND_805 = {1{`RANDOM}};
  rob_flits_returned_32 = _RAND_805[3:0];
  _RAND_806 = {1{`RANDOM}};
  rob_flits_returned_33 = _RAND_806[3:0];
  _RAND_807 = {1{`RANDOM}};
  rob_flits_returned_34 = _RAND_807[3:0];
  _RAND_808 = {1{`RANDOM}};
  rob_flits_returned_35 = _RAND_808[3:0];
  _RAND_809 = {1{`RANDOM}};
  rob_flits_returned_36 = _RAND_809[3:0];
  _RAND_810 = {1{`RANDOM}};
  rob_flits_returned_37 = _RAND_810[3:0];
  _RAND_811 = {1{`RANDOM}};
  rob_flits_returned_38 = _RAND_811[3:0];
  _RAND_812 = {1{`RANDOM}};
  rob_flits_returned_39 = _RAND_812[3:0];
  _RAND_813 = {1{`RANDOM}};
  rob_flits_returned_40 = _RAND_813[3:0];
  _RAND_814 = {1{`RANDOM}};
  rob_flits_returned_41 = _RAND_814[3:0];
  _RAND_815 = {1{`RANDOM}};
  rob_flits_returned_42 = _RAND_815[3:0];
  _RAND_816 = {1{`RANDOM}};
  rob_flits_returned_43 = _RAND_816[3:0];
  _RAND_817 = {1{`RANDOM}};
  rob_flits_returned_44 = _RAND_817[3:0];
  _RAND_818 = {1{`RANDOM}};
  rob_flits_returned_45 = _RAND_818[3:0];
  _RAND_819 = {1{`RANDOM}};
  rob_flits_returned_46 = _RAND_819[3:0];
  _RAND_820 = {1{`RANDOM}};
  rob_flits_returned_47 = _RAND_820[3:0];
  _RAND_821 = {1{`RANDOM}};
  rob_flits_returned_48 = _RAND_821[3:0];
  _RAND_822 = {1{`RANDOM}};
  rob_flits_returned_49 = _RAND_822[3:0];
  _RAND_823 = {1{`RANDOM}};
  rob_flits_returned_50 = _RAND_823[3:0];
  _RAND_824 = {1{`RANDOM}};
  rob_flits_returned_51 = _RAND_824[3:0];
  _RAND_825 = {1{`RANDOM}};
  rob_flits_returned_52 = _RAND_825[3:0];
  _RAND_826 = {1{`RANDOM}};
  rob_flits_returned_53 = _RAND_826[3:0];
  _RAND_827 = {1{`RANDOM}};
  rob_flits_returned_54 = _RAND_827[3:0];
  _RAND_828 = {1{`RANDOM}};
  rob_flits_returned_55 = _RAND_828[3:0];
  _RAND_829 = {1{`RANDOM}};
  rob_flits_returned_56 = _RAND_829[3:0];
  _RAND_830 = {1{`RANDOM}};
  rob_flits_returned_57 = _RAND_830[3:0];
  _RAND_831 = {1{`RANDOM}};
  rob_flits_returned_58 = _RAND_831[3:0];
  _RAND_832 = {1{`RANDOM}};
  rob_flits_returned_59 = _RAND_832[3:0];
  _RAND_833 = {1{`RANDOM}};
  rob_flits_returned_60 = _RAND_833[3:0];
  _RAND_834 = {1{`RANDOM}};
  rob_flits_returned_61 = _RAND_834[3:0];
  _RAND_835 = {1{`RANDOM}};
  rob_flits_returned_62 = _RAND_835[3:0];
  _RAND_836 = {1{`RANDOM}};
  rob_flits_returned_63 = _RAND_836[3:0];
  _RAND_837 = {1{`RANDOM}};
  rob_flits_returned_64 = _RAND_837[3:0];
  _RAND_838 = {1{`RANDOM}};
  rob_flits_returned_65 = _RAND_838[3:0];
  _RAND_839 = {1{`RANDOM}};
  rob_flits_returned_66 = _RAND_839[3:0];
  _RAND_840 = {1{`RANDOM}};
  rob_flits_returned_67 = _RAND_840[3:0];
  _RAND_841 = {1{`RANDOM}};
  rob_flits_returned_68 = _RAND_841[3:0];
  _RAND_842 = {1{`RANDOM}};
  rob_flits_returned_69 = _RAND_842[3:0];
  _RAND_843 = {1{`RANDOM}};
  rob_flits_returned_70 = _RAND_843[3:0];
  _RAND_844 = {1{`RANDOM}};
  rob_flits_returned_71 = _RAND_844[3:0];
  _RAND_845 = {1{`RANDOM}};
  rob_flits_returned_72 = _RAND_845[3:0];
  _RAND_846 = {1{`RANDOM}};
  rob_flits_returned_73 = _RAND_846[3:0];
  _RAND_847 = {1{`RANDOM}};
  rob_flits_returned_74 = _RAND_847[3:0];
  _RAND_848 = {1{`RANDOM}};
  rob_flits_returned_75 = _RAND_848[3:0];
  _RAND_849 = {1{`RANDOM}};
  rob_flits_returned_76 = _RAND_849[3:0];
  _RAND_850 = {1{`RANDOM}};
  rob_flits_returned_77 = _RAND_850[3:0];
  _RAND_851 = {1{`RANDOM}};
  rob_flits_returned_78 = _RAND_851[3:0];
  _RAND_852 = {1{`RANDOM}};
  rob_flits_returned_79 = _RAND_852[3:0];
  _RAND_853 = {1{`RANDOM}};
  rob_flits_returned_80 = _RAND_853[3:0];
  _RAND_854 = {1{`RANDOM}};
  rob_flits_returned_81 = _RAND_854[3:0];
  _RAND_855 = {1{`RANDOM}};
  rob_flits_returned_82 = _RAND_855[3:0];
  _RAND_856 = {1{`RANDOM}};
  rob_flits_returned_83 = _RAND_856[3:0];
  _RAND_857 = {1{`RANDOM}};
  rob_flits_returned_84 = _RAND_857[3:0];
  _RAND_858 = {1{`RANDOM}};
  rob_flits_returned_85 = _RAND_858[3:0];
  _RAND_859 = {1{`RANDOM}};
  rob_flits_returned_86 = _RAND_859[3:0];
  _RAND_860 = {1{`RANDOM}};
  rob_flits_returned_87 = _RAND_860[3:0];
  _RAND_861 = {1{`RANDOM}};
  rob_flits_returned_88 = _RAND_861[3:0];
  _RAND_862 = {1{`RANDOM}};
  rob_flits_returned_89 = _RAND_862[3:0];
  _RAND_863 = {1{`RANDOM}};
  rob_flits_returned_90 = _RAND_863[3:0];
  _RAND_864 = {1{`RANDOM}};
  rob_flits_returned_91 = _RAND_864[3:0];
  _RAND_865 = {1{`RANDOM}};
  rob_flits_returned_92 = _RAND_865[3:0];
  _RAND_866 = {1{`RANDOM}};
  rob_flits_returned_93 = _RAND_866[3:0];
  _RAND_867 = {1{`RANDOM}};
  rob_flits_returned_94 = _RAND_867[3:0];
  _RAND_868 = {1{`RANDOM}};
  rob_flits_returned_95 = _RAND_868[3:0];
  _RAND_869 = {1{`RANDOM}};
  rob_flits_returned_96 = _RAND_869[3:0];
  _RAND_870 = {1{`RANDOM}};
  rob_flits_returned_97 = _RAND_870[3:0];
  _RAND_871 = {1{`RANDOM}};
  rob_flits_returned_98 = _RAND_871[3:0];
  _RAND_872 = {1{`RANDOM}};
  rob_flits_returned_99 = _RAND_872[3:0];
  _RAND_873 = {1{`RANDOM}};
  rob_flits_returned_100 = _RAND_873[3:0];
  _RAND_874 = {1{`RANDOM}};
  rob_flits_returned_101 = _RAND_874[3:0];
  _RAND_875 = {1{`RANDOM}};
  rob_flits_returned_102 = _RAND_875[3:0];
  _RAND_876 = {1{`RANDOM}};
  rob_flits_returned_103 = _RAND_876[3:0];
  _RAND_877 = {1{`RANDOM}};
  rob_flits_returned_104 = _RAND_877[3:0];
  _RAND_878 = {1{`RANDOM}};
  rob_flits_returned_105 = _RAND_878[3:0];
  _RAND_879 = {1{`RANDOM}};
  rob_flits_returned_106 = _RAND_879[3:0];
  _RAND_880 = {1{`RANDOM}};
  rob_flits_returned_107 = _RAND_880[3:0];
  _RAND_881 = {1{`RANDOM}};
  rob_flits_returned_108 = _RAND_881[3:0];
  _RAND_882 = {1{`RANDOM}};
  rob_flits_returned_109 = _RAND_882[3:0];
  _RAND_883 = {1{`RANDOM}};
  rob_flits_returned_110 = _RAND_883[3:0];
  _RAND_884 = {1{`RANDOM}};
  rob_flits_returned_111 = _RAND_884[3:0];
  _RAND_885 = {1{`RANDOM}};
  rob_flits_returned_112 = _RAND_885[3:0];
  _RAND_886 = {1{`RANDOM}};
  rob_flits_returned_113 = _RAND_886[3:0];
  _RAND_887 = {1{`RANDOM}};
  rob_flits_returned_114 = _RAND_887[3:0];
  _RAND_888 = {1{`RANDOM}};
  rob_flits_returned_115 = _RAND_888[3:0];
  _RAND_889 = {1{`RANDOM}};
  rob_flits_returned_116 = _RAND_889[3:0];
  _RAND_890 = {1{`RANDOM}};
  rob_flits_returned_117 = _RAND_890[3:0];
  _RAND_891 = {1{`RANDOM}};
  rob_flits_returned_118 = _RAND_891[3:0];
  _RAND_892 = {1{`RANDOM}};
  rob_flits_returned_119 = _RAND_892[3:0];
  _RAND_893 = {1{`RANDOM}};
  rob_flits_returned_120 = _RAND_893[3:0];
  _RAND_894 = {1{`RANDOM}};
  rob_flits_returned_121 = _RAND_894[3:0];
  _RAND_895 = {1{`RANDOM}};
  rob_flits_returned_122 = _RAND_895[3:0];
  _RAND_896 = {1{`RANDOM}};
  rob_flits_returned_123 = _RAND_896[3:0];
  _RAND_897 = {1{`RANDOM}};
  rob_flits_returned_124 = _RAND_897[3:0];
  _RAND_898 = {1{`RANDOM}};
  rob_flits_returned_125 = _RAND_898[3:0];
  _RAND_899 = {1{`RANDOM}};
  rob_flits_returned_126 = _RAND_899[3:0];
  _RAND_900 = {1{`RANDOM}};
  rob_flits_returned_127 = _RAND_900[3:0];
  _RAND_901 = {2{`RANDOM}};
  rob_tscs_0 = _RAND_901[63:0];
  _RAND_902 = {2{`RANDOM}};
  rob_tscs_1 = _RAND_902[63:0];
  _RAND_903 = {2{`RANDOM}};
  rob_tscs_2 = _RAND_903[63:0];
  _RAND_904 = {2{`RANDOM}};
  rob_tscs_3 = _RAND_904[63:0];
  _RAND_905 = {2{`RANDOM}};
  rob_tscs_4 = _RAND_905[63:0];
  _RAND_906 = {2{`RANDOM}};
  rob_tscs_5 = _RAND_906[63:0];
  _RAND_907 = {2{`RANDOM}};
  rob_tscs_6 = _RAND_907[63:0];
  _RAND_908 = {2{`RANDOM}};
  rob_tscs_7 = _RAND_908[63:0];
  _RAND_909 = {2{`RANDOM}};
  rob_tscs_8 = _RAND_909[63:0];
  _RAND_910 = {2{`RANDOM}};
  rob_tscs_9 = _RAND_910[63:0];
  _RAND_911 = {2{`RANDOM}};
  rob_tscs_10 = _RAND_911[63:0];
  _RAND_912 = {2{`RANDOM}};
  rob_tscs_11 = _RAND_912[63:0];
  _RAND_913 = {2{`RANDOM}};
  rob_tscs_12 = _RAND_913[63:0];
  _RAND_914 = {2{`RANDOM}};
  rob_tscs_13 = _RAND_914[63:0];
  _RAND_915 = {2{`RANDOM}};
  rob_tscs_14 = _RAND_915[63:0];
  _RAND_916 = {2{`RANDOM}};
  rob_tscs_15 = _RAND_916[63:0];
  _RAND_917 = {2{`RANDOM}};
  rob_tscs_16 = _RAND_917[63:0];
  _RAND_918 = {2{`RANDOM}};
  rob_tscs_17 = _RAND_918[63:0];
  _RAND_919 = {2{`RANDOM}};
  rob_tscs_18 = _RAND_919[63:0];
  _RAND_920 = {2{`RANDOM}};
  rob_tscs_19 = _RAND_920[63:0];
  _RAND_921 = {2{`RANDOM}};
  rob_tscs_20 = _RAND_921[63:0];
  _RAND_922 = {2{`RANDOM}};
  rob_tscs_21 = _RAND_922[63:0];
  _RAND_923 = {2{`RANDOM}};
  rob_tscs_22 = _RAND_923[63:0];
  _RAND_924 = {2{`RANDOM}};
  rob_tscs_23 = _RAND_924[63:0];
  _RAND_925 = {2{`RANDOM}};
  rob_tscs_24 = _RAND_925[63:0];
  _RAND_926 = {2{`RANDOM}};
  rob_tscs_25 = _RAND_926[63:0];
  _RAND_927 = {2{`RANDOM}};
  rob_tscs_26 = _RAND_927[63:0];
  _RAND_928 = {2{`RANDOM}};
  rob_tscs_27 = _RAND_928[63:0];
  _RAND_929 = {2{`RANDOM}};
  rob_tscs_28 = _RAND_929[63:0];
  _RAND_930 = {2{`RANDOM}};
  rob_tscs_29 = _RAND_930[63:0];
  _RAND_931 = {2{`RANDOM}};
  rob_tscs_30 = _RAND_931[63:0];
  _RAND_932 = {2{`RANDOM}};
  rob_tscs_31 = _RAND_932[63:0];
  _RAND_933 = {2{`RANDOM}};
  rob_tscs_32 = _RAND_933[63:0];
  _RAND_934 = {2{`RANDOM}};
  rob_tscs_33 = _RAND_934[63:0];
  _RAND_935 = {2{`RANDOM}};
  rob_tscs_34 = _RAND_935[63:0];
  _RAND_936 = {2{`RANDOM}};
  rob_tscs_35 = _RAND_936[63:0];
  _RAND_937 = {2{`RANDOM}};
  rob_tscs_36 = _RAND_937[63:0];
  _RAND_938 = {2{`RANDOM}};
  rob_tscs_37 = _RAND_938[63:0];
  _RAND_939 = {2{`RANDOM}};
  rob_tscs_38 = _RAND_939[63:0];
  _RAND_940 = {2{`RANDOM}};
  rob_tscs_39 = _RAND_940[63:0];
  _RAND_941 = {2{`RANDOM}};
  rob_tscs_40 = _RAND_941[63:0];
  _RAND_942 = {2{`RANDOM}};
  rob_tscs_41 = _RAND_942[63:0];
  _RAND_943 = {2{`RANDOM}};
  rob_tscs_42 = _RAND_943[63:0];
  _RAND_944 = {2{`RANDOM}};
  rob_tscs_43 = _RAND_944[63:0];
  _RAND_945 = {2{`RANDOM}};
  rob_tscs_44 = _RAND_945[63:0];
  _RAND_946 = {2{`RANDOM}};
  rob_tscs_45 = _RAND_946[63:0];
  _RAND_947 = {2{`RANDOM}};
  rob_tscs_46 = _RAND_947[63:0];
  _RAND_948 = {2{`RANDOM}};
  rob_tscs_47 = _RAND_948[63:0];
  _RAND_949 = {2{`RANDOM}};
  rob_tscs_48 = _RAND_949[63:0];
  _RAND_950 = {2{`RANDOM}};
  rob_tscs_49 = _RAND_950[63:0];
  _RAND_951 = {2{`RANDOM}};
  rob_tscs_50 = _RAND_951[63:0];
  _RAND_952 = {2{`RANDOM}};
  rob_tscs_51 = _RAND_952[63:0];
  _RAND_953 = {2{`RANDOM}};
  rob_tscs_52 = _RAND_953[63:0];
  _RAND_954 = {2{`RANDOM}};
  rob_tscs_53 = _RAND_954[63:0];
  _RAND_955 = {2{`RANDOM}};
  rob_tscs_54 = _RAND_955[63:0];
  _RAND_956 = {2{`RANDOM}};
  rob_tscs_55 = _RAND_956[63:0];
  _RAND_957 = {2{`RANDOM}};
  rob_tscs_56 = _RAND_957[63:0];
  _RAND_958 = {2{`RANDOM}};
  rob_tscs_57 = _RAND_958[63:0];
  _RAND_959 = {2{`RANDOM}};
  rob_tscs_58 = _RAND_959[63:0];
  _RAND_960 = {2{`RANDOM}};
  rob_tscs_59 = _RAND_960[63:0];
  _RAND_961 = {2{`RANDOM}};
  rob_tscs_60 = _RAND_961[63:0];
  _RAND_962 = {2{`RANDOM}};
  rob_tscs_61 = _RAND_962[63:0];
  _RAND_963 = {2{`RANDOM}};
  rob_tscs_62 = _RAND_963[63:0];
  _RAND_964 = {2{`RANDOM}};
  rob_tscs_63 = _RAND_964[63:0];
  _RAND_965 = {2{`RANDOM}};
  rob_tscs_64 = _RAND_965[63:0];
  _RAND_966 = {2{`RANDOM}};
  rob_tscs_65 = _RAND_966[63:0];
  _RAND_967 = {2{`RANDOM}};
  rob_tscs_66 = _RAND_967[63:0];
  _RAND_968 = {2{`RANDOM}};
  rob_tscs_67 = _RAND_968[63:0];
  _RAND_969 = {2{`RANDOM}};
  rob_tscs_68 = _RAND_969[63:0];
  _RAND_970 = {2{`RANDOM}};
  rob_tscs_69 = _RAND_970[63:0];
  _RAND_971 = {2{`RANDOM}};
  rob_tscs_70 = _RAND_971[63:0];
  _RAND_972 = {2{`RANDOM}};
  rob_tscs_71 = _RAND_972[63:0];
  _RAND_973 = {2{`RANDOM}};
  rob_tscs_72 = _RAND_973[63:0];
  _RAND_974 = {2{`RANDOM}};
  rob_tscs_73 = _RAND_974[63:0];
  _RAND_975 = {2{`RANDOM}};
  rob_tscs_74 = _RAND_975[63:0];
  _RAND_976 = {2{`RANDOM}};
  rob_tscs_75 = _RAND_976[63:0];
  _RAND_977 = {2{`RANDOM}};
  rob_tscs_76 = _RAND_977[63:0];
  _RAND_978 = {2{`RANDOM}};
  rob_tscs_77 = _RAND_978[63:0];
  _RAND_979 = {2{`RANDOM}};
  rob_tscs_78 = _RAND_979[63:0];
  _RAND_980 = {2{`RANDOM}};
  rob_tscs_79 = _RAND_980[63:0];
  _RAND_981 = {2{`RANDOM}};
  rob_tscs_80 = _RAND_981[63:0];
  _RAND_982 = {2{`RANDOM}};
  rob_tscs_81 = _RAND_982[63:0];
  _RAND_983 = {2{`RANDOM}};
  rob_tscs_82 = _RAND_983[63:0];
  _RAND_984 = {2{`RANDOM}};
  rob_tscs_83 = _RAND_984[63:0];
  _RAND_985 = {2{`RANDOM}};
  rob_tscs_84 = _RAND_985[63:0];
  _RAND_986 = {2{`RANDOM}};
  rob_tscs_85 = _RAND_986[63:0];
  _RAND_987 = {2{`RANDOM}};
  rob_tscs_86 = _RAND_987[63:0];
  _RAND_988 = {2{`RANDOM}};
  rob_tscs_87 = _RAND_988[63:0];
  _RAND_989 = {2{`RANDOM}};
  rob_tscs_88 = _RAND_989[63:0];
  _RAND_990 = {2{`RANDOM}};
  rob_tscs_89 = _RAND_990[63:0];
  _RAND_991 = {2{`RANDOM}};
  rob_tscs_90 = _RAND_991[63:0];
  _RAND_992 = {2{`RANDOM}};
  rob_tscs_91 = _RAND_992[63:0];
  _RAND_993 = {2{`RANDOM}};
  rob_tscs_92 = _RAND_993[63:0];
  _RAND_994 = {2{`RANDOM}};
  rob_tscs_93 = _RAND_994[63:0];
  _RAND_995 = {2{`RANDOM}};
  rob_tscs_94 = _RAND_995[63:0];
  _RAND_996 = {2{`RANDOM}};
  rob_tscs_95 = _RAND_996[63:0];
  _RAND_997 = {2{`RANDOM}};
  rob_tscs_96 = _RAND_997[63:0];
  _RAND_998 = {2{`RANDOM}};
  rob_tscs_97 = _RAND_998[63:0];
  _RAND_999 = {2{`RANDOM}};
  rob_tscs_98 = _RAND_999[63:0];
  _RAND_1000 = {2{`RANDOM}};
  rob_tscs_99 = _RAND_1000[63:0];
  _RAND_1001 = {2{`RANDOM}};
  rob_tscs_100 = _RAND_1001[63:0];
  _RAND_1002 = {2{`RANDOM}};
  rob_tscs_101 = _RAND_1002[63:0];
  _RAND_1003 = {2{`RANDOM}};
  rob_tscs_102 = _RAND_1003[63:0];
  _RAND_1004 = {2{`RANDOM}};
  rob_tscs_103 = _RAND_1004[63:0];
  _RAND_1005 = {2{`RANDOM}};
  rob_tscs_104 = _RAND_1005[63:0];
  _RAND_1006 = {2{`RANDOM}};
  rob_tscs_105 = _RAND_1006[63:0];
  _RAND_1007 = {2{`RANDOM}};
  rob_tscs_106 = _RAND_1007[63:0];
  _RAND_1008 = {2{`RANDOM}};
  rob_tscs_107 = _RAND_1008[63:0];
  _RAND_1009 = {2{`RANDOM}};
  rob_tscs_108 = _RAND_1009[63:0];
  _RAND_1010 = {2{`RANDOM}};
  rob_tscs_109 = _RAND_1010[63:0];
  _RAND_1011 = {2{`RANDOM}};
  rob_tscs_110 = _RAND_1011[63:0];
  _RAND_1012 = {2{`RANDOM}};
  rob_tscs_111 = _RAND_1012[63:0];
  _RAND_1013 = {2{`RANDOM}};
  rob_tscs_112 = _RAND_1013[63:0];
  _RAND_1014 = {2{`RANDOM}};
  rob_tscs_113 = _RAND_1014[63:0];
  _RAND_1015 = {2{`RANDOM}};
  rob_tscs_114 = _RAND_1015[63:0];
  _RAND_1016 = {2{`RANDOM}};
  rob_tscs_115 = _RAND_1016[63:0];
  _RAND_1017 = {2{`RANDOM}};
  rob_tscs_116 = _RAND_1017[63:0];
  _RAND_1018 = {2{`RANDOM}};
  rob_tscs_117 = _RAND_1018[63:0];
  _RAND_1019 = {2{`RANDOM}};
  rob_tscs_118 = _RAND_1019[63:0];
  _RAND_1020 = {2{`RANDOM}};
  rob_tscs_119 = _RAND_1020[63:0];
  _RAND_1021 = {2{`RANDOM}};
  rob_tscs_120 = _RAND_1021[63:0];
  _RAND_1022 = {2{`RANDOM}};
  rob_tscs_121 = _RAND_1022[63:0];
  _RAND_1023 = {2{`RANDOM}};
  rob_tscs_122 = _RAND_1023[63:0];
  _RAND_1024 = {2{`RANDOM}};
  rob_tscs_123 = _RAND_1024[63:0];
  _RAND_1025 = {2{`RANDOM}};
  rob_tscs_124 = _RAND_1025[63:0];
  _RAND_1026 = {2{`RANDOM}};
  rob_tscs_125 = _RAND_1026[63:0];
  _RAND_1027 = {2{`RANDOM}};
  rob_tscs_126 = _RAND_1027[63:0];
  _RAND_1028 = {2{`RANDOM}};
  rob_tscs_127 = _RAND_1028[63:0];
  _RAND_1029 = {1{`RANDOM}};
  io_success_REG = _RAND_1029[0:0];
  _RAND_1030 = {1{`RANDOM}};
  packet_valid = _RAND_1030[0:0];
  _RAND_1031 = {1{`RANDOM}};
  packet_rob_idx = _RAND_1031[6:0];
  _RAND_1032 = {1{`RANDOM}};
  packet_valid_1 = _RAND_1032[0:0];
  _RAND_1033 = {1{`RANDOM}};
  packet_rob_idx_1 = _RAND_1033[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(~idle_counter[10]); // @[TestHarness.scala 148:9]
    end
    //
    if (_T_84 & _T_3) begin
      assert(_T_42[0]); // @[TestHarness.scala 201:13]
    end
    //
    if (_T_84 & _T_3) begin
      assert(_T_48 == io_from_noc_0_flit_bits_payload); // @[TestHarness.scala 202:13]
    end
    //
    if (_T_84 & _T_3) begin
      assert(io_from_noc_0_flit_bits_ingress_id == _GEN_4608); // @[TestHarness.scala 203:13]
    end
    //
    if (_T_84 & _T_3) begin
      assert(~_GEN_4736); // @[TestHarness.scala 204:13]
    end
    //
    if (_T_84 & _T_3) begin
      assert(_GEN_4864 < _GEN_4992); // @[TestHarness.scala 205:13]
    end
    //
    if (_T_84 & _T_3) begin
      assert(~packet_valid & io_from_noc_0_flit_bits_head | out_payload_rob_idx == _GEN_7819); // @[TestHarness.scala 206:13]
    end
    //
    if (_T_131 & _T_3) begin
      assert(_T_89[0]); // @[TestHarness.scala 201:13]
    end
    //
    if (_T_131 & _T_3) begin
      assert(_T_95 == io_from_noc_1_flit_bits_payload); // @[TestHarness.scala 202:13]
    end
    //
    if (_T_131 & _T_3) begin
      assert(io_from_noc_1_flit_bits_ingress_id == _GEN_6405); // @[TestHarness.scala 203:13]
    end
    //
    if (_T_131 & _T_3) begin
      assert(7'h7f == out_payload_1_rob_idx[6:0] ? rob_egress_id_127 : _GEN_6532); // @[TestHarness.scala 204:13]
    end
    //
    if (_T_131 & _T_3) begin
      assert(_GEN_6661 < _GEN_6789); // @[TestHarness.scala 205:13]
    end
    //
    if (_T_131 & _T_3) begin
      assert(~packet_valid_1 & io_from_noc_1_flit_bits_head | out_payload_1_rob_idx == _GEN_7820); // @[TestHarness.scala 206:13]
    end
    //
    if (rob_valids[0] & _T_3) begin
      assert(_T_136 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[1] & _T_3) begin
      assert(_T_143 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[2] & _T_3) begin
      assert(_T_150 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[3] & _T_3) begin
      assert(_T_157 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[4] & _T_3) begin
      assert(_T_164 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[5] & _T_3) begin
      assert(_T_171 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[6] & _T_3) begin
      assert(_T_178 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[7] & _T_3) begin
      assert(_T_185 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[8] & _T_3) begin
      assert(_T_192 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[9] & _T_3) begin
      assert(_T_199 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[10] & _T_3) begin
      assert(_T_206 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[11] & _T_3) begin
      assert(_T_213 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[12] & _T_3) begin
      assert(_T_220 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[13] & _T_3) begin
      assert(_T_227 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[14] & _T_3) begin
      assert(_T_234 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[15] & _T_3) begin
      assert(_T_241 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[16] & _T_3) begin
      assert(_T_248 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[17] & _T_3) begin
      assert(_T_255 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[18] & _T_3) begin
      assert(_T_262 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[19] & _T_3) begin
      assert(_T_269 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[20] & _T_3) begin
      assert(_T_276 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[21] & _T_3) begin
      assert(_T_283 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[22] & _T_3) begin
      assert(_T_290 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[23] & _T_3) begin
      assert(_T_297 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[24] & _T_3) begin
      assert(_T_304 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[25] & _T_3) begin
      assert(_T_311 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[26] & _T_3) begin
      assert(_T_318 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[27] & _T_3) begin
      assert(_T_325 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[28] & _T_3) begin
      assert(_T_332 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[29] & _T_3) begin
      assert(_T_339 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[30] & _T_3) begin
      assert(_T_346 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[31] & _T_3) begin
      assert(_T_353 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[32] & _T_3) begin
      assert(_T_360 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[33] & _T_3) begin
      assert(_T_367 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[34] & _T_3) begin
      assert(_T_374 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[35] & _T_3) begin
      assert(_T_381 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[36] & _T_3) begin
      assert(_T_388 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[37] & _T_3) begin
      assert(_T_395 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[38] & _T_3) begin
      assert(_T_402 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[39] & _T_3) begin
      assert(_T_409 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[40] & _T_3) begin
      assert(_T_416 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[41] & _T_3) begin
      assert(_T_423 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[42] & _T_3) begin
      assert(_T_430 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[43] & _T_3) begin
      assert(_T_437 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[44] & _T_3) begin
      assert(_T_444 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[45] & _T_3) begin
      assert(_T_451 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[46] & _T_3) begin
      assert(_T_458 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[47] & _T_3) begin
      assert(_T_465 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[48] & _T_3) begin
      assert(_T_472 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[49] & _T_3) begin
      assert(_T_479 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[50] & _T_3) begin
      assert(_T_486 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[51] & _T_3) begin
      assert(_T_493 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[52] & _T_3) begin
      assert(_T_500 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[53] & _T_3) begin
      assert(_T_507 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[54] & _T_3) begin
      assert(_T_514 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[55] & _T_3) begin
      assert(_T_521 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[56] & _T_3) begin
      assert(_T_528 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[57] & _T_3) begin
      assert(_T_535 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[58] & _T_3) begin
      assert(_T_542 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[59] & _T_3) begin
      assert(_T_549 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[60] & _T_3) begin
      assert(_T_556 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[61] & _T_3) begin
      assert(_T_563 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[62] & _T_3) begin
      assert(_T_570 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[63] & _T_3) begin
      assert(_T_577 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[64] & _T_3) begin
      assert(_T_584 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[65] & _T_3) begin
      assert(_T_591 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[66] & _T_3) begin
      assert(_T_598 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[67] & _T_3) begin
      assert(_T_605 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[68] & _T_3) begin
      assert(_T_612 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[69] & _T_3) begin
      assert(_T_619 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[70] & _T_3) begin
      assert(_T_626 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[71] & _T_3) begin
      assert(_T_633 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[72] & _T_3) begin
      assert(_T_640 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[73] & _T_3) begin
      assert(_T_647 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[74] & _T_3) begin
      assert(_T_654 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[75] & _T_3) begin
      assert(_T_661 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[76] & _T_3) begin
      assert(_T_668 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[77] & _T_3) begin
      assert(_T_675 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[78] & _T_3) begin
      assert(_T_682 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[79] & _T_3) begin
      assert(_T_689 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[80] & _T_3) begin
      assert(_T_696 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[81] & _T_3) begin
      assert(_T_703 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[82] & _T_3) begin
      assert(_T_710 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[83] & _T_3) begin
      assert(_T_717 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[84] & _T_3) begin
      assert(_T_724 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[85] & _T_3) begin
      assert(_T_731 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[86] & _T_3) begin
      assert(_T_738 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[87] & _T_3) begin
      assert(_T_745 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[88] & _T_3) begin
      assert(_T_752 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[89] & _T_3) begin
      assert(_T_759 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[90] & _T_3) begin
      assert(_T_766 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[91] & _T_3) begin
      assert(_T_773 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[92] & _T_3) begin
      assert(_T_780 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[93] & _T_3) begin
      assert(_T_787 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[94] & _T_3) begin
      assert(_T_794 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[95] & _T_3) begin
      assert(_T_801 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[96] & _T_3) begin
      assert(_T_808 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[97] & _T_3) begin
      assert(_T_815 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[98] & _T_3) begin
      assert(_T_822 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[99] & _T_3) begin
      assert(_T_829 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[100] & _T_3) begin
      assert(_T_836 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[101] & _T_3) begin
      assert(_T_843 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[102] & _T_3) begin
      assert(_T_850 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[103] & _T_3) begin
      assert(_T_857 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[104] & _T_3) begin
      assert(_T_864 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[105] & _T_3) begin
      assert(_T_871 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[106] & _T_3) begin
      assert(_T_878 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[107] & _T_3) begin
      assert(_T_885 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[108] & _T_3) begin
      assert(_T_892 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[109] & _T_3) begin
      assert(_T_899 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[110] & _T_3) begin
      assert(_T_906 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[111] & _T_3) begin
      assert(_T_913 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[112] & _T_3) begin
      assert(_T_920 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[113] & _T_3) begin
      assert(_T_927 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[114] & _T_3) begin
      assert(_T_934 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[115] & _T_3) begin
      assert(_T_941 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[116] & _T_3) begin
      assert(_T_948 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[117] & _T_3) begin
      assert(_T_955 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[118] & _T_3) begin
      assert(_T_962 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[119] & _T_3) begin
      assert(_T_969 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[120] & _T_3) begin
      assert(_T_976 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[121] & _T_3) begin
      assert(_T_983 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[122] & _T_3) begin
      assert(_T_990 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[123] & _T_3) begin
      assert(_T_997 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[124] & _T_3) begin
      assert(_T_1004 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[125] & _T_3) begin
      assert(_T_1011 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[126] & _T_3) begin
      assert(_T_1018 < 64'h4000); // @[TestHarness.scala 229:13]
    end
    //
    if (rob_valids[127] & _T_3) begin
      assert(_T_1025 < 64'h4000); // @[TestHarness.scala 229:13]
    end
  end
endmodule
module TestHarness(
  input   clock,
  input   reset,
  output  io_success
);
  wire  lazyNoC_clock; // @[TestHarness.scala 238:19]
  wire  lazyNoC_reset; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_ingress_1_flit_ready; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_ingress_1_flit_valid; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_ingress_1_flit_bits_head; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_ingress_1_flit_bits_tail; // @[TestHarness.scala 238:19]
  wire [63:0] lazyNoC_io_ingress_1_flit_bits_payload; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_ingress_1_flit_bits_egress_id; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_ingress_0_flit_ready; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_ingress_0_flit_valid; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_ingress_0_flit_bits_head; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_ingress_0_flit_bits_tail; // @[TestHarness.scala 238:19]
  wire [63:0] lazyNoC_io_ingress_0_flit_bits_payload; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_ingress_0_flit_bits_egress_id; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_egress_1_flit_valid; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_egress_1_flit_bits_head; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_egress_1_flit_bits_tail; // @[TestHarness.scala 238:19]
  wire [63:0] lazyNoC_io_egress_1_flit_bits_payload; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_egress_1_flit_bits_ingress_id; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_egress_0_flit_valid; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_egress_0_flit_bits_head; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_egress_0_flit_bits_tail; // @[TestHarness.scala 238:19]
  wire [63:0] lazyNoC_io_egress_0_flit_bits_payload; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_egress_0_flit_bits_ingress_id; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_router_clocks_0_clock; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_router_clocks_0_reset; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_router_clocks_1_clock; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_router_clocks_1_reset; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_router_clocks_2_clock; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_router_clocks_2_reset; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_router_clocks_3_clock; // @[TestHarness.scala 238:19]
  wire  lazyNoC_io_router_clocks_3_reset; // @[TestHarness.scala 238:19]
  wire  noc_tester_clock; // @[TestHarness.scala 269:26]
  wire  noc_tester_reset; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_to_noc_1_flit_ready; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_to_noc_1_flit_valid; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_to_noc_1_flit_bits_head; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_to_noc_1_flit_bits_tail; // @[TestHarness.scala 269:26]
  wire [63:0] noc_tester_io_to_noc_1_flit_bits_payload; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_to_noc_1_flit_bits_egress_id; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_to_noc_0_flit_ready; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_to_noc_0_flit_valid; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_to_noc_0_flit_bits_head; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_to_noc_0_flit_bits_tail; // @[TestHarness.scala 269:26]
  wire [63:0] noc_tester_io_to_noc_0_flit_bits_payload; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_to_noc_0_flit_bits_egress_id; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_from_noc_1_flit_ready; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_from_noc_1_flit_valid; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_from_noc_1_flit_bits_head; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_from_noc_1_flit_bits_tail; // @[TestHarness.scala 269:26]
  wire [63:0] noc_tester_io_from_noc_1_flit_bits_payload; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_from_noc_1_flit_bits_ingress_id; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_from_noc_0_flit_ready; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_from_noc_0_flit_valid; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_from_noc_0_flit_bits_head; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_from_noc_0_flit_bits_tail; // @[TestHarness.scala 269:26]
  wire [63:0] noc_tester_io_from_noc_0_flit_bits_payload; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_from_noc_0_flit_bits_ingress_id; // @[TestHarness.scala 269:26]
  wire  noc_tester_io_success; // @[TestHarness.scala 269:26]
  NoC lazyNoC ( // @[TestHarness.scala 238:19]
    .clock(lazyNoC_clock),
    .reset(lazyNoC_reset),
    .io_ingress_1_flit_ready(lazyNoC_io_ingress_1_flit_ready),
    .io_ingress_1_flit_valid(lazyNoC_io_ingress_1_flit_valid),
    .io_ingress_1_flit_bits_head(lazyNoC_io_ingress_1_flit_bits_head),
    .io_ingress_1_flit_bits_tail(lazyNoC_io_ingress_1_flit_bits_tail),
    .io_ingress_1_flit_bits_payload(lazyNoC_io_ingress_1_flit_bits_payload),
    .io_ingress_1_flit_bits_egress_id(lazyNoC_io_ingress_1_flit_bits_egress_id),
    .io_ingress_0_flit_ready(lazyNoC_io_ingress_0_flit_ready),
    .io_ingress_0_flit_valid(lazyNoC_io_ingress_0_flit_valid),
    .io_ingress_0_flit_bits_head(lazyNoC_io_ingress_0_flit_bits_head),
    .io_ingress_0_flit_bits_tail(lazyNoC_io_ingress_0_flit_bits_tail),
    .io_ingress_0_flit_bits_payload(lazyNoC_io_ingress_0_flit_bits_payload),
    .io_ingress_0_flit_bits_egress_id(lazyNoC_io_ingress_0_flit_bits_egress_id),
    .io_egress_1_flit_valid(lazyNoC_io_egress_1_flit_valid),
    .io_egress_1_flit_bits_head(lazyNoC_io_egress_1_flit_bits_head),
    .io_egress_1_flit_bits_tail(lazyNoC_io_egress_1_flit_bits_tail),
    .io_egress_1_flit_bits_payload(lazyNoC_io_egress_1_flit_bits_payload),
    .io_egress_1_flit_bits_ingress_id(lazyNoC_io_egress_1_flit_bits_ingress_id),
    .io_egress_0_flit_valid(lazyNoC_io_egress_0_flit_valid),
    .io_egress_0_flit_bits_head(lazyNoC_io_egress_0_flit_bits_head),
    .io_egress_0_flit_bits_tail(lazyNoC_io_egress_0_flit_bits_tail),
    .io_egress_0_flit_bits_payload(lazyNoC_io_egress_0_flit_bits_payload),
    .io_egress_0_flit_bits_ingress_id(lazyNoC_io_egress_0_flit_bits_ingress_id),
    .io_router_clocks_0_clock(lazyNoC_io_router_clocks_0_clock),
    .io_router_clocks_0_reset(lazyNoC_io_router_clocks_0_reset),
    .io_router_clocks_1_clock(lazyNoC_io_router_clocks_1_clock),
    .io_router_clocks_1_reset(lazyNoC_io_router_clocks_1_reset),
    .io_router_clocks_2_clock(lazyNoC_io_router_clocks_2_clock),
    .io_router_clocks_2_reset(lazyNoC_io_router_clocks_2_reset),
    .io_router_clocks_3_clock(lazyNoC_io_router_clocks_3_clock),
    .io_router_clocks_3_reset(lazyNoC_io_router_clocks_3_reset)
  );
  NoCTester noc_tester ( // @[TestHarness.scala 269:26]
    .clock(noc_tester_clock),
    .reset(noc_tester_reset),
    .io_to_noc_1_flit_ready(noc_tester_io_to_noc_1_flit_ready),
    .io_to_noc_1_flit_valid(noc_tester_io_to_noc_1_flit_valid),
    .io_to_noc_1_flit_bits_head(noc_tester_io_to_noc_1_flit_bits_head),
    .io_to_noc_1_flit_bits_tail(noc_tester_io_to_noc_1_flit_bits_tail),
    .io_to_noc_1_flit_bits_payload(noc_tester_io_to_noc_1_flit_bits_payload),
    .io_to_noc_1_flit_bits_egress_id(noc_tester_io_to_noc_1_flit_bits_egress_id),
    .io_to_noc_0_flit_ready(noc_tester_io_to_noc_0_flit_ready),
    .io_to_noc_0_flit_valid(noc_tester_io_to_noc_0_flit_valid),
    .io_to_noc_0_flit_bits_head(noc_tester_io_to_noc_0_flit_bits_head),
    .io_to_noc_0_flit_bits_tail(noc_tester_io_to_noc_0_flit_bits_tail),
    .io_to_noc_0_flit_bits_payload(noc_tester_io_to_noc_0_flit_bits_payload),
    .io_to_noc_0_flit_bits_egress_id(noc_tester_io_to_noc_0_flit_bits_egress_id),
    .io_from_noc_1_flit_ready(noc_tester_io_from_noc_1_flit_ready),
    .io_from_noc_1_flit_valid(noc_tester_io_from_noc_1_flit_valid),
    .io_from_noc_1_flit_bits_head(noc_tester_io_from_noc_1_flit_bits_head),
    .io_from_noc_1_flit_bits_tail(noc_tester_io_from_noc_1_flit_bits_tail),
    .io_from_noc_1_flit_bits_payload(noc_tester_io_from_noc_1_flit_bits_payload),
    .io_from_noc_1_flit_bits_ingress_id(noc_tester_io_from_noc_1_flit_bits_ingress_id),
    .io_from_noc_0_flit_ready(noc_tester_io_from_noc_0_flit_ready),
    .io_from_noc_0_flit_valid(noc_tester_io_from_noc_0_flit_valid),
    .io_from_noc_0_flit_bits_head(noc_tester_io_from_noc_0_flit_bits_head),
    .io_from_noc_0_flit_bits_tail(noc_tester_io_from_noc_0_flit_bits_tail),
    .io_from_noc_0_flit_bits_payload(noc_tester_io_from_noc_0_flit_bits_payload),
    .io_from_noc_0_flit_bits_ingress_id(noc_tester_io_from_noc_0_flit_bits_ingress_id),
    .io_success(noc_tester_io_success)
  );
  assign io_success = noc_tester_io_success; // @[TestHarness.scala 272:14]
  assign lazyNoC_clock = clock;
  assign lazyNoC_reset = reset;
  assign lazyNoC_io_ingress_1_flit_valid = noc_tester_io_to_noc_1_flit_valid; // @[TestHarness.scala 270:18]
  assign lazyNoC_io_ingress_1_flit_bits_head = noc_tester_io_to_noc_1_flit_bits_head; // @[TestHarness.scala 270:18]
  assign lazyNoC_io_ingress_1_flit_bits_tail = noc_tester_io_to_noc_1_flit_bits_tail; // @[TestHarness.scala 270:18]
  assign lazyNoC_io_ingress_1_flit_bits_payload = noc_tester_io_to_noc_1_flit_bits_payload; // @[TestHarness.scala 270:18]
  assign lazyNoC_io_ingress_1_flit_bits_egress_id = noc_tester_io_to_noc_1_flit_bits_egress_id; // @[TestHarness.scala 270:18]
  assign lazyNoC_io_ingress_0_flit_valid = noc_tester_io_to_noc_0_flit_valid; // @[TestHarness.scala 270:18]
  assign lazyNoC_io_ingress_0_flit_bits_head = noc_tester_io_to_noc_0_flit_bits_head; // @[TestHarness.scala 270:18]
  assign lazyNoC_io_ingress_0_flit_bits_tail = noc_tester_io_to_noc_0_flit_bits_tail; // @[TestHarness.scala 270:18]
  assign lazyNoC_io_ingress_0_flit_bits_payload = noc_tester_io_to_noc_0_flit_bits_payload; // @[TestHarness.scala 270:18]
  assign lazyNoC_io_ingress_0_flit_bits_egress_id = noc_tester_io_to_noc_0_flit_bits_egress_id; // @[TestHarness.scala 270:18]
  assign lazyNoC_io_router_clocks_0_clock = clock; // @[TestHarness.scala 239:40]
  assign lazyNoC_io_router_clocks_0_reset = reset; // @[TestHarness.scala 240:40]
  assign lazyNoC_io_router_clocks_1_clock = clock; // @[TestHarness.scala 239:40]
  assign lazyNoC_io_router_clocks_1_reset = reset; // @[TestHarness.scala 240:40]
  assign lazyNoC_io_router_clocks_2_clock = clock; // @[TestHarness.scala 239:40]
  assign lazyNoC_io_router_clocks_2_reset = reset; // @[TestHarness.scala 240:40]
  assign lazyNoC_io_router_clocks_3_clock = clock; // @[TestHarness.scala 239:40]
  assign lazyNoC_io_router_clocks_3_reset = reset; // @[TestHarness.scala 240:40]
  assign noc_tester_clock = clock;
  assign noc_tester_reset = reset;
  assign noc_tester_io_to_noc_1_flit_ready = lazyNoC_io_ingress_1_flit_ready; // @[TestHarness.scala 270:18]
  assign noc_tester_io_to_noc_0_flit_ready = lazyNoC_io_ingress_0_flit_ready; // @[TestHarness.scala 270:18]
  assign noc_tester_io_from_noc_1_flit_valid = lazyNoC_io_egress_1_flit_valid; // @[TestHarness.scala 271:26]
  assign noc_tester_io_from_noc_1_flit_bits_head = lazyNoC_io_egress_1_flit_bits_head; // @[TestHarness.scala 271:26]
  assign noc_tester_io_from_noc_1_flit_bits_tail = lazyNoC_io_egress_1_flit_bits_tail; // @[TestHarness.scala 271:26]
  assign noc_tester_io_from_noc_1_flit_bits_payload = lazyNoC_io_egress_1_flit_bits_payload; // @[TestHarness.scala 271:26]
  assign noc_tester_io_from_noc_1_flit_bits_ingress_id = lazyNoC_io_egress_1_flit_bits_ingress_id; // @[TestHarness.scala 271:26]
  assign noc_tester_io_from_noc_0_flit_valid = lazyNoC_io_egress_0_flit_valid; // @[TestHarness.scala 271:26]
  assign noc_tester_io_from_noc_0_flit_bits_head = lazyNoC_io_egress_0_flit_bits_head; // @[TestHarness.scala 271:26]
  assign noc_tester_io_from_noc_0_flit_bits_tail = lazyNoC_io_egress_0_flit_bits_tail; // @[TestHarness.scala 271:26]
  assign noc_tester_io_from_noc_0_flit_bits_payload = lazyNoC_io_egress_0_flit_bits_payload; // @[TestHarness.scala 271:26]
  assign noc_tester_io_from_noc_0_flit_bits_ingress_id = lazyNoC_io_egress_0_flit_bits_ingress_id; // @[TestHarness.scala 271:26]
endmodule
module NoCChiselTester(
  input   clock,
  input   reset
);
  wire  th_clock; // @[NocTests.scala 11:18]
  wire  th_reset; // @[NocTests.scala 11:18]
  wire  th_io_success; // @[NocTests.scala 11:18]
  TestHarness th ( // @[NocTests.scala 11:18]
    .clock(th_clock),
    .reset(th_reset),
    .io_success(th_io_success)
  );
  assign th_clock = clock;
  assign th_reset = reset;
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (th_io_success & ~reset) begin
          $finish; // @[NocTests.scala 12:30]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
